magic
tech scmos
timestamp
<< pdiffusion >>
rect	92	57	98	63
rect	20	149	26	155
rect	20	9	26	15
rect	53	149	59	155
rect	79	82	85	88
rect	26	101	32	107
rect	98	82	104	88
rect	70	130	76	136
rect	13	9	19	15
rect	0	101	6	107
rect	10	101	16	107
rect	22	82	28	88
rect	76	57	82	63
rect	16	26	22	32
rect	30	149	36	155
rect	10	149	16	155
rect	0	57	6	63
rect	60	9	66	15
rect	3	130	9	136
rect	41	82	47	88
rect	77	130	83	136
rect	33	9	39	15
rect	35	130	41	136
rect	16	57	22	63
rect	42	26	48	32
rect	57	82	63	88
rect	23	26	29	32
rect	16	130	22	136
rect	0	26	6	32
rect	3	82	9	88
rect	51	57	57	63
rect	45	130	51	136
rect	38	57	44	63
rect	78	26	84	32
rect	46	9	52	15
rect	55	101	61	107
rect	68	26	74	32
rect	83	101	89	107
rect	46	149	52	155
rect	108	57	114	63
rect	53	9	59	15
rect	0	149	6	155
rect	0	9	6	15
rect	58	26	64	32
rect	45	101	51	107
rect	9	130	12	136
rect	82	57	85	63
rect	57	57	60	63
rect	85	57	88	63
rect	60	57	63	63
rect	47	82	50	88
rect	51	130	54	136
rect	63	82	66	88
rect	36	149	39	155
rect	54	130	57	136
rect	57	130	60	136
rect	63	57	66	63
rect	22	130	25	136
rect	44	57	47	63
rect	12	130	15	136
rect	85	82	88	88
rect	26	9	29	15
rect	60	130	63	136
rect	22	57	25	63
rect	66	82	69	88
rect	9	82	12	88
rect	6	9	9	15
rect	6	26	9	32
rect	63	130	66	136
rect	12	82	15	88
rect	9	26	12	32
rect	48	26	51	32
rect	25	130	28	136
rect	29	9	32	15
rect	29	26	32	32
rect	26	149	29	155
rect	16	149	19	155
rect	104	101	107	107
rect	16	101	19	107
rect	88	57	91	63
rect	98	57	101	63
rect	32	101	35	107
rect	64	26	67	32
rect	69	82	72	88
rect	72	82	75	88
rect	61	101	64	107
rect	64	101	67	107
rect	66	130	69	136
rect	67	101	70	107
rect	70	101	73	107
rect	51	26	54	32
rect	35	101	38	107
rect	19	101	22	107
rect	66	57	69	63
rect	73	101	76	107
rect	28	82	31	88
rect	69	57	72	63
rect	25	57	28	63
rect	6	57	9	63
rect	76	101	79	107
rect	28	57	31	63
rect	22	101	25	107
rect	28	130	31	136
rect	126	82	129	88
rect	15	82	18	88
rect	89	26	92	32
rect	99	26	102	32
rect	79	101	82	107
rect	50	82	53	88
rect	41	130	44	136
rect	51	101	54	107
rect	88	82	91	88
rect	91	82	94	88
rect	39	9	42	15
rect	31	82	34	88
rect	34	82	37	88
rect	94	82	97	88
rect	38	101	41	107
rect	32	26	35	32
rect	0	82	3	88
rect	75	82	78	88
rect	37	82	40	88
rect	18	82	21	88
rect	148	57	151	63
rect	9	57	12	63
rect	94	9	97	15
rect	39	149	42	155
rect	53	82	56	88
rect	101	57	104	63
rect	104	57	107	63
rect	31	57	34	63
rect	34	57	37	63
rect	31	130	34	136
rect	42	9	45	15
rect	6	101	9	107
rect	72	57	75	63
rect	41	101	44	107
rect	12	57	15	63
rect	47	57	50	63
rect	117	26	120	32
rect	35	26	38	32
rect	38	26	41	32
rect	42	149	45	155
rect	0	130	3	136
rect	74	26	77	32
rect	12	26	15	32
rect	54	26	57	32
rect	6	149	9	155
rect	78	9	81	15
rect	9	9	12	15
