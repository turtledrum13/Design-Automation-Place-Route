magic
tech scmos
timestamp
<< pdiffusion >>
rect	0	11	6	17
rect	0	105	6	111
rect	17	11	23	17
rect	56	105	62	111
rect	0	51	6	57
rect	0	159	6	165
rect	29	51	35	57
rect	20	159	26	165
rect	10	11	16	17
rect	31	105	37	111
rect	27	11	33	17
rect	78	105	84	111
rect	13	51	19	57
rect	10	159	16	165
rect	54	51	60	57
rect	27	159	33	165
rect	0	26	6	32
rect	0	134	6	140
rect	17	26	23	32
rect	35	134	41	140
rect	0	78	6	84
rect	3	178	9	184
rect	35	78	41	84
rect	37	11	43	17
rect	94	105	100	111
rect	60	11	66	17
rect	123	105	129	111
rect	82	51	88	57
rect	37	159	43	165
rect	105	51	111	57
rect	51	159	57	165
rect	47	11	53	17
rect	107	105	113	111
rect	73	11	79	17
rect	130	105	136	111
rect	95	51	101	57
rect	44	159	50	165
rect	112	51	118	57
rect	67	159	73	165
rect	46	26	52	32
rect	82	134	88	140
rect	75	26	81	32
rect	105	134	111	140
rect	67	78	73	84
rect	31	178	37	184
rect	65	26	68	32
rect	6	51	9	57
rect	23	26	26	32
rect	111	134	114	140
rect	6	11	9	17
rect	9	51	12	57
rect	55	134	58	140
rect	41	134	44	140
rect	66	11	69	17
rect	57	159	60	165
rect	53	11	56	17
rect	113	105	116	111
rect	101	134	104	140
rect	31	26	34	32
rect	41	78	44	84
rect	60	51	63	57
rect	116	105	119	111
rect	6	105	9	111
rect	19	51	22	57
rect	23	11	26	17
rect	44	78	47	84
rect	16	159	19	165
rect	88	51	91	57
rect	127	78	130	84
rect	26	26	29	32
rect	14	134	17	140
rect	34	26	37	32
rect	37	105	40	111
rect	33	11	36	17
rect	59	134	62	140
rect	28	134	31	140
rect	100	105	103	111
rect	40	105	43	111
rect	0	178	3	184
rect	69	134	72	140
rect	62	134	65	140
rect	9	105	12	111
rect	33	159	36	165
rect	31	134	34	140
rect	56	11	59	17
rect	6	159	9	165
rect	91	51	94	57
rect	63	51	66	57
rect	66	51	69	57
rect	10	78	13	84
rect	22	51	25	57
rect	136	105	139	111
rect	7	26	10	32
rect	13	78	16	84
rect	62	105	65	111
rect	65	105	68	111
rect	68	26	71	32
rect	88	134	91	140
rect	93	134	96	140
rect	119	105	122	111
rect	35	51	38	57
rect	73	78	76	84
rect	117	78	120	84
rect	7	134	10	140
rect	38	51	41	57
rect	23	134	26	140
rect	107	78	110	84
rect	41	51	44	57
rect	12	105	15	111
rect	44	51	47	57
rect	84	105	87	111
rect	15	105	18	111
rect	72	134	75	140
rect	87	105	90	111
rect	16	78	19	84
rect	44	134	47	140
rect	43	105	46	111
rect	60	26	63	32
rect	10	134	13	140
rect	113	78	116	84
rect	88	78	91	84
rect	91	78	94	84
rect	18	105	21	111
rect	47	78	50	84
rect	140	78	143	84
rect	21	105	24	111
rect	76	78	79	84
rect	69	51	72	57
rect	90	105	93	111
rect	91	159	94	165
rect	123	78	126	84
rect	101	51	104	57
rect	24	105	27	111
rect	57	78	60	84
rect	19	78	22	84
rect	79	78	82	84
rect	6	78	9	84
rect	60	159	63	165
rect	46	105	49	111
rect	50	78	53	84
rect	72	51	75	57
rect	27	105	30	111
rect	103	105	106	111
rect	68	105	71	111
rect	71	105	74	111
rect	19	134	22	140
rect	49	105	52	111
rect	75	51	78	57
rect	82	78	85	84
rect	94	78	97	84
rect	127	51	130	57
rect	102	26	105	32
rect	25	78	28	84
rect	52	105	55	111
rect	25	51	28	57
rect	53	78	56	84
rect	78	51	81	57
rect	28	78	31	84
rect	75	134	78	140
rect	78	134	81	140
rect	50	134	53	140
rect	71	26	74	32
rect	74	105	77	111
rect	131	26	134	32
rect	47	51	50	57
rect	82	26	85	32
rect	50	51	53	57
rect	76	159	79	165
rect	79	159	82	165
rect	69	11	72	17
rect	65	134	68	140
rect	52	26	55	32
rect	42	26	45	32
rect	77	178	80	184
rect	63	159	66	165
rect	43	11	46	17
