magic
tech scmos
timestamp
<< pdiffusion >>
rect	8	0	9	1
rect	8	1	9	2
rect	8	2	9	3
rect	8	3	9	4
rect	8	4	9	5
rect	8	5	9	6
rect	8	6	9	7
rect	8	7	9	8
rect	8	8	9	9
rect	8	9	9	10
rect	8	10	9	11
rect	8	11	9	12
rect	8	13	9	14
rect	8	14	9	15
rect	8	15	9	16
rect	8	18	9	19
rect	8	21	9	22
rect	8	24	9	25
rect	8	27	9	28
rect	8	28	9	29
rect	8	29	9	30
rect	8	30	9	31
rect	8	31	9	32
rect	8	32	9	33
rect	8	33	9	34
rect	8	36	9	37
rect	8	37	9	38
rect	8	38	9	39
rect	8	39	9	40
rect	8	40	9	41
rect	8	41	9	42
rect	8	42	9	43
rect	8	43	9	44
rect	8	44	9	45
rect	8	45	9	46
rect	8	46	9	47
rect	8	47	9	48
rect	8	49	9	50
rect	8	50	9	51
rect	8	51	9	52
rect	8	52	9	53
rect	8	56	9	57
rect	8	57	9	58
rect	8	60	9	61
rect	8	61	9	62
rect	8	62	9	63
rect	8	63	9	64
rect	8	64	9	65
rect	8	65	9	66
rect	8	66	9	67
rect	8	67	9	68
rect	8	69	9	70
rect	8	70	9	71
rect	8	71	9	72
rect	8	76	9	77
rect	8	77	9	78
rect	8	78	9	79
rect	8	79	9	80
rect	8	82	9	83
rect	8	86	9	87
rect	8	87	9	88
rect	8	88	9	89
rect	8	89	9	90
rect	8	90	9	91
rect	8	91	9	92
rect	8	92	9	93
rect	8	93	9	94
rect	8	94	9	95
rect	8	96	9	97
rect	8	97	9	98
rect	8	98	9	99
rect	8	99	9	100
rect	8	100	9	101
rect	8	101	9	102
rect	8	102	9	103
rect	8	103	9	104
rect	8	104	9	105
rect	9	0	10	1
rect	9	1	10	2
rect	9	2	10	3
rect	9	3	10	4
rect	9	4	10	5
rect	9	5	10	6
rect	9	6	10	7
rect	9	7	10	8
rect	9	8	10	9
rect	9	9	10	10
rect	9	10	10	11
rect	9	11	10	12
rect	9	13	10	14
rect	9	14	10	15
rect	9	15	10	16
rect	9	18	10	19
rect	9	21	10	22
rect	9	24	10	25
rect	9	27	10	28
rect	9	28	10	29
rect	9	29	10	30
rect	9	30	10	31
rect	9	31	10	32
rect	9	32	10	33
rect	9	33	10	34
rect	9	36	10	37
rect	9	37	10	38
rect	9	38	10	39
rect	9	39	10	40
rect	9	40	10	41
rect	9	41	10	42
rect	9	42	10	43
rect	9	43	10	44
rect	9	44	10	45
rect	9	45	10	46
rect	9	46	10	47
rect	9	47	10	48
rect	9	49	10	50
rect	9	50	10	51
rect	9	51	10	52
rect	9	52	10	53
rect	9	56	10	57
rect	9	57	10	58
rect	9	60	10	61
rect	9	61	10	62
rect	9	62	10	63
rect	9	63	10	64
rect	9	64	10	65
rect	9	65	10	66
rect	9	66	10	67
rect	9	67	10	68
rect	9	69	10	70
rect	9	70	10	71
rect	9	71	10	72
rect	9	76	10	77
rect	9	77	10	78
rect	9	78	10	79
rect	9	79	10	80
rect	9	82	10	83
rect	9	86	10	87
rect	9	87	10	88
rect	9	88	10	89
rect	9	89	10	90
rect	9	90	10	91
rect	9	91	10	92
rect	9	92	10	93
rect	9	93	10	94
rect	9	94	10	95
rect	9	96	10	97
rect	9	97	10	98
rect	9	98	10	99
rect	9	99	10	100
rect	9	100	10	101
rect	9	101	10	102
rect	9	102	10	103
rect	9	103	10	104
rect	9	104	10	105
rect	10	0	11	1
rect	10	1	11	2
rect	10	2	11	3
rect	10	3	11	4
rect	10	4	11	5
rect	10	5	11	6
rect	10	6	11	7
rect	10	7	11	8
rect	10	8	11	9
rect	10	9	11	10
rect	10	10	11	11
rect	10	11	11	12
rect	10	13	11	14
rect	10	14	11	15
rect	10	15	11	16
rect	10	18	11	19
rect	10	21	11	22
rect	10	24	11	25
rect	10	27	11	28
rect	10	28	11	29
rect	10	29	11	30
rect	10	30	11	31
rect	10	31	11	32
rect	10	32	11	33
rect	10	33	11	34
rect	10	36	11	37
rect	10	37	11	38
rect	10	38	11	39
rect	10	39	11	40
rect	10	40	11	41
rect	10	41	11	42
rect	10	42	11	43
rect	10	43	11	44
rect	10	44	11	45
rect	10	45	11	46
rect	10	46	11	47
rect	10	47	11	48
rect	10	49	11	50
rect	10	50	11	51
rect	10	51	11	52
rect	10	52	11	53
rect	10	56	11	57
rect	10	57	11	58
rect	10	60	11	61
rect	10	61	11	62
rect	10	62	11	63
rect	10	63	11	64
rect	10	64	11	65
rect	10	65	11	66
rect	10	66	11	67
rect	10	67	11	68
rect	10	69	11	70
rect	10	70	11	71
rect	10	71	11	72
rect	10	76	11	77
rect	10	77	11	78
rect	10	78	11	79
rect	10	79	11	80
rect	10	82	11	83
rect	10	86	11	87
rect	10	87	11	88
rect	10	88	11	89
rect	10	89	11	90
rect	10	90	11	91
rect	10	91	11	92
rect	10	92	11	93
rect	10	93	11	94
rect	10	94	11	95
rect	10	96	11	97
rect	10	97	11	98
rect	10	98	11	99
rect	10	99	11	100
rect	10	100	11	101
rect	10	101	11	102
rect	10	102	11	103
rect	10	103	11	104
rect	10	104	11	105
rect	11	0	12	1
rect	11	1	12	2
rect	11	2	12	3
rect	11	3	12	4
rect	11	4	12	5
rect	11	5	12	6
rect	11	6	12	7
rect	11	7	12	8
rect	11	8	12	9
rect	11	9	12	10
rect	11	10	12	11
rect	11	11	12	12
rect	11	13	12	14
rect	11	14	12	15
rect	11	15	12	16
rect	11	18	12	19
rect	11	21	12	22
rect	11	24	12	25
rect	11	27	12	28
rect	11	28	12	29
rect	11	29	12	30
rect	11	30	12	31
rect	11	31	12	32
rect	11	32	12	33
rect	11	33	12	34
rect	11	36	12	37
rect	11	37	12	38
rect	11	38	12	39
rect	11	39	12	40
rect	11	40	12	41
rect	11	41	12	42
rect	11	42	12	43
rect	11	43	12	44
rect	11	44	12	45
rect	11	45	12	46
rect	11	46	12	47
rect	11	47	12	48
rect	11	49	12	50
rect	11	50	12	51
rect	11	51	12	52
rect	11	52	12	53
rect	11	56	12	57
rect	11	57	12	58
rect	11	60	12	61
rect	11	61	12	62
rect	11	62	12	63
rect	11	63	12	64
rect	11	64	12	65
rect	11	65	12	66
rect	11	66	12	67
rect	11	67	12	68
rect	11	69	12	70
rect	11	70	12	71
rect	11	71	12	72
rect	11	76	12	77
rect	11	77	12	78
rect	11	78	12	79
rect	11	79	12	80
rect	11	82	12	83
rect	11	86	12	87
rect	11	87	12	88
rect	11	88	12	89
rect	11	89	12	90
rect	11	90	12	91
rect	11	91	12	92
rect	11	92	12	93
rect	11	93	12	94
rect	11	94	12	95
rect	11	96	12	97
rect	11	97	12	98
rect	11	98	12	99
rect	11	99	12	100
rect	11	100	12	101
rect	11	101	12	102
rect	11	102	12	103
rect	11	103	12	104
rect	11	104	12	105
rect	12	0	13	1
rect	12	1	13	2
rect	12	2	13	3
rect	12	3	13	4
rect	12	4	13	5
rect	12	5	13	6
rect	12	6	13	7
rect	12	7	13	8
rect	12	8	13	9
rect	12	9	13	10
rect	12	10	13	11
rect	12	11	13	12
rect	12	13	13	14
rect	12	14	13	15
rect	12	15	13	16
rect	12	18	13	19
rect	12	21	13	22
rect	12	24	13	25
rect	12	27	13	28
rect	12	28	13	29
rect	12	29	13	30
rect	12	30	13	31
rect	12	31	13	32
rect	12	32	13	33
rect	12	33	13	34
rect	12	36	13	37
rect	12	37	13	38
rect	12	38	13	39
rect	12	39	13	40
rect	12	40	13	41
rect	12	41	13	42
rect	12	42	13	43
rect	12	43	13	44
rect	12	44	13	45
rect	12	45	13	46
rect	12	46	13	47
rect	12	47	13	48
rect	12	49	13	50
rect	12	50	13	51
rect	12	51	13	52
rect	12	52	13	53
rect	12	56	13	57
rect	12	57	13	58
rect	12	60	13	61
rect	12	61	13	62
rect	12	62	13	63
rect	12	63	13	64
rect	12	64	13	65
rect	12	65	13	66
rect	12	66	13	67
rect	12	67	13	68
rect	12	69	13	70
rect	12	70	13	71
rect	12	71	13	72
rect	12	76	13	77
rect	12	77	13	78
rect	12	78	13	79
rect	12	79	13	80
rect	12	82	13	83
rect	12	86	13	87
rect	12	87	13	88
rect	12	88	13	89
rect	12	89	13	90
rect	12	90	13	91
rect	12	91	13	92
rect	12	92	13	93
rect	12	93	13	94
rect	12	94	13	95
rect	12	96	13	97
rect	12	97	13	98
rect	12	98	13	99
rect	12	99	13	100
rect	12	100	13	101
rect	12	101	13	102
rect	12	102	13	103
rect	12	103	13	104
rect	12	104	13	105
rect	13	0	14	1
rect	13	1	14	2
rect	13	2	14	3
rect	13	3	14	4
rect	13	4	14	5
rect	13	5	14	6
rect	13	6	14	7
rect	13	7	14	8
rect	13	8	14	9
rect	13	9	14	10
rect	13	10	14	11
rect	13	11	14	12
rect	13	13	14	14
rect	13	14	14	15
rect	13	15	14	16
rect	13	18	14	19
rect	13	21	14	22
rect	13	24	14	25
rect	13	27	14	28
rect	13	28	14	29
rect	13	29	14	30
rect	13	30	14	31
rect	13	31	14	32
rect	13	32	14	33
rect	13	33	14	34
rect	13	36	14	37
rect	13	37	14	38
rect	13	38	14	39
rect	13	39	14	40
rect	13	40	14	41
rect	13	41	14	42
rect	13	42	14	43
rect	13	43	14	44
rect	13	44	14	45
rect	13	45	14	46
rect	13	46	14	47
rect	13	47	14	48
rect	13	49	14	50
rect	13	50	14	51
rect	13	51	14	52
rect	13	52	14	53
rect	13	56	14	57
rect	13	57	14	58
rect	13	60	14	61
rect	13	61	14	62
rect	13	62	14	63
rect	13	63	14	64
rect	13	64	14	65
rect	13	65	14	66
rect	13	66	14	67
rect	13	67	14	68
rect	13	69	14	70
rect	13	70	14	71
rect	13	71	14	72
rect	13	76	14	77
rect	13	77	14	78
rect	13	78	14	79
rect	13	79	14	80
rect	13	82	14	83
rect	13	86	14	87
rect	13	87	14	88
rect	13	88	14	89
rect	13	89	14	90
rect	13	90	14	91
rect	13	91	14	92
rect	13	92	14	93
rect	13	93	14	94
rect	13	94	14	95
rect	13	96	14	97
rect	13	97	14	98
rect	13	98	14	99
rect	13	99	14	100
rect	13	100	14	101
rect	13	101	14	102
rect	13	102	14	103
rect	13	103	14	104
rect	13	104	14	105
rect	31	0	32	1
rect	31	1	32	2
rect	31	2	32	3
rect	31	3	32	4
rect	31	4	32	5
rect	31	5	32	6
rect	31	6	32	7
rect	31	7	32	8
rect	31	8	32	9
rect	31	10	32	11
rect	31	11	32	12
rect	31	12	32	13
rect	31	13	32	14
rect	31	14	32	15
rect	31	15	32	16
rect	31	18	32	19
rect	31	21	32	22
rect	31	24	32	25
rect	31	27	32	28
rect	31	28	32	29
rect	31	29	32	30
rect	31	30	32	31
rect	31	31	32	32
rect	31	32	32	33
rect	31	33	32	34
rect	31	36	32	37
rect	31	37	32	38
rect	31	38	32	39
rect	31	39	32	40
rect	31	40	32	41
rect	31	41	32	42
rect	31	42	32	43
rect	31	43	32	44
rect	31	45	32	46
rect	31	46	32	47
rect	31	47	32	48
rect	31	48	32	49
rect	31	49	32	50
rect	31	50	32	51
rect	31	51	32	52
rect	31	52	32	53
rect	31	55	32	56
rect	31	56	32	57
rect	31	57	32	58
rect	31	60	32	61
rect	31	61	32	62
rect	31	62	32	63
rect	31	63	32	64
rect	31	64	32	65
rect	31	65	32	66
rect	31	67	32	68
rect	31	68	32	69
rect	31	69	32	70
rect	31	70	32	71
rect	31	71	32	72
rect	31	76	32	77
rect	31	77	32	78
rect	31	78	32	79
rect	31	79	32	80
rect	31	82	32	83
rect	31	86	32	87
rect	31	87	32	88
rect	31	88	32	89
rect	31	89	32	90
rect	31	90	32	91
rect	31	91	32	92
rect	31	92	32	93
rect	31	93	32	94
rect	31	94	32	95
rect	31	95	32	96
rect	31	96	32	97
rect	31	97	32	98
rect	31	98	32	99
rect	31	99	32	100
rect	31	100	32	101
rect	31	101	32	102
rect	31	102	32	103
rect	31	103	32	104
rect	31	105	32	106
rect	31	106	32	107
rect	31	107	32	108
rect	31	108	32	109
rect	31	109	32	110
rect	31	110	32	111
rect	31	111	32	112
rect	31	112	32	113
rect	31	113	32	114
rect	31	114	32	115
rect	31	115	32	116
rect	31	116	32	117
rect	31	118	32	119
rect	31	119	32	120
rect	31	120	32	121
rect	31	121	32	122
rect	31	122	32	123
rect	31	123	32	124
rect	31	125	32	126
rect	31	126	32	127
rect	31	127	32	128
rect	31	128	32	129
rect	31	129	32	130
rect	31	130	32	131
rect	31	131	32	132
rect	31	132	32	133
rect	31	133	32	134
rect	31	135	32	136
rect	31	136	32	137
rect	31	137	32	138
rect	31	138	32	139
rect	31	139	32	140
rect	31	140	32	141
rect	31	141	32	142
rect	31	142	32	143
rect	31	143	32	144
rect	32	0	33	1
rect	32	1	33	2
rect	32	2	33	3
rect	32	3	33	4
rect	32	4	33	5
rect	32	5	33	6
rect	32	6	33	7
rect	32	7	33	8
rect	32	8	33	9
rect	32	10	33	11
rect	32	11	33	12
rect	32	12	33	13
rect	32	13	33	14
rect	32	14	33	15
rect	32	15	33	16
rect	32	18	33	19
rect	32	21	33	22
rect	32	24	33	25
rect	32	27	33	28
rect	32	28	33	29
rect	32	29	33	30
rect	32	30	33	31
rect	32	31	33	32
rect	32	32	33	33
rect	32	33	33	34
rect	32	36	33	37
rect	32	37	33	38
rect	32	38	33	39
rect	32	39	33	40
rect	32	40	33	41
rect	32	41	33	42
rect	32	42	33	43
rect	32	43	33	44
rect	32	45	33	46
rect	32	46	33	47
rect	32	47	33	48
rect	32	48	33	49
rect	32	49	33	50
rect	32	50	33	51
rect	32	51	33	52
rect	32	52	33	53
rect	32	55	33	56
rect	32	56	33	57
rect	32	57	33	58
rect	32	60	33	61
rect	32	61	33	62
rect	32	62	33	63
rect	32	63	33	64
rect	32	64	33	65
rect	32	65	33	66
rect	32	67	33	68
rect	32	68	33	69
rect	32	69	33	70
rect	32	70	33	71
rect	32	71	33	72
rect	32	76	33	77
rect	32	77	33	78
rect	32	78	33	79
rect	32	79	33	80
rect	32	82	33	83
rect	32	86	33	87
rect	32	87	33	88
rect	32	88	33	89
rect	32	89	33	90
rect	32	90	33	91
rect	32	91	33	92
rect	32	92	33	93
rect	32	93	33	94
rect	32	94	33	95
rect	32	95	33	96
rect	32	96	33	97
rect	32	97	33	98
rect	32	98	33	99
rect	32	99	33	100
rect	32	100	33	101
rect	32	101	33	102
rect	32	102	33	103
rect	32	103	33	104
rect	32	105	33	106
rect	32	106	33	107
rect	32	107	33	108
rect	32	108	33	109
rect	32	109	33	110
rect	32	110	33	111
rect	32	111	33	112
rect	32	112	33	113
rect	32	113	33	114
rect	32	114	33	115
rect	32	115	33	116
rect	32	116	33	117
rect	32	118	33	119
rect	32	119	33	120
rect	32	120	33	121
rect	32	121	33	122
rect	32	122	33	123
rect	32	123	33	124
rect	32	125	33	126
rect	32	126	33	127
rect	32	127	33	128
rect	32	128	33	129
rect	32	129	33	130
rect	32	130	33	131
rect	32	131	33	132
rect	32	132	33	133
rect	32	133	33	134
rect	32	135	33	136
rect	32	136	33	137
rect	32	137	33	138
rect	32	138	33	139
rect	32	139	33	140
rect	32	140	33	141
rect	32	141	33	142
rect	32	142	33	143
rect	32	143	33	144
rect	33	0	34	1
rect	33	1	34	2
rect	33	2	34	3
rect	33	3	34	4
rect	33	4	34	5
rect	33	5	34	6
rect	33	6	34	7
rect	33	7	34	8
rect	33	8	34	9
rect	33	10	34	11
rect	33	11	34	12
rect	33	12	34	13
rect	33	13	34	14
rect	33	14	34	15
rect	33	15	34	16
rect	33	18	34	19
rect	33	21	34	22
rect	33	24	34	25
rect	33	27	34	28
rect	33	28	34	29
rect	33	29	34	30
rect	33	30	34	31
rect	33	31	34	32
rect	33	32	34	33
rect	33	33	34	34
rect	33	36	34	37
rect	33	37	34	38
rect	33	38	34	39
rect	33	39	34	40
rect	33	40	34	41
rect	33	41	34	42
rect	33	42	34	43
rect	33	43	34	44
rect	33	45	34	46
rect	33	46	34	47
rect	33	47	34	48
rect	33	48	34	49
rect	33	49	34	50
rect	33	50	34	51
rect	33	51	34	52
rect	33	52	34	53
rect	33	55	34	56
rect	33	56	34	57
rect	33	57	34	58
rect	33	60	34	61
rect	33	61	34	62
rect	33	62	34	63
rect	33	63	34	64
rect	33	64	34	65
rect	33	65	34	66
rect	33	67	34	68
rect	33	68	34	69
rect	33	69	34	70
rect	33	70	34	71
rect	33	71	34	72
rect	33	76	34	77
rect	33	77	34	78
rect	33	78	34	79
rect	33	79	34	80
rect	33	82	34	83
rect	33	86	34	87
rect	33	87	34	88
rect	33	88	34	89
rect	33	89	34	90
rect	33	90	34	91
rect	33	91	34	92
rect	33	92	34	93
rect	33	93	34	94
rect	33	94	34	95
rect	33	95	34	96
rect	33	96	34	97
rect	33	97	34	98
rect	33	98	34	99
rect	33	99	34	100
rect	33	100	34	101
rect	33	101	34	102
rect	33	102	34	103
rect	33	103	34	104
rect	33	105	34	106
rect	33	106	34	107
rect	33	107	34	108
rect	33	108	34	109
rect	33	109	34	110
rect	33	110	34	111
rect	33	111	34	112
rect	33	112	34	113
rect	33	113	34	114
rect	33	114	34	115
rect	33	115	34	116
rect	33	116	34	117
rect	33	118	34	119
rect	33	119	34	120
rect	33	120	34	121
rect	33	121	34	122
rect	33	122	34	123
rect	33	123	34	124
rect	33	125	34	126
rect	33	126	34	127
rect	33	127	34	128
rect	33	128	34	129
rect	33	129	34	130
rect	33	130	34	131
rect	33	131	34	132
rect	33	132	34	133
rect	33	133	34	134
rect	33	135	34	136
rect	33	136	34	137
rect	33	137	34	138
rect	33	138	34	139
rect	33	139	34	140
rect	33	140	34	141
rect	33	141	34	142
rect	33	142	34	143
rect	33	143	34	144
rect	34	0	35	1
rect	34	1	35	2
rect	34	2	35	3
rect	34	3	35	4
rect	34	4	35	5
rect	34	5	35	6
rect	34	6	35	7
rect	34	7	35	8
rect	34	8	35	9
rect	34	10	35	11
rect	34	11	35	12
rect	34	12	35	13
rect	34	13	35	14
rect	34	14	35	15
rect	34	15	35	16
rect	34	18	35	19
rect	34	21	35	22
rect	34	24	35	25
rect	34	27	35	28
rect	34	28	35	29
rect	34	29	35	30
rect	34	30	35	31
rect	34	31	35	32
rect	34	32	35	33
rect	34	33	35	34
rect	34	36	35	37
rect	34	37	35	38
rect	34	38	35	39
rect	34	39	35	40
rect	34	40	35	41
rect	34	41	35	42
rect	34	42	35	43
rect	34	43	35	44
rect	34	45	35	46
rect	34	46	35	47
rect	34	47	35	48
rect	34	48	35	49
rect	34	49	35	50
rect	34	50	35	51
rect	34	51	35	52
rect	34	52	35	53
rect	34	55	35	56
rect	34	56	35	57
rect	34	57	35	58
rect	34	60	35	61
rect	34	61	35	62
rect	34	62	35	63
rect	34	63	35	64
rect	34	64	35	65
rect	34	65	35	66
rect	34	67	35	68
rect	34	68	35	69
rect	34	69	35	70
rect	34	70	35	71
rect	34	71	35	72
rect	34	76	35	77
rect	34	77	35	78
rect	34	78	35	79
rect	34	79	35	80
rect	34	82	35	83
rect	34	86	35	87
rect	34	87	35	88
rect	34	88	35	89
rect	34	89	35	90
rect	34	90	35	91
rect	34	91	35	92
rect	34	92	35	93
rect	34	93	35	94
rect	34	94	35	95
rect	34	95	35	96
rect	34	96	35	97
rect	34	97	35	98
rect	34	98	35	99
rect	34	99	35	100
rect	34	100	35	101
rect	34	101	35	102
rect	34	102	35	103
rect	34	103	35	104
rect	34	105	35	106
rect	34	106	35	107
rect	34	107	35	108
rect	34	108	35	109
rect	34	109	35	110
rect	34	110	35	111
rect	34	111	35	112
rect	34	112	35	113
rect	34	113	35	114
rect	34	114	35	115
rect	34	115	35	116
rect	34	116	35	117
rect	34	118	35	119
rect	34	119	35	120
rect	34	120	35	121
rect	34	121	35	122
rect	34	122	35	123
rect	34	123	35	124
rect	34	125	35	126
rect	34	126	35	127
rect	34	127	35	128
rect	34	128	35	129
rect	34	129	35	130
rect	34	130	35	131
rect	34	131	35	132
rect	34	132	35	133
rect	34	133	35	134
rect	34	135	35	136
rect	34	136	35	137
rect	34	137	35	138
rect	34	138	35	139
rect	34	139	35	140
rect	34	140	35	141
rect	34	141	35	142
rect	34	142	35	143
rect	34	143	35	144
rect	35	0	36	1
rect	35	1	36	2
rect	35	2	36	3
rect	35	3	36	4
rect	35	4	36	5
rect	35	5	36	6
rect	35	6	36	7
rect	35	7	36	8
rect	35	8	36	9
rect	35	10	36	11
rect	35	11	36	12
rect	35	12	36	13
rect	35	13	36	14
rect	35	14	36	15
rect	35	15	36	16
rect	35	18	36	19
rect	35	21	36	22
rect	35	24	36	25
rect	35	27	36	28
rect	35	28	36	29
rect	35	29	36	30
rect	35	30	36	31
rect	35	31	36	32
rect	35	32	36	33
rect	35	33	36	34
rect	35	36	36	37
rect	35	37	36	38
rect	35	38	36	39
rect	35	39	36	40
rect	35	40	36	41
rect	35	41	36	42
rect	35	42	36	43
rect	35	43	36	44
rect	35	45	36	46
rect	35	46	36	47
rect	35	47	36	48
rect	35	48	36	49
rect	35	49	36	50
rect	35	50	36	51
rect	35	51	36	52
rect	35	52	36	53
rect	35	55	36	56
rect	35	56	36	57
rect	35	57	36	58
rect	35	60	36	61
rect	35	61	36	62
rect	35	62	36	63
rect	35	63	36	64
rect	35	64	36	65
rect	35	65	36	66
rect	35	67	36	68
rect	35	68	36	69
rect	35	69	36	70
rect	35	70	36	71
rect	35	71	36	72
rect	35	76	36	77
rect	35	77	36	78
rect	35	78	36	79
rect	35	79	36	80
rect	35	82	36	83
rect	35	86	36	87
rect	35	87	36	88
rect	35	88	36	89
rect	35	89	36	90
rect	35	90	36	91
rect	35	91	36	92
rect	35	92	36	93
rect	35	93	36	94
rect	35	94	36	95
rect	35	95	36	96
rect	35	96	36	97
rect	35	97	36	98
rect	35	98	36	99
rect	35	99	36	100
rect	35	100	36	101
rect	35	101	36	102
rect	35	102	36	103
rect	35	103	36	104
rect	35	105	36	106
rect	35	106	36	107
rect	35	107	36	108
rect	35	108	36	109
rect	35	109	36	110
rect	35	110	36	111
rect	35	111	36	112
rect	35	112	36	113
rect	35	113	36	114
rect	35	114	36	115
rect	35	115	36	116
rect	35	116	36	117
rect	35	118	36	119
rect	35	119	36	120
rect	35	120	36	121
rect	35	121	36	122
rect	35	122	36	123
rect	35	123	36	124
rect	35	125	36	126
rect	35	126	36	127
rect	35	127	36	128
rect	35	128	36	129
rect	35	129	36	130
rect	35	130	36	131
rect	35	131	36	132
rect	35	132	36	133
rect	35	133	36	134
rect	35	135	36	136
rect	35	136	36	137
rect	35	137	36	138
rect	35	138	36	139
rect	35	139	36	140
rect	35	140	36	141
rect	35	141	36	142
rect	35	142	36	143
rect	35	143	36	144
rect	36	0	37	1
rect	36	1	37	2
rect	36	2	37	3
rect	36	3	37	4
rect	36	4	37	5
rect	36	5	37	6
rect	36	6	37	7
rect	36	7	37	8
rect	36	8	37	9
rect	36	10	37	11
rect	36	11	37	12
rect	36	12	37	13
rect	36	13	37	14
rect	36	14	37	15
rect	36	15	37	16
rect	36	18	37	19
rect	36	21	37	22
rect	36	24	37	25
rect	36	27	37	28
rect	36	28	37	29
rect	36	29	37	30
rect	36	30	37	31
rect	36	31	37	32
rect	36	32	37	33
rect	36	33	37	34
rect	36	36	37	37
rect	36	37	37	38
rect	36	38	37	39
rect	36	39	37	40
rect	36	40	37	41
rect	36	41	37	42
rect	36	42	37	43
rect	36	43	37	44
rect	36	45	37	46
rect	36	46	37	47
rect	36	47	37	48
rect	36	48	37	49
rect	36	49	37	50
rect	36	50	37	51
rect	36	51	37	52
rect	36	52	37	53
rect	36	55	37	56
rect	36	56	37	57
rect	36	57	37	58
rect	36	60	37	61
rect	36	61	37	62
rect	36	62	37	63
rect	36	63	37	64
rect	36	64	37	65
rect	36	65	37	66
rect	36	67	37	68
rect	36	68	37	69
rect	36	69	37	70
rect	36	70	37	71
rect	36	71	37	72
rect	36	76	37	77
rect	36	77	37	78
rect	36	78	37	79
rect	36	79	37	80
rect	36	82	37	83
rect	36	86	37	87
rect	36	87	37	88
rect	36	88	37	89
rect	36	89	37	90
rect	36	90	37	91
rect	36	91	37	92
rect	36	92	37	93
rect	36	93	37	94
rect	36	94	37	95
rect	36	95	37	96
rect	36	96	37	97
rect	36	97	37	98
rect	36	98	37	99
rect	36	99	37	100
rect	36	100	37	101
rect	36	101	37	102
rect	36	102	37	103
rect	36	103	37	104
rect	36	105	37	106
rect	36	106	37	107
rect	36	107	37	108
rect	36	108	37	109
rect	36	109	37	110
rect	36	110	37	111
rect	36	111	37	112
rect	36	112	37	113
rect	36	113	37	114
rect	36	114	37	115
rect	36	115	37	116
rect	36	116	37	117
rect	36	118	37	119
rect	36	119	37	120
rect	36	120	37	121
rect	36	121	37	122
rect	36	122	37	123
rect	36	123	37	124
rect	36	125	37	126
rect	36	126	37	127
rect	36	127	37	128
rect	36	128	37	129
rect	36	129	37	130
rect	36	130	37	131
rect	36	131	37	132
rect	36	132	37	133
rect	36	133	37	134
rect	36	135	37	136
rect	36	136	37	137
rect	36	137	37	138
rect	36	138	37	139
rect	36	139	37	140
rect	36	140	37	141
rect	36	141	37	142
rect	36	142	37	143
rect	36	143	37	144
rect	56	0	57	1
rect	56	1	57	2
rect	56	2	57	3
rect	56	3	57	4
rect	56	4	57	5
rect	56	5	57	6
rect	56	6	57	7
rect	56	7	57	8
rect	56	8	57	9
rect	56	9	57	10
rect	56	10	57	11
rect	56	11	57	12
rect	56	12	57	13
rect	56	13	57	14
rect	56	14	57	15
rect	56	18	57	19
rect	56	21	57	22
rect	56	24	57	25
rect	56	27	57	28
rect	56	28	57	29
rect	56	29	57	30
rect	56	30	57	31
rect	56	32	57	33
rect	56	33	57	34
rect	56	36	57	37
rect	56	37	57	38
rect	56	38	57	39
rect	56	39	57	40
rect	56	40	57	41
rect	56	41	57	42
rect	56	42	57	43
rect	56	43	57	44
rect	56	44	57	45
rect	56	45	57	46
rect	56	46	57	47
rect	56	48	57	49
rect	56	49	57	50
rect	56	50	57	51
rect	56	51	57	52
rect	56	52	57	53
rect	56	55	57	56
rect	56	56	57	57
rect	56	57	57	58
rect	56	60	57	61
rect	56	61	57	62
rect	56	62	57	63
rect	56	63	57	64
rect	56	64	57	65
rect	56	65	57	66
rect	56	66	57	67
rect	56	67	57	68
rect	56	68	57	69
rect	56	69	57	70
rect	56	70	57	71
rect	56	71	57	72
rect	56	76	57	77
rect	56	77	57	78
rect	56	79	57	80
rect	56	82	57	83
rect	56	85	57	86
rect	56	86	57	87
rect	56	87	57	88
rect	56	88	57	89
rect	56	89	57	90
rect	56	90	57	91
rect	56	91	57	92
rect	56	92	57	93
rect	56	93	57	94
rect	56	95	57	96
rect	56	96	57	97
rect	56	97	57	98
rect	56	98	57	99
rect	56	99	57	100
rect	56	100	57	101
rect	56	101	57	102
rect	56	102	57	103
rect	56	103	57	104
rect	56	104	57	105
rect	56	105	57	106
rect	56	106	57	107
rect	56	107	57	108
rect	56	108	57	109
rect	56	109	57	110
rect	56	110	57	111
rect	56	111	57	112
rect	56	112	57	113
rect	56	114	57	115
rect	56	115	57	116
rect	56	116	57	117
rect	56	117	57	118
rect	56	118	57	119
rect	56	119	57	120
rect	56	120	57	121
rect	56	121	57	122
rect	56	122	57	123
rect	56	123	57	124
rect	56	124	57	125
rect	56	125	57	126
rect	56	127	57	128
rect	56	128	57	129
rect	56	129	57	130
rect	56	130	57	131
rect	56	131	57	132
rect	56	132	57	133
rect	56	133	57	134
rect	56	134	57	135
rect	56	135	57	136
rect	56	136	57	137
rect	56	137	57	138
rect	56	138	57	139
rect	56	140	57	141
rect	56	141	57	142
rect	56	142	57	143
rect	56	143	57	144
rect	56	144	57	145
rect	56	145	57	146
rect	56	146	57	147
rect	56	147	57	148
rect	56	148	57	149
rect	56	149	57	150
rect	56	150	57	151
rect	56	151	57	152
rect	56	153	57	154
rect	56	154	57	155
rect	56	155	57	156
rect	56	156	57	157
rect	56	157	57	158
rect	56	158	57	159
rect	56	159	57	160
rect	56	160	57	161
rect	56	161	57	162
rect	56	162	57	163
rect	56	163	57	164
rect	56	164	57	165
rect	56	165	57	166
rect	56	166	57	167
rect	56	167	57	168
rect	57	0	58	1
rect	57	1	58	2
rect	57	2	58	3
rect	57	3	58	4
rect	57	4	58	5
rect	57	5	58	6
rect	57	6	58	7
rect	57	7	58	8
rect	57	8	58	9
rect	57	9	58	10
rect	57	10	58	11
rect	57	11	58	12
rect	57	12	58	13
rect	57	13	58	14
rect	57	14	58	15
rect	57	18	58	19
rect	57	21	58	22
rect	57	24	58	25
rect	57	27	58	28
rect	57	28	58	29
rect	57	29	58	30
rect	57	30	58	31
rect	57	32	58	33
rect	57	33	58	34
rect	57	36	58	37
rect	57	37	58	38
rect	57	38	58	39
rect	57	39	58	40
rect	57	40	58	41
rect	57	41	58	42
rect	57	42	58	43
rect	57	43	58	44
rect	57	44	58	45
rect	57	45	58	46
rect	57	46	58	47
rect	57	48	58	49
rect	57	49	58	50
rect	57	50	58	51
rect	57	51	58	52
rect	57	52	58	53
rect	57	55	58	56
rect	57	56	58	57
rect	57	57	58	58
rect	57	60	58	61
rect	57	61	58	62
rect	57	62	58	63
rect	57	63	58	64
rect	57	64	58	65
rect	57	65	58	66
rect	57	66	58	67
rect	57	67	58	68
rect	57	68	58	69
rect	57	69	58	70
rect	57	70	58	71
rect	57	71	58	72
rect	57	76	58	77
rect	57	77	58	78
rect	57	79	58	80
rect	57	82	58	83
rect	57	85	58	86
rect	57	86	58	87
rect	57	87	58	88
rect	57	88	58	89
rect	57	89	58	90
rect	57	90	58	91
rect	57	91	58	92
rect	57	92	58	93
rect	57	93	58	94
rect	57	95	58	96
rect	57	96	58	97
rect	57	97	58	98
rect	57	98	58	99
rect	57	99	58	100
rect	57	100	58	101
rect	57	101	58	102
rect	57	102	58	103
rect	57	103	58	104
rect	57	104	58	105
rect	57	105	58	106
rect	57	106	58	107
rect	57	107	58	108
rect	57	108	58	109
rect	57	109	58	110
rect	57	110	58	111
rect	57	111	58	112
rect	57	112	58	113
rect	57	114	58	115
rect	57	115	58	116
rect	57	116	58	117
rect	57	117	58	118
rect	57	118	58	119
rect	57	119	58	120
rect	57	120	58	121
rect	57	121	58	122
rect	57	122	58	123
rect	57	123	58	124
rect	57	124	58	125
rect	57	125	58	126
rect	57	127	58	128
rect	57	128	58	129
rect	57	129	58	130
rect	57	130	58	131
rect	57	131	58	132
rect	57	132	58	133
rect	57	133	58	134
rect	57	134	58	135
rect	57	135	58	136
rect	57	136	58	137
rect	57	137	58	138
rect	57	138	58	139
rect	57	140	58	141
rect	57	141	58	142
rect	57	142	58	143
rect	57	143	58	144
rect	57	144	58	145
rect	57	145	58	146
rect	57	146	58	147
rect	57	147	58	148
rect	57	148	58	149
rect	57	149	58	150
rect	57	150	58	151
rect	57	151	58	152
rect	57	153	58	154
rect	57	154	58	155
rect	57	155	58	156
rect	57	156	58	157
rect	57	157	58	158
rect	57	158	58	159
rect	57	159	58	160
rect	57	160	58	161
rect	57	161	58	162
rect	57	162	58	163
rect	57	163	58	164
rect	57	164	58	165
rect	57	165	58	166
rect	57	166	58	167
rect	57	167	58	168
rect	58	0	59	1
rect	58	1	59	2
rect	58	2	59	3
rect	58	3	59	4
rect	58	4	59	5
rect	58	5	59	6
rect	58	6	59	7
rect	58	7	59	8
rect	58	8	59	9
rect	58	9	59	10
rect	58	10	59	11
rect	58	11	59	12
rect	58	12	59	13
rect	58	13	59	14
rect	58	14	59	15
rect	58	18	59	19
rect	58	21	59	22
rect	58	24	59	25
rect	58	27	59	28
rect	58	28	59	29
rect	58	29	59	30
rect	58	30	59	31
rect	58	32	59	33
rect	58	33	59	34
rect	58	36	59	37
rect	58	37	59	38
rect	58	38	59	39
rect	58	39	59	40
rect	58	40	59	41
rect	58	41	59	42
rect	58	42	59	43
rect	58	43	59	44
rect	58	44	59	45
rect	58	45	59	46
rect	58	46	59	47
rect	58	48	59	49
rect	58	49	59	50
rect	58	50	59	51
rect	58	51	59	52
rect	58	52	59	53
rect	58	55	59	56
rect	58	56	59	57
rect	58	57	59	58
rect	58	60	59	61
rect	58	61	59	62
rect	58	62	59	63
rect	58	63	59	64
rect	58	64	59	65
rect	58	65	59	66
rect	58	66	59	67
rect	58	67	59	68
rect	58	68	59	69
rect	58	69	59	70
rect	58	70	59	71
rect	58	71	59	72
rect	58	76	59	77
rect	58	77	59	78
rect	58	79	59	80
rect	58	82	59	83
rect	58	85	59	86
rect	58	86	59	87
rect	58	87	59	88
rect	58	88	59	89
rect	58	89	59	90
rect	58	90	59	91
rect	58	91	59	92
rect	58	92	59	93
rect	58	93	59	94
rect	58	95	59	96
rect	58	96	59	97
rect	58	97	59	98
rect	58	98	59	99
rect	58	99	59	100
rect	58	100	59	101
rect	58	101	59	102
rect	58	102	59	103
rect	58	103	59	104
rect	58	104	59	105
rect	58	105	59	106
rect	58	106	59	107
rect	58	107	59	108
rect	58	108	59	109
rect	58	109	59	110
rect	58	110	59	111
rect	58	111	59	112
rect	58	112	59	113
rect	58	114	59	115
rect	58	115	59	116
rect	58	116	59	117
rect	58	117	59	118
rect	58	118	59	119
rect	58	119	59	120
rect	58	120	59	121
rect	58	121	59	122
rect	58	122	59	123
rect	58	123	59	124
rect	58	124	59	125
rect	58	125	59	126
rect	58	127	59	128
rect	58	128	59	129
rect	58	129	59	130
rect	58	130	59	131
rect	58	131	59	132
rect	58	132	59	133
rect	58	133	59	134
rect	58	134	59	135
rect	58	135	59	136
rect	58	136	59	137
rect	58	137	59	138
rect	58	138	59	139
rect	58	140	59	141
rect	58	141	59	142
rect	58	142	59	143
rect	58	143	59	144
rect	58	144	59	145
rect	58	145	59	146
rect	58	146	59	147
rect	58	147	59	148
rect	58	148	59	149
rect	58	149	59	150
rect	58	150	59	151
rect	58	151	59	152
rect	58	153	59	154
rect	58	154	59	155
rect	58	155	59	156
rect	58	156	59	157
rect	58	157	59	158
rect	58	158	59	159
rect	58	159	59	160
rect	58	160	59	161
rect	58	161	59	162
rect	58	162	59	163
rect	58	163	59	164
rect	58	164	59	165
rect	58	165	59	166
rect	58	166	59	167
rect	58	167	59	168
rect	59	0	60	1
rect	59	1	60	2
rect	59	2	60	3
rect	59	3	60	4
rect	59	4	60	5
rect	59	5	60	6
rect	59	6	60	7
rect	59	7	60	8
rect	59	8	60	9
rect	59	9	60	10
rect	59	10	60	11
rect	59	11	60	12
rect	59	12	60	13
rect	59	13	60	14
rect	59	14	60	15
rect	59	18	60	19
rect	59	21	60	22
rect	59	24	60	25
rect	59	27	60	28
rect	59	28	60	29
rect	59	29	60	30
rect	59	30	60	31
rect	59	32	60	33
rect	59	33	60	34
rect	59	36	60	37
rect	59	37	60	38
rect	59	38	60	39
rect	59	39	60	40
rect	59	40	60	41
rect	59	41	60	42
rect	59	42	60	43
rect	59	43	60	44
rect	59	44	60	45
rect	59	45	60	46
rect	59	46	60	47
rect	59	48	60	49
rect	59	49	60	50
rect	59	50	60	51
rect	59	51	60	52
rect	59	52	60	53
rect	59	55	60	56
rect	59	56	60	57
rect	59	57	60	58
rect	59	60	60	61
rect	59	61	60	62
rect	59	62	60	63
rect	59	63	60	64
rect	59	64	60	65
rect	59	65	60	66
rect	59	66	60	67
rect	59	67	60	68
rect	59	68	60	69
rect	59	69	60	70
rect	59	70	60	71
rect	59	71	60	72
rect	59	76	60	77
rect	59	77	60	78
rect	59	79	60	80
rect	59	82	60	83
rect	59	85	60	86
rect	59	86	60	87
rect	59	87	60	88
rect	59	88	60	89
rect	59	89	60	90
rect	59	90	60	91
rect	59	91	60	92
rect	59	92	60	93
rect	59	93	60	94
rect	59	95	60	96
rect	59	96	60	97
rect	59	97	60	98
rect	59	98	60	99
rect	59	99	60	100
rect	59	100	60	101
rect	59	101	60	102
rect	59	102	60	103
rect	59	103	60	104
rect	59	104	60	105
rect	59	105	60	106
rect	59	106	60	107
rect	59	107	60	108
rect	59	108	60	109
rect	59	109	60	110
rect	59	110	60	111
rect	59	111	60	112
rect	59	112	60	113
rect	59	114	60	115
rect	59	115	60	116
rect	59	116	60	117
rect	59	117	60	118
rect	59	118	60	119
rect	59	119	60	120
rect	59	120	60	121
rect	59	121	60	122
rect	59	122	60	123
rect	59	123	60	124
rect	59	124	60	125
rect	59	125	60	126
rect	59	127	60	128
rect	59	128	60	129
rect	59	129	60	130
rect	59	130	60	131
rect	59	131	60	132
rect	59	132	60	133
rect	59	133	60	134
rect	59	134	60	135
rect	59	135	60	136
rect	59	136	60	137
rect	59	137	60	138
rect	59	138	60	139
rect	59	140	60	141
rect	59	141	60	142
rect	59	142	60	143
rect	59	143	60	144
rect	59	144	60	145
rect	59	145	60	146
rect	59	146	60	147
rect	59	147	60	148
rect	59	148	60	149
rect	59	149	60	150
rect	59	150	60	151
rect	59	151	60	152
rect	59	153	60	154
rect	59	154	60	155
rect	59	155	60	156
rect	59	156	60	157
rect	59	157	60	158
rect	59	158	60	159
rect	59	159	60	160
rect	59	160	60	161
rect	59	161	60	162
rect	59	162	60	163
rect	59	163	60	164
rect	59	164	60	165
rect	59	165	60	166
rect	59	166	60	167
rect	59	167	60	168
rect	60	0	61	1
rect	60	1	61	2
rect	60	2	61	3
rect	60	3	61	4
rect	60	4	61	5
rect	60	5	61	6
rect	60	6	61	7
rect	60	7	61	8
rect	60	8	61	9
rect	60	9	61	10
rect	60	10	61	11
rect	60	11	61	12
rect	60	12	61	13
rect	60	13	61	14
rect	60	14	61	15
rect	60	18	61	19
rect	60	21	61	22
rect	60	24	61	25
rect	60	27	61	28
rect	60	28	61	29
rect	60	29	61	30
rect	60	30	61	31
rect	60	32	61	33
rect	60	33	61	34
rect	60	36	61	37
rect	60	37	61	38
rect	60	38	61	39
rect	60	39	61	40
rect	60	40	61	41
rect	60	41	61	42
rect	60	42	61	43
rect	60	43	61	44
rect	60	44	61	45
rect	60	45	61	46
rect	60	46	61	47
rect	60	48	61	49
rect	60	49	61	50
rect	60	50	61	51
rect	60	51	61	52
rect	60	52	61	53
rect	60	55	61	56
rect	60	56	61	57
rect	60	57	61	58
rect	60	60	61	61
rect	60	61	61	62
rect	60	62	61	63
rect	60	63	61	64
rect	60	64	61	65
rect	60	65	61	66
rect	60	66	61	67
rect	60	67	61	68
rect	60	68	61	69
rect	60	69	61	70
rect	60	70	61	71
rect	60	71	61	72
rect	60	76	61	77
rect	60	77	61	78
rect	60	79	61	80
rect	60	82	61	83
rect	60	85	61	86
rect	60	86	61	87
rect	60	87	61	88
rect	60	88	61	89
rect	60	89	61	90
rect	60	90	61	91
rect	60	91	61	92
rect	60	92	61	93
rect	60	93	61	94
rect	60	95	61	96
rect	60	96	61	97
rect	60	97	61	98
rect	60	98	61	99
rect	60	99	61	100
rect	60	100	61	101
rect	60	101	61	102
rect	60	102	61	103
rect	60	103	61	104
rect	60	104	61	105
rect	60	105	61	106
rect	60	106	61	107
rect	60	107	61	108
rect	60	108	61	109
rect	60	109	61	110
rect	60	110	61	111
rect	60	111	61	112
rect	60	112	61	113
rect	60	114	61	115
rect	60	115	61	116
rect	60	116	61	117
rect	60	117	61	118
rect	60	118	61	119
rect	60	119	61	120
rect	60	120	61	121
rect	60	121	61	122
rect	60	122	61	123
rect	60	123	61	124
rect	60	124	61	125
rect	60	125	61	126
rect	60	127	61	128
rect	60	128	61	129
rect	60	129	61	130
rect	60	130	61	131
rect	60	131	61	132
rect	60	132	61	133
rect	60	133	61	134
rect	60	134	61	135
rect	60	135	61	136
rect	60	136	61	137
rect	60	137	61	138
rect	60	138	61	139
rect	60	140	61	141
rect	60	141	61	142
rect	60	142	61	143
rect	60	143	61	144
rect	60	144	61	145
rect	60	145	61	146
rect	60	146	61	147
rect	60	147	61	148
rect	60	148	61	149
rect	60	149	61	150
rect	60	150	61	151
rect	60	151	61	152
rect	60	153	61	154
rect	60	154	61	155
rect	60	155	61	156
rect	60	156	61	157
rect	60	157	61	158
rect	60	158	61	159
rect	60	159	61	160
rect	60	160	61	161
rect	60	161	61	162
rect	60	162	61	163
rect	60	163	61	164
rect	60	164	61	165
rect	60	165	61	166
rect	60	166	61	167
rect	60	167	61	168
rect	61	0	62	1
rect	61	1	62	2
rect	61	2	62	3
rect	61	3	62	4
rect	61	4	62	5
rect	61	5	62	6
rect	61	6	62	7
rect	61	7	62	8
rect	61	8	62	9
rect	61	9	62	10
rect	61	10	62	11
rect	61	11	62	12
rect	61	12	62	13
rect	61	13	62	14
rect	61	14	62	15
rect	61	18	62	19
rect	61	21	62	22
rect	61	24	62	25
rect	61	27	62	28
rect	61	28	62	29
rect	61	29	62	30
rect	61	30	62	31
rect	61	32	62	33
rect	61	33	62	34
rect	61	36	62	37
rect	61	37	62	38
rect	61	38	62	39
rect	61	39	62	40
rect	61	40	62	41
rect	61	41	62	42
rect	61	42	62	43
rect	61	43	62	44
rect	61	44	62	45
rect	61	45	62	46
rect	61	46	62	47
rect	61	48	62	49
rect	61	49	62	50
rect	61	50	62	51
rect	61	51	62	52
rect	61	52	62	53
rect	61	55	62	56
rect	61	56	62	57
rect	61	57	62	58
rect	61	60	62	61
rect	61	61	62	62
rect	61	62	62	63
rect	61	63	62	64
rect	61	64	62	65
rect	61	65	62	66
rect	61	66	62	67
rect	61	67	62	68
rect	61	68	62	69
rect	61	69	62	70
rect	61	70	62	71
rect	61	71	62	72
rect	61	76	62	77
rect	61	77	62	78
rect	61	79	62	80
rect	61	82	62	83
rect	61	85	62	86
rect	61	86	62	87
rect	61	87	62	88
rect	61	88	62	89
rect	61	89	62	90
rect	61	90	62	91
rect	61	91	62	92
rect	61	92	62	93
rect	61	93	62	94
rect	61	95	62	96
rect	61	96	62	97
rect	61	97	62	98
rect	61	98	62	99
rect	61	99	62	100
rect	61	100	62	101
rect	61	101	62	102
rect	61	102	62	103
rect	61	103	62	104
rect	61	104	62	105
rect	61	105	62	106
rect	61	106	62	107
rect	61	107	62	108
rect	61	108	62	109
rect	61	109	62	110
rect	61	110	62	111
rect	61	111	62	112
rect	61	112	62	113
rect	61	114	62	115
rect	61	115	62	116
rect	61	116	62	117
rect	61	117	62	118
rect	61	118	62	119
rect	61	119	62	120
rect	61	120	62	121
rect	61	121	62	122
rect	61	122	62	123
rect	61	123	62	124
rect	61	124	62	125
rect	61	125	62	126
rect	61	127	62	128
rect	61	128	62	129
rect	61	129	62	130
rect	61	130	62	131
rect	61	131	62	132
rect	61	132	62	133
rect	61	133	62	134
rect	61	134	62	135
rect	61	135	62	136
rect	61	136	62	137
rect	61	137	62	138
rect	61	138	62	139
rect	61	140	62	141
rect	61	141	62	142
rect	61	142	62	143
rect	61	143	62	144
rect	61	144	62	145
rect	61	145	62	146
rect	61	146	62	147
rect	61	147	62	148
rect	61	148	62	149
rect	61	149	62	150
rect	61	150	62	151
rect	61	151	62	152
rect	61	153	62	154
rect	61	154	62	155
rect	61	155	62	156
rect	61	156	62	157
rect	61	157	62	158
rect	61	158	62	159
rect	61	159	62	160
rect	61	160	62	161
rect	61	161	62	162
rect	61	162	62	163
rect	61	163	62	164
rect	61	164	62	165
rect	61	165	62	166
rect	61	166	62	167
rect	61	167	62	168
rect	89	0	90	1
rect	89	1	90	2
rect	89	2	90	3
rect	89	3	90	4
rect	89	4	90	5
rect	89	5	90	6
rect	89	7	90	8
rect	89	8	90	9
rect	89	9	90	10
rect	89	10	90	11
rect	89	11	90	12
rect	89	12	90	13
rect	89	13	90	14
rect	89	14	90	15
rect	89	15	90	16
rect	89	18	90	19
rect	89	21	90	22
rect	89	24	90	25
rect	89	27	90	28
rect	89	28	90	29
rect	89	29	90	30
rect	89	30	90	31
rect	89	32	90	33
rect	89	33	90	34
rect	89	36	90	37
rect	89	37	90	38
rect	89	38	90	39
rect	89	39	90	40
rect	89	40	90	41
rect	89	41	90	42
rect	89	42	90	43
rect	89	43	90	44
rect	89	45	90	46
rect	89	46	90	47
rect	89	47	90	48
rect	89	48	90	49
rect	89	49	90	50
rect	89	50	90	51
rect	89	51	90	52
rect	89	52	90	53
rect	89	55	90	56
rect	89	56	90	57
rect	89	57	90	58
rect	89	60	90	61
rect	89	61	90	62
rect	89	62	90	63
rect	89	63	90	64
rect	89	64	90	65
rect	89	65	90	66
rect	89	66	90	67
rect	89	67	90	68
rect	89	68	90	69
rect	89	69	90	70
rect	89	70	90	71
rect	89	71	90	72
rect	89	76	90	77
rect	89	77	90	78
rect	89	78	90	79
rect	89	79	90	80
rect	89	82	90	83
rect	89	86	90	87
rect	89	87	90	88
rect	89	88	90	89
rect	89	89	90	90
rect	89	90	90	91
rect	89	91	90	92
rect	89	92	90	93
rect	89	93	90	94
rect	89	94	90	95
rect	89	96	90	97
rect	89	97	90	98
rect	89	98	90	99
rect	89	99	90	100
rect	89	100	90	101
rect	89	101	90	102
rect	89	102	90	103
rect	89	103	90	104
rect	89	104	90	105
rect	89	105	90	106
rect	89	106	90	107
rect	89	107	90	108
rect	89	108	90	109
rect	89	109	90	110
rect	89	110	90	111
rect	89	111	90	112
rect	89	112	90	113
rect	89	113	90	114
rect	89	114	90	115
rect	89	115	90	116
rect	89	116	90	117
rect	89	118	90	119
rect	89	119	90	120
rect	89	120	90	121
rect	89	121	90	122
rect	89	122	90	123
rect	89	123	90	124
rect	89	124	90	125
rect	89	125	90	126
rect	89	126	90	127
rect	89	127	90	128
rect	89	128	90	129
rect	89	129	90	130
rect	89	130	90	131
rect	89	131	90	132
rect	89	132	90	133
rect	89	133	90	134
rect	89	134	90	135
rect	89	135	90	136
rect	89	136	90	137
rect	89	137	90	138
rect	89	138	90	139
rect	89	139	90	140
rect	89	140	90	141
rect	89	141	90	142
rect	89	143	90	144
rect	89	144	90	145
rect	89	145	90	146
rect	89	146	90	147
rect	89	147	90	148
rect	89	148	90	149
rect	89	149	90	150
rect	89	150	90	151
rect	89	151	90	152
rect	89	152	90	153
rect	89	153	90	154
rect	89	154	90	155
rect	89	155	90	156
rect	89	156	90	157
rect	89	157	90	158
rect	89	159	90	160
rect	89	160	90	161
rect	89	161	90	162
rect	89	162	90	163
rect	89	163	90	164
rect	89	164	90	165
rect	89	165	90	166
rect	89	166	90	167
rect	89	167	90	168
rect	89	168	90	169
rect	89	169	90	170
rect	89	170	90	171
rect	89	171	90	172
rect	89	172	90	173
rect	89	173	90	174
rect	89	174	90	175
rect	89	175	90	176
rect	89	176	90	177
rect	89	177	90	178
rect	89	178	90	179
rect	89	179	90	180
rect	89	207	90	208
rect	89	208	90	209
rect	89	209	90	210
rect	90	0	91	1
rect	90	1	91	2
rect	90	2	91	3
rect	90	3	91	4
rect	90	4	91	5
rect	90	5	91	6
rect	90	7	91	8
rect	90	8	91	9
rect	90	9	91	10
rect	90	10	91	11
rect	90	11	91	12
rect	90	12	91	13
rect	90	13	91	14
rect	90	14	91	15
rect	90	15	91	16
rect	90	18	91	19
rect	90	21	91	22
rect	90	24	91	25
rect	90	27	91	28
rect	90	28	91	29
rect	90	29	91	30
rect	90	30	91	31
rect	90	32	91	33
rect	90	33	91	34
rect	90	36	91	37
rect	90	37	91	38
rect	90	38	91	39
rect	90	39	91	40
rect	90	40	91	41
rect	90	41	91	42
rect	90	42	91	43
rect	90	43	91	44
rect	90	45	91	46
rect	90	46	91	47
rect	90	47	91	48
rect	90	48	91	49
rect	90	49	91	50
rect	90	50	91	51
rect	90	51	91	52
rect	90	52	91	53
rect	90	55	91	56
rect	90	56	91	57
rect	90	57	91	58
rect	90	60	91	61
rect	90	61	91	62
rect	90	62	91	63
rect	90	63	91	64
rect	90	64	91	65
rect	90	65	91	66
rect	90	66	91	67
rect	90	67	91	68
rect	90	68	91	69
rect	90	69	91	70
rect	90	70	91	71
rect	90	71	91	72
rect	90	76	91	77
rect	90	77	91	78
rect	90	78	91	79
rect	90	79	91	80
rect	90	82	91	83
rect	90	86	91	87
rect	90	87	91	88
rect	90	88	91	89
rect	90	89	91	90
rect	90	90	91	91
rect	90	91	91	92
rect	90	92	91	93
rect	90	93	91	94
rect	90	94	91	95
rect	90	96	91	97
rect	90	97	91	98
rect	90	98	91	99
rect	90	99	91	100
rect	90	100	91	101
rect	90	101	91	102
rect	90	102	91	103
rect	90	103	91	104
rect	90	104	91	105
rect	90	105	91	106
rect	90	106	91	107
rect	90	107	91	108
rect	90	108	91	109
rect	90	109	91	110
rect	90	110	91	111
rect	90	111	91	112
rect	90	112	91	113
rect	90	113	91	114
rect	90	114	91	115
rect	90	115	91	116
rect	90	116	91	117
rect	90	118	91	119
rect	90	119	91	120
rect	90	120	91	121
rect	90	121	91	122
rect	90	122	91	123
rect	90	123	91	124
rect	90	124	91	125
rect	90	125	91	126
rect	90	126	91	127
rect	90	127	91	128
rect	90	128	91	129
rect	90	129	91	130
rect	90	130	91	131
rect	90	131	91	132
rect	90	132	91	133
rect	90	133	91	134
rect	90	134	91	135
rect	90	135	91	136
rect	90	136	91	137
rect	90	137	91	138
rect	90	138	91	139
rect	90	139	91	140
rect	90	140	91	141
rect	90	141	91	142
rect	90	143	91	144
rect	90	144	91	145
rect	90	145	91	146
rect	90	146	91	147
rect	90	147	91	148
rect	90	148	91	149
rect	90	149	91	150
rect	90	150	91	151
rect	90	151	91	152
rect	90	152	91	153
rect	90	153	91	154
rect	90	154	91	155
rect	90	155	91	156
rect	90	156	91	157
rect	90	157	91	158
rect	90	159	91	160
rect	90	160	91	161
rect	90	161	91	162
rect	90	162	91	163
rect	90	163	91	164
rect	90	164	91	165
rect	90	165	91	166
rect	90	166	91	167
rect	90	167	91	168
rect	90	168	91	169
rect	90	169	91	170
rect	90	170	91	171
rect	90	171	91	172
rect	90	172	91	173
rect	90	173	91	174
rect	90	174	91	175
rect	90	175	91	176
rect	90	176	91	177
rect	90	177	91	178
rect	90	178	91	179
rect	90	179	91	180
rect	90	207	91	208
rect	90	208	91	209
rect	90	209	91	210
rect	91	0	92	1
rect	91	1	92	2
rect	91	2	92	3
rect	91	3	92	4
rect	91	4	92	5
rect	91	5	92	6
rect	91	7	92	8
rect	91	8	92	9
rect	91	9	92	10
rect	91	10	92	11
rect	91	11	92	12
rect	91	12	92	13
rect	91	13	92	14
rect	91	14	92	15
rect	91	15	92	16
rect	91	18	92	19
rect	91	21	92	22
rect	91	24	92	25
rect	91	27	92	28
rect	91	28	92	29
rect	91	29	92	30
rect	91	30	92	31
rect	91	32	92	33
rect	91	33	92	34
rect	91	36	92	37
rect	91	37	92	38
rect	91	38	92	39
rect	91	39	92	40
rect	91	40	92	41
rect	91	41	92	42
rect	91	42	92	43
rect	91	43	92	44
rect	91	45	92	46
rect	91	46	92	47
rect	91	47	92	48
rect	91	48	92	49
rect	91	49	92	50
rect	91	50	92	51
rect	91	51	92	52
rect	91	52	92	53
rect	91	55	92	56
rect	91	56	92	57
rect	91	57	92	58
rect	91	60	92	61
rect	91	61	92	62
rect	91	62	92	63
rect	91	63	92	64
rect	91	64	92	65
rect	91	65	92	66
rect	91	66	92	67
rect	91	67	92	68
rect	91	68	92	69
rect	91	69	92	70
rect	91	70	92	71
rect	91	71	92	72
rect	91	76	92	77
rect	91	77	92	78
rect	91	78	92	79
rect	91	79	92	80
rect	91	82	92	83
rect	91	86	92	87
rect	91	87	92	88
rect	91	88	92	89
rect	91	89	92	90
rect	91	90	92	91
rect	91	91	92	92
rect	91	92	92	93
rect	91	93	92	94
rect	91	94	92	95
rect	91	96	92	97
rect	91	97	92	98
rect	91	98	92	99
rect	91	99	92	100
rect	91	100	92	101
rect	91	101	92	102
rect	91	102	92	103
rect	91	103	92	104
rect	91	104	92	105
rect	91	105	92	106
rect	91	106	92	107
rect	91	107	92	108
rect	91	108	92	109
rect	91	109	92	110
rect	91	110	92	111
rect	91	111	92	112
rect	91	112	92	113
rect	91	113	92	114
rect	91	114	92	115
rect	91	115	92	116
rect	91	116	92	117
rect	91	118	92	119
rect	91	119	92	120
rect	91	120	92	121
rect	91	121	92	122
rect	91	122	92	123
rect	91	123	92	124
rect	91	124	92	125
rect	91	125	92	126
rect	91	126	92	127
rect	91	127	92	128
rect	91	128	92	129
rect	91	129	92	130
rect	91	130	92	131
rect	91	131	92	132
rect	91	132	92	133
rect	91	133	92	134
rect	91	134	92	135
rect	91	135	92	136
rect	91	136	92	137
rect	91	137	92	138
rect	91	138	92	139
rect	91	139	92	140
rect	91	140	92	141
rect	91	141	92	142
rect	91	143	92	144
rect	91	144	92	145
rect	91	145	92	146
rect	91	146	92	147
rect	91	147	92	148
rect	91	148	92	149
rect	91	149	92	150
rect	91	150	92	151
rect	91	151	92	152
rect	91	152	92	153
rect	91	153	92	154
rect	91	154	92	155
rect	91	155	92	156
rect	91	156	92	157
rect	91	157	92	158
rect	91	159	92	160
rect	91	160	92	161
rect	91	161	92	162
rect	91	162	92	163
rect	91	163	92	164
rect	91	164	92	165
rect	91	165	92	166
rect	91	166	92	167
rect	91	167	92	168
rect	91	168	92	169
rect	91	169	92	170
rect	91	170	92	171
rect	91	171	92	172
rect	91	172	92	173
rect	91	173	92	174
rect	91	174	92	175
rect	91	175	92	176
rect	91	176	92	177
rect	91	177	92	178
rect	91	178	92	179
rect	91	179	92	180
rect	91	207	92	208
rect	91	208	92	209
rect	91	209	92	210
rect	92	0	93	1
rect	92	1	93	2
rect	92	2	93	3
rect	92	3	93	4
rect	92	4	93	5
rect	92	5	93	6
rect	92	7	93	8
rect	92	8	93	9
rect	92	9	93	10
rect	92	10	93	11
rect	92	11	93	12
rect	92	12	93	13
rect	92	13	93	14
rect	92	14	93	15
rect	92	15	93	16
rect	92	18	93	19
rect	92	21	93	22
rect	92	24	93	25
rect	92	27	93	28
rect	92	28	93	29
rect	92	29	93	30
rect	92	30	93	31
rect	92	32	93	33
rect	92	33	93	34
rect	92	36	93	37
rect	92	37	93	38
rect	92	38	93	39
rect	92	39	93	40
rect	92	40	93	41
rect	92	41	93	42
rect	92	42	93	43
rect	92	43	93	44
rect	92	45	93	46
rect	92	46	93	47
rect	92	47	93	48
rect	92	48	93	49
rect	92	49	93	50
rect	92	50	93	51
rect	92	51	93	52
rect	92	52	93	53
rect	92	55	93	56
rect	92	56	93	57
rect	92	57	93	58
rect	92	60	93	61
rect	92	61	93	62
rect	92	62	93	63
rect	92	63	93	64
rect	92	64	93	65
rect	92	65	93	66
rect	92	66	93	67
rect	92	67	93	68
rect	92	68	93	69
rect	92	69	93	70
rect	92	70	93	71
rect	92	71	93	72
rect	92	76	93	77
rect	92	77	93	78
rect	92	78	93	79
rect	92	79	93	80
rect	92	82	93	83
rect	92	86	93	87
rect	92	87	93	88
rect	92	88	93	89
rect	92	89	93	90
rect	92	90	93	91
rect	92	91	93	92
rect	92	92	93	93
rect	92	93	93	94
rect	92	94	93	95
rect	92	96	93	97
rect	92	97	93	98
rect	92	98	93	99
rect	92	99	93	100
rect	92	100	93	101
rect	92	101	93	102
rect	92	102	93	103
rect	92	103	93	104
rect	92	104	93	105
rect	92	105	93	106
rect	92	106	93	107
rect	92	107	93	108
rect	92	108	93	109
rect	92	109	93	110
rect	92	110	93	111
rect	92	111	93	112
rect	92	112	93	113
rect	92	113	93	114
rect	92	114	93	115
rect	92	115	93	116
rect	92	116	93	117
rect	92	118	93	119
rect	92	119	93	120
rect	92	120	93	121
rect	92	121	93	122
rect	92	122	93	123
rect	92	123	93	124
rect	92	124	93	125
rect	92	125	93	126
rect	92	126	93	127
rect	92	127	93	128
rect	92	128	93	129
rect	92	129	93	130
rect	92	130	93	131
rect	92	131	93	132
rect	92	132	93	133
rect	92	133	93	134
rect	92	134	93	135
rect	92	135	93	136
rect	92	136	93	137
rect	92	137	93	138
rect	92	138	93	139
rect	92	139	93	140
rect	92	140	93	141
rect	92	141	93	142
rect	92	143	93	144
rect	92	144	93	145
rect	92	145	93	146
rect	92	146	93	147
rect	92	147	93	148
rect	92	148	93	149
rect	92	149	93	150
rect	92	150	93	151
rect	92	151	93	152
rect	92	152	93	153
rect	92	153	93	154
rect	92	154	93	155
rect	92	155	93	156
rect	92	156	93	157
rect	92	157	93	158
rect	92	159	93	160
rect	92	160	93	161
rect	92	161	93	162
rect	92	162	93	163
rect	92	163	93	164
rect	92	164	93	165
rect	92	165	93	166
rect	92	166	93	167
rect	92	167	93	168
rect	92	168	93	169
rect	92	169	93	170
rect	92	170	93	171
rect	92	171	93	172
rect	92	172	93	173
rect	92	173	93	174
rect	92	174	93	175
rect	92	175	93	176
rect	92	176	93	177
rect	92	177	93	178
rect	92	178	93	179
rect	92	179	93	180
rect	92	207	93	208
rect	92	208	93	209
rect	92	209	93	210
rect	93	0	94	1
rect	93	1	94	2
rect	93	2	94	3
rect	93	3	94	4
rect	93	4	94	5
rect	93	5	94	6
rect	93	7	94	8
rect	93	8	94	9
rect	93	9	94	10
rect	93	10	94	11
rect	93	11	94	12
rect	93	12	94	13
rect	93	13	94	14
rect	93	14	94	15
rect	93	15	94	16
rect	93	18	94	19
rect	93	21	94	22
rect	93	24	94	25
rect	93	27	94	28
rect	93	28	94	29
rect	93	29	94	30
rect	93	30	94	31
rect	93	32	94	33
rect	93	33	94	34
rect	93	36	94	37
rect	93	37	94	38
rect	93	38	94	39
rect	93	39	94	40
rect	93	40	94	41
rect	93	41	94	42
rect	93	42	94	43
rect	93	43	94	44
rect	93	45	94	46
rect	93	46	94	47
rect	93	47	94	48
rect	93	48	94	49
rect	93	49	94	50
rect	93	50	94	51
rect	93	51	94	52
rect	93	52	94	53
rect	93	55	94	56
rect	93	56	94	57
rect	93	57	94	58
rect	93	60	94	61
rect	93	61	94	62
rect	93	62	94	63
rect	93	63	94	64
rect	93	64	94	65
rect	93	65	94	66
rect	93	66	94	67
rect	93	67	94	68
rect	93	68	94	69
rect	93	69	94	70
rect	93	70	94	71
rect	93	71	94	72
rect	93	76	94	77
rect	93	77	94	78
rect	93	78	94	79
rect	93	79	94	80
rect	93	82	94	83
rect	93	86	94	87
rect	93	87	94	88
rect	93	88	94	89
rect	93	89	94	90
rect	93	90	94	91
rect	93	91	94	92
rect	93	92	94	93
rect	93	93	94	94
rect	93	94	94	95
rect	93	96	94	97
rect	93	97	94	98
rect	93	98	94	99
rect	93	99	94	100
rect	93	100	94	101
rect	93	101	94	102
rect	93	102	94	103
rect	93	103	94	104
rect	93	104	94	105
rect	93	105	94	106
rect	93	106	94	107
rect	93	107	94	108
rect	93	108	94	109
rect	93	109	94	110
rect	93	110	94	111
rect	93	111	94	112
rect	93	112	94	113
rect	93	113	94	114
rect	93	114	94	115
rect	93	115	94	116
rect	93	116	94	117
rect	93	118	94	119
rect	93	119	94	120
rect	93	120	94	121
rect	93	121	94	122
rect	93	122	94	123
rect	93	123	94	124
rect	93	124	94	125
rect	93	125	94	126
rect	93	126	94	127
rect	93	127	94	128
rect	93	128	94	129
rect	93	129	94	130
rect	93	130	94	131
rect	93	131	94	132
rect	93	132	94	133
rect	93	133	94	134
rect	93	134	94	135
rect	93	135	94	136
rect	93	136	94	137
rect	93	137	94	138
rect	93	138	94	139
rect	93	139	94	140
rect	93	140	94	141
rect	93	141	94	142
rect	93	143	94	144
rect	93	144	94	145
rect	93	145	94	146
rect	93	146	94	147
rect	93	147	94	148
rect	93	148	94	149
rect	93	149	94	150
rect	93	150	94	151
rect	93	151	94	152
rect	93	152	94	153
rect	93	153	94	154
rect	93	154	94	155
rect	93	155	94	156
rect	93	156	94	157
rect	93	157	94	158
rect	93	159	94	160
rect	93	160	94	161
rect	93	161	94	162
rect	93	162	94	163
rect	93	163	94	164
rect	93	164	94	165
rect	93	165	94	166
rect	93	166	94	167
rect	93	167	94	168
rect	93	168	94	169
rect	93	169	94	170
rect	93	170	94	171
rect	93	171	94	172
rect	93	172	94	173
rect	93	173	94	174
rect	93	174	94	175
rect	93	175	94	176
rect	93	176	94	177
rect	93	177	94	178
rect	93	178	94	179
rect	93	179	94	180
rect	93	207	94	208
rect	93	208	94	209
rect	93	209	94	210
rect	94	0	95	1
rect	94	1	95	2
rect	94	2	95	3
rect	94	3	95	4
rect	94	4	95	5
rect	94	5	95	6
rect	94	7	95	8
rect	94	8	95	9
rect	94	9	95	10
rect	94	10	95	11
rect	94	11	95	12
rect	94	12	95	13
rect	94	13	95	14
rect	94	14	95	15
rect	94	15	95	16
rect	94	18	95	19
rect	94	21	95	22
rect	94	24	95	25
rect	94	27	95	28
rect	94	28	95	29
rect	94	29	95	30
rect	94	30	95	31
rect	94	32	95	33
rect	94	33	95	34
rect	94	36	95	37
rect	94	37	95	38
rect	94	38	95	39
rect	94	39	95	40
rect	94	40	95	41
rect	94	41	95	42
rect	94	42	95	43
rect	94	43	95	44
rect	94	45	95	46
rect	94	46	95	47
rect	94	47	95	48
rect	94	48	95	49
rect	94	49	95	50
rect	94	50	95	51
rect	94	51	95	52
rect	94	52	95	53
rect	94	55	95	56
rect	94	56	95	57
rect	94	57	95	58
rect	94	60	95	61
rect	94	61	95	62
rect	94	62	95	63
rect	94	63	95	64
rect	94	64	95	65
rect	94	65	95	66
rect	94	66	95	67
rect	94	67	95	68
rect	94	68	95	69
rect	94	69	95	70
rect	94	70	95	71
rect	94	71	95	72
rect	94	74	95	75
rect	94	76	95	77
rect	94	77	95	78
rect	94	78	95	79
rect	94	79	95	80
rect	94	80	95	81
rect	94	82	95	83
rect	94	86	95	87
rect	94	87	95	88
rect	94	88	95	89
rect	94	89	95	90
rect	94	90	95	91
rect	94	91	95	92
rect	94	92	95	93
rect	94	93	95	94
rect	94	94	95	95
rect	94	96	95	97
rect	94	97	95	98
rect	94	98	95	99
rect	94	99	95	100
rect	94	100	95	101
rect	94	101	95	102
rect	94	102	95	103
rect	94	103	95	104
rect	94	104	95	105
rect	94	105	95	106
rect	94	106	95	107
rect	94	107	95	108
rect	94	108	95	109
rect	94	109	95	110
rect	94	110	95	111
rect	94	111	95	112
rect	94	112	95	113
rect	94	113	95	114
rect	94	114	95	115
rect	94	115	95	116
rect	94	116	95	117
rect	94	118	95	119
rect	94	119	95	120
rect	94	120	95	121
rect	94	121	95	122
rect	94	122	95	123
rect	94	123	95	124
rect	94	124	95	125
rect	94	125	95	126
rect	94	126	95	127
rect	94	127	95	128
rect	94	128	95	129
rect	94	129	95	130
rect	94	130	95	131
rect	94	131	95	132
rect	94	132	95	133
rect	94	133	95	134
rect	94	134	95	135
rect	94	135	95	136
rect	94	136	95	137
rect	94	137	95	138
rect	94	138	95	139
rect	94	139	95	140
rect	94	140	95	141
rect	94	141	95	142
rect	94	143	95	144
rect	94	144	95	145
rect	94	145	95	146
rect	94	146	95	147
rect	94	147	95	148
rect	94	148	95	149
rect	94	149	95	150
rect	94	150	95	151
rect	94	151	95	152
rect	94	152	95	153
rect	94	153	95	154
rect	94	154	95	155
rect	94	155	95	156
rect	94	156	95	157
rect	94	157	95	158
rect	94	159	95	160
rect	94	160	95	161
rect	94	161	95	162
rect	94	162	95	163
rect	94	163	95	164
rect	94	164	95	165
rect	94	165	95	166
rect	94	166	95	167
rect	94	167	95	168
rect	94	168	95	169
rect	94	169	95	170
rect	94	170	95	171
rect	94	171	95	172
rect	94	172	95	173
rect	94	173	95	174
rect	94	174	95	175
rect	94	175	95	176
rect	94	176	95	177
rect	94	177	95	178
rect	94	178	95	179
rect	94	179	95	180
rect	94	207	95	208
rect	94	208	95	209
rect	94	209	95	210
rect	126	0	127	1
rect	126	1	127	2
rect	126	2	127	3
rect	126	3	127	4
rect	126	4	127	5
rect	126	5	127	6
rect	126	6	127	7
rect	126	7	127	8
rect	126	8	127	9
rect	126	9	127	10
rect	126	10	127	11
rect	126	11	127	12
rect	126	12	127	13
rect	126	13	127	14
rect	126	14	127	15
rect	126	15	127	16
rect	126	18	127	19
rect	126	21	127	22
rect	126	24	127	25
rect	126	27	127	28
rect	126	28	127	29
rect	126	29	127	30
rect	126	30	127	31
rect	126	31	127	32
rect	126	32	127	33
rect	126	33	127	34
rect	126	37	127	38
rect	126	38	127	39
rect	126	39	127	40
rect	126	40	127	41
rect	126	41	127	42
rect	126	42	127	43
rect	126	43	127	44
rect	126	44	127	45
rect	126	45	127	46
rect	126	46	127	47
rect	126	47	127	48
rect	126	48	127	49
rect	126	50	127	51
rect	126	51	127	52
rect	126	52	127	53
rect	126	55	127	56
rect	126	56	127	57
rect	126	57	127	58
rect	126	60	127	61
rect	126	61	127	62
rect	126	62	127	63
rect	126	63	127	64
rect	126	64	127	65
rect	126	65	127	66
rect	126	66	127	67
rect	126	67	127	68
rect	126	68	127	69
rect	126	69	127	70
rect	126	70	127	71
rect	126	71	127	72
rect	126	74	127	75
rect	126	75	127	76
rect	126	76	127	77
rect	126	77	127	78
rect	126	78	127	79
rect	126	79	127	80
rect	126	80	127	81
rect	126	81	127	82
rect	126	82	127	83
rect	126	85	127	86
rect	126	87	127	88
rect	126	88	127	89
rect	126	89	127	90
rect	126	90	127	91
rect	126	91	127	92
rect	126	92	127	93
rect	126	93	127	94
rect	126	94	127	95
rect	126	95	127	96
rect	126	96	127	97
rect	126	97	127	98
rect	126	98	127	99
rect	126	99	127	100
rect	126	100	127	101
rect	126	101	127	102
rect	126	103	127	104
rect	126	104	127	105
rect	126	105	127	106
rect	126	106	127	107
rect	126	107	127	108
rect	126	108	127	109
rect	126	109	127	110
rect	126	110	127	111
rect	126	111	127	112
rect	126	112	127	113
rect	126	113	127	114
rect	126	114	127	115
rect	126	115	127	116
rect	126	116	127	117
rect	126	117	127	118
rect	126	119	127	120
rect	126	120	127	121
rect	126	121	127	122
rect	126	122	127	123
rect	126	123	127	124
rect	126	124	127	125
rect	126	125	127	126
rect	126	126	127	127
rect	126	127	127	128
rect	126	128	127	129
rect	126	129	127	130
rect	126	130	127	131
rect	126	131	127	132
rect	126	132	127	133
rect	126	133	127	134
rect	126	134	127	135
rect	126	135	127	136
rect	126	136	127	137
rect	126	137	127	138
rect	126	138	127	139
rect	126	139	127	140
rect	126	141	127	142
rect	126	142	127	143
rect	126	143	127	144
rect	126	144	127	145
rect	126	145	127	146
rect	126	146	127	147
rect	126	147	127	148
rect	126	148	127	149
rect	126	149	127	150
rect	126	150	127	151
rect	126	151	127	152
rect	126	152	127	153
rect	126	153	127	154
rect	126	154	127	155
rect	126	155	127	156
rect	126	156	127	157
rect	126	157	127	158
rect	126	158	127	159
rect	126	160	127	161
rect	126	161	127	162
rect	126	162	127	163
rect	126	163	127	164
rect	126	164	127	165
rect	126	165	127	166
rect	126	166	127	167
rect	126	167	127	168
rect	126	168	127	169
rect	126	169	127	170
rect	126	170	127	171
rect	126	171	127	172
rect	126	172	127	173
rect	126	173	127	174
rect	126	174	127	175
rect	126	175	127	176
rect	126	176	127	177
rect	126	177	127	178
rect	126	178	127	179
rect	126	179	127	180
rect	126	180	127	181
rect	126	181	127	182
rect	126	182	127	183
rect	126	183	127	184
rect	126	185	127	186
rect	126	186	127	187
rect	126	187	127	188
rect	126	188	127	189
rect	126	189	127	190
rect	126	190	127	191
rect	126	192	127	193
rect	126	193	127	194
rect	126	194	127	195
rect	126	195	127	196
rect	126	196	127	197
rect	126	197	127	198
rect	127	0	128	1
rect	127	1	128	2
rect	127	2	128	3
rect	127	3	128	4
rect	127	4	128	5
rect	127	5	128	6
rect	127	6	128	7
rect	127	7	128	8
rect	127	8	128	9
rect	127	9	128	10
rect	127	10	128	11
rect	127	11	128	12
rect	127	12	128	13
rect	127	13	128	14
rect	127	14	128	15
rect	127	15	128	16
rect	127	18	128	19
rect	127	21	128	22
rect	127	24	128	25
rect	127	27	128	28
rect	127	28	128	29
rect	127	29	128	30
rect	127	30	128	31
rect	127	31	128	32
rect	127	32	128	33
rect	127	33	128	34
rect	127	37	128	38
rect	127	38	128	39
rect	127	39	128	40
rect	127	40	128	41
rect	127	41	128	42
rect	127	42	128	43
rect	127	43	128	44
rect	127	44	128	45
rect	127	45	128	46
rect	127	46	128	47
rect	127	47	128	48
rect	127	48	128	49
rect	127	50	128	51
rect	127	51	128	52
rect	127	52	128	53
rect	127	55	128	56
rect	127	56	128	57
rect	127	57	128	58
rect	127	60	128	61
rect	127	61	128	62
rect	127	62	128	63
rect	127	63	128	64
rect	127	64	128	65
rect	127	65	128	66
rect	127	66	128	67
rect	127	67	128	68
rect	127	68	128	69
rect	127	69	128	70
rect	127	70	128	71
rect	127	71	128	72
rect	127	74	128	75
rect	127	75	128	76
rect	127	76	128	77
rect	127	77	128	78
rect	127	78	128	79
rect	127	79	128	80
rect	127	80	128	81
rect	127	81	128	82
rect	127	82	128	83
rect	127	85	128	86
rect	127	87	128	88
rect	127	88	128	89
rect	127	89	128	90
rect	127	90	128	91
rect	127	91	128	92
rect	127	92	128	93
rect	127	93	128	94
rect	127	94	128	95
rect	127	95	128	96
rect	127	96	128	97
rect	127	97	128	98
rect	127	98	128	99
rect	127	99	128	100
rect	127	100	128	101
rect	127	101	128	102
rect	127	103	128	104
rect	127	104	128	105
rect	127	105	128	106
rect	127	106	128	107
rect	127	107	128	108
rect	127	108	128	109
rect	127	109	128	110
rect	127	110	128	111
rect	127	111	128	112
rect	127	112	128	113
rect	127	113	128	114
rect	127	114	128	115
rect	127	115	128	116
rect	127	116	128	117
rect	127	117	128	118
rect	127	119	128	120
rect	127	120	128	121
rect	127	121	128	122
rect	127	122	128	123
rect	127	123	128	124
rect	127	124	128	125
rect	127	125	128	126
rect	127	126	128	127
rect	127	127	128	128
rect	127	128	128	129
rect	127	129	128	130
rect	127	130	128	131
rect	127	131	128	132
rect	127	132	128	133
rect	127	133	128	134
rect	127	134	128	135
rect	127	135	128	136
rect	127	136	128	137
rect	127	137	128	138
rect	127	138	128	139
rect	127	139	128	140
rect	127	141	128	142
rect	127	142	128	143
rect	127	143	128	144
rect	127	144	128	145
rect	127	145	128	146
rect	127	146	128	147
rect	127	147	128	148
rect	127	148	128	149
rect	127	149	128	150
rect	127	150	128	151
rect	127	151	128	152
rect	127	152	128	153
rect	127	153	128	154
rect	127	154	128	155
rect	127	155	128	156
rect	127	156	128	157
rect	127	157	128	158
rect	127	158	128	159
rect	127	160	128	161
rect	127	161	128	162
rect	127	162	128	163
rect	127	163	128	164
rect	127	164	128	165
rect	127	165	128	166
rect	127	166	128	167
rect	127	167	128	168
rect	127	168	128	169
rect	127	169	128	170
rect	127	170	128	171
rect	127	171	128	172
rect	127	172	128	173
rect	127	173	128	174
rect	127	174	128	175
rect	127	175	128	176
rect	127	176	128	177
rect	127	177	128	178
rect	127	178	128	179
rect	127	179	128	180
rect	127	180	128	181
rect	127	181	128	182
rect	127	182	128	183
rect	127	183	128	184
rect	127	185	128	186
rect	127	186	128	187
rect	127	187	128	188
rect	127	188	128	189
rect	127	189	128	190
rect	127	190	128	191
rect	127	192	128	193
rect	127	193	128	194
rect	127	194	128	195
rect	127	195	128	196
rect	127	196	128	197
rect	127	197	128	198
rect	128	0	129	1
rect	128	1	129	2
rect	128	2	129	3
rect	128	3	129	4
rect	128	4	129	5
rect	128	5	129	6
rect	128	6	129	7
rect	128	7	129	8
rect	128	8	129	9
rect	128	9	129	10
rect	128	10	129	11
rect	128	11	129	12
rect	128	12	129	13
rect	128	13	129	14
rect	128	14	129	15
rect	128	15	129	16
rect	128	18	129	19
rect	128	21	129	22
rect	128	24	129	25
rect	128	27	129	28
rect	128	28	129	29
rect	128	29	129	30
rect	128	30	129	31
rect	128	31	129	32
rect	128	32	129	33
rect	128	33	129	34
rect	128	37	129	38
rect	128	38	129	39
rect	128	39	129	40
rect	128	40	129	41
rect	128	41	129	42
rect	128	42	129	43
rect	128	43	129	44
rect	128	44	129	45
rect	128	45	129	46
rect	128	46	129	47
rect	128	47	129	48
rect	128	48	129	49
rect	128	50	129	51
rect	128	51	129	52
rect	128	52	129	53
rect	128	55	129	56
rect	128	56	129	57
rect	128	57	129	58
rect	128	60	129	61
rect	128	61	129	62
rect	128	62	129	63
rect	128	63	129	64
rect	128	64	129	65
rect	128	65	129	66
rect	128	66	129	67
rect	128	67	129	68
rect	128	68	129	69
rect	128	69	129	70
rect	128	70	129	71
rect	128	71	129	72
rect	128	74	129	75
rect	128	75	129	76
rect	128	76	129	77
rect	128	77	129	78
rect	128	78	129	79
rect	128	79	129	80
rect	128	80	129	81
rect	128	81	129	82
rect	128	82	129	83
rect	128	85	129	86
rect	128	87	129	88
rect	128	88	129	89
rect	128	89	129	90
rect	128	90	129	91
rect	128	91	129	92
rect	128	92	129	93
rect	128	93	129	94
rect	128	94	129	95
rect	128	95	129	96
rect	128	96	129	97
rect	128	97	129	98
rect	128	98	129	99
rect	128	99	129	100
rect	128	100	129	101
rect	128	101	129	102
rect	128	103	129	104
rect	128	104	129	105
rect	128	105	129	106
rect	128	106	129	107
rect	128	107	129	108
rect	128	108	129	109
rect	128	109	129	110
rect	128	110	129	111
rect	128	111	129	112
rect	128	112	129	113
rect	128	113	129	114
rect	128	114	129	115
rect	128	115	129	116
rect	128	116	129	117
rect	128	117	129	118
rect	128	119	129	120
rect	128	120	129	121
rect	128	121	129	122
rect	128	122	129	123
rect	128	123	129	124
rect	128	124	129	125
rect	128	125	129	126
rect	128	126	129	127
rect	128	127	129	128
rect	128	128	129	129
rect	128	129	129	130
rect	128	130	129	131
rect	128	131	129	132
rect	128	132	129	133
rect	128	133	129	134
rect	128	134	129	135
rect	128	135	129	136
rect	128	136	129	137
rect	128	137	129	138
rect	128	138	129	139
rect	128	139	129	140
rect	128	141	129	142
rect	128	142	129	143
rect	128	143	129	144
rect	128	144	129	145
rect	128	145	129	146
rect	128	146	129	147
rect	128	147	129	148
rect	128	148	129	149
rect	128	149	129	150
rect	128	150	129	151
rect	128	151	129	152
rect	128	152	129	153
rect	128	153	129	154
rect	128	154	129	155
rect	128	155	129	156
rect	128	156	129	157
rect	128	157	129	158
rect	128	158	129	159
rect	128	160	129	161
rect	128	161	129	162
rect	128	162	129	163
rect	128	163	129	164
rect	128	164	129	165
rect	128	165	129	166
rect	128	166	129	167
rect	128	167	129	168
rect	128	168	129	169
rect	128	169	129	170
rect	128	170	129	171
rect	128	171	129	172
rect	128	172	129	173
rect	128	173	129	174
rect	128	174	129	175
rect	128	175	129	176
rect	128	176	129	177
rect	128	177	129	178
rect	128	178	129	179
rect	128	179	129	180
rect	128	180	129	181
rect	128	181	129	182
rect	128	182	129	183
rect	128	183	129	184
rect	128	185	129	186
rect	128	186	129	187
rect	128	187	129	188
rect	128	188	129	189
rect	128	189	129	190
rect	128	190	129	191
rect	128	192	129	193
rect	128	193	129	194
rect	128	194	129	195
rect	128	195	129	196
rect	128	196	129	197
rect	128	197	129	198
rect	129	0	130	1
rect	129	1	130	2
rect	129	2	130	3
rect	129	3	130	4
rect	129	4	130	5
rect	129	5	130	6
rect	129	6	130	7
rect	129	7	130	8
rect	129	8	130	9
rect	129	9	130	10
rect	129	10	130	11
rect	129	11	130	12
rect	129	12	130	13
rect	129	13	130	14
rect	129	14	130	15
rect	129	15	130	16
rect	129	18	130	19
rect	129	21	130	22
rect	129	24	130	25
rect	129	27	130	28
rect	129	28	130	29
rect	129	29	130	30
rect	129	30	130	31
rect	129	31	130	32
rect	129	32	130	33
rect	129	33	130	34
rect	129	37	130	38
rect	129	38	130	39
rect	129	39	130	40
rect	129	40	130	41
rect	129	41	130	42
rect	129	42	130	43
rect	129	43	130	44
rect	129	44	130	45
rect	129	45	130	46
rect	129	46	130	47
rect	129	47	130	48
rect	129	48	130	49
rect	129	50	130	51
rect	129	51	130	52
rect	129	52	130	53
rect	129	55	130	56
rect	129	56	130	57
rect	129	57	130	58
rect	129	60	130	61
rect	129	61	130	62
rect	129	62	130	63
rect	129	63	130	64
rect	129	64	130	65
rect	129	65	130	66
rect	129	66	130	67
rect	129	67	130	68
rect	129	68	130	69
rect	129	69	130	70
rect	129	70	130	71
rect	129	71	130	72
rect	129	74	130	75
rect	129	75	130	76
rect	129	76	130	77
rect	129	77	130	78
rect	129	78	130	79
rect	129	79	130	80
rect	129	80	130	81
rect	129	81	130	82
rect	129	82	130	83
rect	129	85	130	86
rect	129	87	130	88
rect	129	88	130	89
rect	129	89	130	90
rect	129	90	130	91
rect	129	91	130	92
rect	129	92	130	93
rect	129	93	130	94
rect	129	94	130	95
rect	129	95	130	96
rect	129	96	130	97
rect	129	97	130	98
rect	129	98	130	99
rect	129	99	130	100
rect	129	100	130	101
rect	129	101	130	102
rect	129	103	130	104
rect	129	104	130	105
rect	129	105	130	106
rect	129	106	130	107
rect	129	107	130	108
rect	129	108	130	109
rect	129	109	130	110
rect	129	110	130	111
rect	129	111	130	112
rect	129	112	130	113
rect	129	113	130	114
rect	129	114	130	115
rect	129	115	130	116
rect	129	116	130	117
rect	129	117	130	118
rect	129	119	130	120
rect	129	120	130	121
rect	129	121	130	122
rect	129	122	130	123
rect	129	123	130	124
rect	129	124	130	125
rect	129	125	130	126
rect	129	126	130	127
rect	129	127	130	128
rect	129	128	130	129
rect	129	129	130	130
rect	129	130	130	131
rect	129	131	130	132
rect	129	132	130	133
rect	129	133	130	134
rect	129	134	130	135
rect	129	135	130	136
rect	129	136	130	137
rect	129	137	130	138
rect	129	138	130	139
rect	129	139	130	140
rect	129	141	130	142
rect	129	142	130	143
rect	129	143	130	144
rect	129	144	130	145
rect	129	145	130	146
rect	129	146	130	147
rect	129	147	130	148
rect	129	148	130	149
rect	129	149	130	150
rect	129	150	130	151
rect	129	151	130	152
rect	129	152	130	153
rect	129	153	130	154
rect	129	154	130	155
rect	129	155	130	156
rect	129	156	130	157
rect	129	157	130	158
rect	129	158	130	159
rect	129	160	130	161
rect	129	161	130	162
rect	129	162	130	163
rect	129	163	130	164
rect	129	164	130	165
rect	129	165	130	166
rect	129	166	130	167
rect	129	167	130	168
rect	129	168	130	169
rect	129	169	130	170
rect	129	170	130	171
rect	129	171	130	172
rect	129	172	130	173
rect	129	173	130	174
rect	129	174	130	175
rect	129	175	130	176
rect	129	176	130	177
rect	129	177	130	178
rect	129	178	130	179
rect	129	179	130	180
rect	129	180	130	181
rect	129	181	130	182
rect	129	182	130	183
rect	129	183	130	184
rect	129	185	130	186
rect	129	186	130	187
rect	129	187	130	188
rect	129	188	130	189
rect	129	189	130	190
rect	129	190	130	191
rect	129	192	130	193
rect	129	193	130	194
rect	129	194	130	195
rect	129	195	130	196
rect	129	196	130	197
rect	129	197	130	198
rect	130	0	131	1
rect	130	1	131	2
rect	130	2	131	3
rect	130	3	131	4
rect	130	4	131	5
rect	130	5	131	6
rect	130	6	131	7
rect	130	7	131	8
rect	130	8	131	9
rect	130	9	131	10
rect	130	10	131	11
rect	130	11	131	12
rect	130	12	131	13
rect	130	13	131	14
rect	130	14	131	15
rect	130	15	131	16
rect	130	18	131	19
rect	130	21	131	22
rect	130	24	131	25
rect	130	27	131	28
rect	130	28	131	29
rect	130	29	131	30
rect	130	30	131	31
rect	130	31	131	32
rect	130	32	131	33
rect	130	33	131	34
rect	130	37	131	38
rect	130	38	131	39
rect	130	39	131	40
rect	130	40	131	41
rect	130	41	131	42
rect	130	42	131	43
rect	130	43	131	44
rect	130	44	131	45
rect	130	45	131	46
rect	130	46	131	47
rect	130	47	131	48
rect	130	48	131	49
rect	130	50	131	51
rect	130	51	131	52
rect	130	52	131	53
rect	130	55	131	56
rect	130	56	131	57
rect	130	57	131	58
rect	130	60	131	61
rect	130	61	131	62
rect	130	62	131	63
rect	130	63	131	64
rect	130	64	131	65
rect	130	65	131	66
rect	130	66	131	67
rect	130	67	131	68
rect	130	68	131	69
rect	130	69	131	70
rect	130	70	131	71
rect	130	71	131	72
rect	130	74	131	75
rect	130	75	131	76
rect	130	76	131	77
rect	130	77	131	78
rect	130	78	131	79
rect	130	79	131	80
rect	130	80	131	81
rect	130	81	131	82
rect	130	82	131	83
rect	130	85	131	86
rect	130	87	131	88
rect	130	88	131	89
rect	130	89	131	90
rect	130	90	131	91
rect	130	91	131	92
rect	130	92	131	93
rect	130	93	131	94
rect	130	94	131	95
rect	130	95	131	96
rect	130	96	131	97
rect	130	97	131	98
rect	130	98	131	99
rect	130	99	131	100
rect	130	100	131	101
rect	130	101	131	102
rect	130	103	131	104
rect	130	104	131	105
rect	130	105	131	106
rect	130	106	131	107
rect	130	107	131	108
rect	130	108	131	109
rect	130	109	131	110
rect	130	110	131	111
rect	130	111	131	112
rect	130	112	131	113
rect	130	113	131	114
rect	130	114	131	115
rect	130	115	131	116
rect	130	116	131	117
rect	130	117	131	118
rect	130	119	131	120
rect	130	120	131	121
rect	130	121	131	122
rect	130	122	131	123
rect	130	123	131	124
rect	130	124	131	125
rect	130	125	131	126
rect	130	126	131	127
rect	130	127	131	128
rect	130	128	131	129
rect	130	129	131	130
rect	130	130	131	131
rect	130	131	131	132
rect	130	132	131	133
rect	130	133	131	134
rect	130	134	131	135
rect	130	135	131	136
rect	130	136	131	137
rect	130	137	131	138
rect	130	138	131	139
rect	130	139	131	140
rect	130	141	131	142
rect	130	142	131	143
rect	130	143	131	144
rect	130	144	131	145
rect	130	145	131	146
rect	130	146	131	147
rect	130	147	131	148
rect	130	148	131	149
rect	130	149	131	150
rect	130	150	131	151
rect	130	151	131	152
rect	130	152	131	153
rect	130	153	131	154
rect	130	154	131	155
rect	130	155	131	156
rect	130	156	131	157
rect	130	157	131	158
rect	130	158	131	159
rect	130	160	131	161
rect	130	161	131	162
rect	130	162	131	163
rect	130	163	131	164
rect	130	164	131	165
rect	130	165	131	166
rect	130	166	131	167
rect	130	167	131	168
rect	130	168	131	169
rect	130	169	131	170
rect	130	170	131	171
rect	130	171	131	172
rect	130	172	131	173
rect	130	173	131	174
rect	130	174	131	175
rect	130	175	131	176
rect	130	176	131	177
rect	130	177	131	178
rect	130	178	131	179
rect	130	179	131	180
rect	130	180	131	181
rect	130	181	131	182
rect	130	182	131	183
rect	130	183	131	184
rect	130	185	131	186
rect	130	186	131	187
rect	130	187	131	188
rect	130	188	131	189
rect	130	189	131	190
rect	130	190	131	191
rect	130	192	131	193
rect	130	193	131	194
rect	130	194	131	195
rect	130	195	131	196
rect	130	196	131	197
rect	130	197	131	198
rect	131	0	132	1
rect	131	1	132	2
rect	131	2	132	3
rect	131	3	132	4
rect	131	4	132	5
rect	131	5	132	6
rect	131	6	132	7
rect	131	7	132	8
rect	131	8	132	9
rect	131	9	132	10
rect	131	10	132	11
rect	131	11	132	12
rect	131	12	132	13
rect	131	13	132	14
rect	131	14	132	15
rect	131	15	132	16
rect	131	18	132	19
rect	131	21	132	22
rect	131	24	132	25
rect	131	27	132	28
rect	131	28	132	29
rect	131	29	132	30
rect	131	30	132	31
rect	131	31	132	32
rect	131	32	132	33
rect	131	33	132	34
rect	131	34	132	35
rect	131	37	132	38
rect	131	38	132	39
rect	131	39	132	40
rect	131	40	132	41
rect	131	41	132	42
rect	131	42	132	43
rect	131	43	132	44
rect	131	44	132	45
rect	131	45	132	46
rect	131	46	132	47
rect	131	47	132	48
rect	131	48	132	49
rect	131	50	132	51
rect	131	51	132	52
rect	131	52	132	53
rect	131	55	132	56
rect	131	56	132	57
rect	131	57	132	58
rect	131	60	132	61
rect	131	61	132	62
rect	131	62	132	63
rect	131	63	132	64
rect	131	64	132	65
rect	131	65	132	66
rect	131	66	132	67
rect	131	67	132	68
rect	131	68	132	69
rect	131	69	132	70
rect	131	70	132	71
rect	131	71	132	72
rect	131	74	132	75
rect	131	75	132	76
rect	131	76	132	77
rect	131	77	132	78
rect	131	78	132	79
rect	131	79	132	80
rect	131	80	132	81
rect	131	81	132	82
rect	131	82	132	83
rect	131	85	132	86
rect	131	87	132	88
rect	131	88	132	89
rect	131	89	132	90
rect	131	90	132	91
rect	131	91	132	92
rect	131	92	132	93
rect	131	93	132	94
rect	131	94	132	95
rect	131	95	132	96
rect	131	96	132	97
rect	131	97	132	98
rect	131	98	132	99
rect	131	99	132	100
rect	131	100	132	101
rect	131	101	132	102
rect	131	103	132	104
rect	131	104	132	105
rect	131	105	132	106
rect	131	106	132	107
rect	131	107	132	108
rect	131	108	132	109
rect	131	109	132	110
rect	131	110	132	111
rect	131	111	132	112
rect	131	112	132	113
rect	131	113	132	114
rect	131	114	132	115
rect	131	115	132	116
rect	131	116	132	117
rect	131	117	132	118
rect	131	119	132	120
rect	131	120	132	121
rect	131	121	132	122
rect	131	122	132	123
rect	131	123	132	124
rect	131	124	132	125
rect	131	125	132	126
rect	131	126	132	127
rect	131	127	132	128
rect	131	128	132	129
rect	131	129	132	130
rect	131	130	132	131
rect	131	131	132	132
rect	131	132	132	133
rect	131	133	132	134
rect	131	134	132	135
rect	131	135	132	136
rect	131	136	132	137
rect	131	137	132	138
rect	131	138	132	139
rect	131	139	132	140
rect	131	141	132	142
rect	131	142	132	143
rect	131	143	132	144
rect	131	144	132	145
rect	131	145	132	146
rect	131	146	132	147
rect	131	147	132	148
rect	131	148	132	149
rect	131	149	132	150
rect	131	150	132	151
rect	131	151	132	152
rect	131	152	132	153
rect	131	153	132	154
rect	131	154	132	155
rect	131	155	132	156
rect	131	156	132	157
rect	131	157	132	158
rect	131	158	132	159
rect	131	160	132	161
rect	131	161	132	162
rect	131	162	132	163
rect	131	163	132	164
rect	131	164	132	165
rect	131	165	132	166
rect	131	166	132	167
rect	131	167	132	168
rect	131	168	132	169
rect	131	169	132	170
rect	131	170	132	171
rect	131	171	132	172
rect	131	172	132	173
rect	131	173	132	174
rect	131	174	132	175
rect	131	175	132	176
rect	131	176	132	177
rect	131	177	132	178
rect	131	178	132	179
rect	131	179	132	180
rect	131	180	132	181
rect	131	181	132	182
rect	131	182	132	183
rect	131	183	132	184
rect	131	185	132	186
rect	131	186	132	187
rect	131	187	132	188
rect	131	188	132	189
rect	131	189	132	190
rect	131	190	132	191
rect	131	192	132	193
rect	131	193	132	194
rect	131	194	132	195
rect	131	195	132	196
rect	131	196	132	197
rect	131	197	132	198
rect	171	0	172	1
rect	171	1	172	2
rect	171	2	172	3
rect	171	3	172	4
rect	171	4	172	5
rect	171	5	172	6
rect	171	6	172	7
rect	171	7	172	8
rect	171	8	172	9
rect	171	9	172	10
rect	171	10	172	11
rect	171	11	172	12
rect	171	12	172	13
rect	171	13	172	14
rect	171	14	172	15
rect	171	15	172	16
rect	171	18	172	19
rect	171	21	172	22
rect	171	24	172	25
rect	171	25	172	26
rect	171	28	172	29
rect	171	29	172	30
rect	171	30	172	31
rect	171	31	172	32
rect	171	32	172	33
rect	171	33	172	34
rect	171	34	172	35
rect	171	35	172	36
rect	171	36	172	37
rect	171	37	172	38
rect	171	38	172	39
rect	171	39	172	40
rect	171	40	172	41
rect	171	41	172	42
rect	171	42	172	43
rect	171	43	172	44
rect	171	44	172	45
rect	171	45	172	46
rect	171	46	172	47
rect	171	47	172	48
rect	171	48	172	49
rect	171	49	172	50
rect	171	50	172	51
rect	171	51	172	52
rect	171	52	172	53
rect	171	55	172	56
rect	171	56	172	57
rect	171	57	172	58
rect	171	60	172	61
rect	171	61	172	62
rect	171	62	172	63
rect	171	63	172	64
rect	171	65	172	66
rect	171	66	172	67
rect	171	67	172	68
rect	171	68	172	69
rect	171	69	172	70
rect	171	70	172	71
rect	171	71	172	72
rect	171	74	172	75
rect	171	75	172	76
rect	171	76	172	77
rect	171	77	172	78
rect	171	78	172	79
rect	171	79	172	80
rect	171	80	172	81
rect	171	81	172	82
rect	171	82	172	83
rect	171	85	172	86
rect	171	86	172	87
rect	171	87	172	88
rect	171	88	172	89
rect	171	89	172	90
rect	171	90	172	91
rect	171	91	172	92
rect	171	93	172	94
rect	171	94	172	95
rect	171	95	172	96
rect	171	96	172	97
rect	171	97	172	98
rect	171	98	172	99
rect	171	99	172	100
rect	171	100	172	101
rect	171	101	172	102
rect	171	102	172	103
rect	171	103	172	104
rect	171	104	172	105
rect	171	105	172	106
rect	171	106	172	107
rect	171	107	172	108
rect	171	109	172	110
rect	171	110	172	111
rect	171	111	172	112
rect	171	112	172	113
rect	171	113	172	114
rect	171	114	172	115
rect	171	115	172	116
rect	171	116	172	117
rect	171	117	172	118
rect	171	118	172	119
rect	171	119	172	120
rect	171	120	172	121
rect	171	122	172	123
rect	171	123	172	124
rect	171	124	172	125
rect	171	125	172	126
rect	171	126	172	127
rect	171	127	172	128
rect	171	128	172	129
rect	171	129	172	130
rect	171	130	172	131
rect	171	131	172	132
rect	171	132	172	133
rect	171	133	172	134
rect	171	134	172	135
rect	171	135	172	136
rect	171	136	172	137
rect	171	138	172	139
rect	171	139	172	140
rect	171	140	172	141
rect	171	141	172	142
rect	171	142	172	143
rect	171	143	172	144
rect	171	144	172	145
rect	171	145	172	146
rect	171	146	172	147
rect	171	147	172	148
rect	171	148	172	149
rect	171	149	172	150
rect	171	150	172	151
rect	171	151	172	152
rect	171	152	172	153
rect	171	153	172	154
rect	171	154	172	155
rect	171	155	172	156
rect	171	156	172	157
rect	171	157	172	158
rect	171	158	172	159
rect	171	160	172	161
rect	171	161	172	162
rect	171	162	172	163
rect	171	163	172	164
rect	171	164	172	165
rect	171	165	172	166
rect	171	166	172	167
rect	171	167	172	168
rect	171	168	172	169
rect	171	169	172	170
rect	171	170	172	171
rect	171	171	172	172
rect	171	173	172	174
rect	171	174	172	175
rect	171	175	172	176
rect	171	176	172	177
rect	171	177	172	178
rect	171	178	172	179
rect	171	179	172	180
rect	171	180	172	181
rect	171	181	172	182
rect	171	182	172	183
rect	171	183	172	184
rect	171	184	172	185
rect	171	186	172	187
rect	171	187	172	188
rect	171	188	172	189
rect	171	189	172	190
rect	171	190	172	191
rect	171	191	172	192
rect	172	0	173	1
rect	172	1	173	2
rect	172	2	173	3
rect	172	3	173	4
rect	172	4	173	5
rect	172	5	173	6
rect	172	6	173	7
rect	172	7	173	8
rect	172	8	173	9
rect	172	9	173	10
rect	172	10	173	11
rect	172	11	173	12
rect	172	12	173	13
rect	172	13	173	14
rect	172	14	173	15
rect	172	15	173	16
rect	172	18	173	19
rect	172	21	173	22
rect	172	24	173	25
rect	172	25	173	26
rect	172	28	173	29
rect	172	29	173	30
rect	172	30	173	31
rect	172	31	173	32
rect	172	32	173	33
rect	172	33	173	34
rect	172	34	173	35
rect	172	35	173	36
rect	172	36	173	37
rect	172	37	173	38
rect	172	38	173	39
rect	172	39	173	40
rect	172	40	173	41
rect	172	41	173	42
rect	172	42	173	43
rect	172	43	173	44
rect	172	44	173	45
rect	172	45	173	46
rect	172	46	173	47
rect	172	47	173	48
rect	172	48	173	49
rect	172	49	173	50
rect	172	50	173	51
rect	172	51	173	52
rect	172	52	173	53
rect	172	55	173	56
rect	172	56	173	57
rect	172	57	173	58
rect	172	60	173	61
rect	172	61	173	62
rect	172	62	173	63
rect	172	63	173	64
rect	172	65	173	66
rect	172	66	173	67
rect	172	67	173	68
rect	172	68	173	69
rect	172	69	173	70
rect	172	70	173	71
rect	172	71	173	72
rect	172	74	173	75
rect	172	75	173	76
rect	172	76	173	77
rect	172	77	173	78
rect	172	78	173	79
rect	172	79	173	80
rect	172	80	173	81
rect	172	81	173	82
rect	172	82	173	83
rect	172	85	173	86
rect	172	86	173	87
rect	172	87	173	88
rect	172	88	173	89
rect	172	89	173	90
rect	172	90	173	91
rect	172	91	173	92
rect	172	93	173	94
rect	172	94	173	95
rect	172	95	173	96
rect	172	96	173	97
rect	172	97	173	98
rect	172	98	173	99
rect	172	99	173	100
rect	172	100	173	101
rect	172	101	173	102
rect	172	102	173	103
rect	172	103	173	104
rect	172	104	173	105
rect	172	105	173	106
rect	172	106	173	107
rect	172	107	173	108
rect	172	109	173	110
rect	172	110	173	111
rect	172	111	173	112
rect	172	112	173	113
rect	172	113	173	114
rect	172	114	173	115
rect	172	115	173	116
rect	172	116	173	117
rect	172	117	173	118
rect	172	118	173	119
rect	172	119	173	120
rect	172	120	173	121
rect	172	122	173	123
rect	172	123	173	124
rect	172	124	173	125
rect	172	125	173	126
rect	172	126	173	127
rect	172	127	173	128
rect	172	128	173	129
rect	172	129	173	130
rect	172	130	173	131
rect	172	131	173	132
rect	172	132	173	133
rect	172	133	173	134
rect	172	134	173	135
rect	172	135	173	136
rect	172	136	173	137
rect	172	138	173	139
rect	172	139	173	140
rect	172	140	173	141
rect	172	141	173	142
rect	172	142	173	143
rect	172	143	173	144
rect	172	144	173	145
rect	172	145	173	146
rect	172	146	173	147
rect	172	147	173	148
rect	172	148	173	149
rect	172	149	173	150
rect	172	150	173	151
rect	172	151	173	152
rect	172	152	173	153
rect	172	153	173	154
rect	172	154	173	155
rect	172	155	173	156
rect	172	156	173	157
rect	172	157	173	158
rect	172	158	173	159
rect	172	160	173	161
rect	172	161	173	162
rect	172	162	173	163
rect	172	163	173	164
rect	172	164	173	165
rect	172	165	173	166
rect	172	166	173	167
rect	172	167	173	168
rect	172	168	173	169
rect	172	169	173	170
rect	172	170	173	171
rect	172	171	173	172
rect	172	173	173	174
rect	172	174	173	175
rect	172	175	173	176
rect	172	176	173	177
rect	172	177	173	178
rect	172	178	173	179
rect	172	179	173	180
rect	172	180	173	181
rect	172	181	173	182
rect	172	182	173	183
rect	172	183	173	184
rect	172	184	173	185
rect	172	186	173	187
rect	172	187	173	188
rect	172	188	173	189
rect	172	189	173	190
rect	172	190	173	191
rect	172	191	173	192
rect	173	0	174	1
rect	173	1	174	2
rect	173	2	174	3
rect	173	3	174	4
rect	173	4	174	5
rect	173	5	174	6
rect	173	6	174	7
rect	173	7	174	8
rect	173	8	174	9
rect	173	9	174	10
rect	173	10	174	11
rect	173	11	174	12
rect	173	12	174	13
rect	173	13	174	14
rect	173	14	174	15
rect	173	15	174	16
rect	173	18	174	19
rect	173	21	174	22
rect	173	24	174	25
rect	173	25	174	26
rect	173	28	174	29
rect	173	29	174	30
rect	173	30	174	31
rect	173	31	174	32
rect	173	32	174	33
rect	173	33	174	34
rect	173	34	174	35
rect	173	35	174	36
rect	173	36	174	37
rect	173	37	174	38
rect	173	38	174	39
rect	173	39	174	40
rect	173	40	174	41
rect	173	41	174	42
rect	173	42	174	43
rect	173	43	174	44
rect	173	44	174	45
rect	173	45	174	46
rect	173	46	174	47
rect	173	47	174	48
rect	173	48	174	49
rect	173	49	174	50
rect	173	50	174	51
rect	173	51	174	52
rect	173	52	174	53
rect	173	55	174	56
rect	173	56	174	57
rect	173	57	174	58
rect	173	60	174	61
rect	173	61	174	62
rect	173	62	174	63
rect	173	63	174	64
rect	173	65	174	66
rect	173	66	174	67
rect	173	67	174	68
rect	173	68	174	69
rect	173	69	174	70
rect	173	70	174	71
rect	173	71	174	72
rect	173	74	174	75
rect	173	75	174	76
rect	173	76	174	77
rect	173	77	174	78
rect	173	78	174	79
rect	173	79	174	80
rect	173	80	174	81
rect	173	81	174	82
rect	173	82	174	83
rect	173	85	174	86
rect	173	86	174	87
rect	173	87	174	88
rect	173	88	174	89
rect	173	89	174	90
rect	173	90	174	91
rect	173	91	174	92
rect	173	93	174	94
rect	173	94	174	95
rect	173	95	174	96
rect	173	96	174	97
rect	173	97	174	98
rect	173	98	174	99
rect	173	99	174	100
rect	173	100	174	101
rect	173	101	174	102
rect	173	102	174	103
rect	173	103	174	104
rect	173	104	174	105
rect	173	105	174	106
rect	173	106	174	107
rect	173	107	174	108
rect	173	109	174	110
rect	173	110	174	111
rect	173	111	174	112
rect	173	112	174	113
rect	173	113	174	114
rect	173	114	174	115
rect	173	115	174	116
rect	173	116	174	117
rect	173	117	174	118
rect	173	118	174	119
rect	173	119	174	120
rect	173	120	174	121
rect	173	122	174	123
rect	173	123	174	124
rect	173	124	174	125
rect	173	125	174	126
rect	173	126	174	127
rect	173	127	174	128
rect	173	128	174	129
rect	173	129	174	130
rect	173	130	174	131
rect	173	131	174	132
rect	173	132	174	133
rect	173	133	174	134
rect	173	134	174	135
rect	173	135	174	136
rect	173	136	174	137
rect	173	138	174	139
rect	173	139	174	140
rect	173	140	174	141
rect	173	141	174	142
rect	173	142	174	143
rect	173	143	174	144
rect	173	144	174	145
rect	173	145	174	146
rect	173	146	174	147
rect	173	147	174	148
rect	173	148	174	149
rect	173	149	174	150
rect	173	150	174	151
rect	173	151	174	152
rect	173	152	174	153
rect	173	153	174	154
rect	173	154	174	155
rect	173	155	174	156
rect	173	156	174	157
rect	173	157	174	158
rect	173	158	174	159
rect	173	160	174	161
rect	173	161	174	162
rect	173	162	174	163
rect	173	163	174	164
rect	173	164	174	165
rect	173	165	174	166
rect	173	166	174	167
rect	173	167	174	168
rect	173	168	174	169
rect	173	169	174	170
rect	173	170	174	171
rect	173	171	174	172
rect	173	173	174	174
rect	173	174	174	175
rect	173	175	174	176
rect	173	176	174	177
rect	173	177	174	178
rect	173	178	174	179
rect	173	179	174	180
rect	173	180	174	181
rect	173	181	174	182
rect	173	182	174	183
rect	173	183	174	184
rect	173	184	174	185
rect	173	186	174	187
rect	173	187	174	188
rect	173	188	174	189
rect	173	189	174	190
rect	173	190	174	191
rect	173	191	174	192
rect	174	0	175	1
rect	174	1	175	2
rect	174	2	175	3
rect	174	3	175	4
rect	174	4	175	5
rect	174	5	175	6
rect	174	6	175	7
rect	174	7	175	8
rect	174	8	175	9
rect	174	9	175	10
rect	174	10	175	11
rect	174	11	175	12
rect	174	12	175	13
rect	174	13	175	14
rect	174	14	175	15
rect	174	15	175	16
rect	174	18	175	19
rect	174	21	175	22
rect	174	24	175	25
rect	174	25	175	26
rect	174	28	175	29
rect	174	29	175	30
rect	174	30	175	31
rect	174	31	175	32
rect	174	32	175	33
rect	174	33	175	34
rect	174	34	175	35
rect	174	35	175	36
rect	174	36	175	37
rect	174	37	175	38
rect	174	38	175	39
rect	174	39	175	40
rect	174	40	175	41
rect	174	41	175	42
rect	174	42	175	43
rect	174	43	175	44
rect	174	44	175	45
rect	174	45	175	46
rect	174	46	175	47
rect	174	47	175	48
rect	174	48	175	49
rect	174	49	175	50
rect	174	50	175	51
rect	174	51	175	52
rect	174	52	175	53
rect	174	55	175	56
rect	174	56	175	57
rect	174	57	175	58
rect	174	60	175	61
rect	174	61	175	62
rect	174	62	175	63
rect	174	63	175	64
rect	174	65	175	66
rect	174	66	175	67
rect	174	67	175	68
rect	174	68	175	69
rect	174	69	175	70
rect	174	70	175	71
rect	174	71	175	72
rect	174	74	175	75
rect	174	75	175	76
rect	174	76	175	77
rect	174	77	175	78
rect	174	78	175	79
rect	174	79	175	80
rect	174	80	175	81
rect	174	81	175	82
rect	174	82	175	83
rect	174	85	175	86
rect	174	86	175	87
rect	174	87	175	88
rect	174	88	175	89
rect	174	89	175	90
rect	174	90	175	91
rect	174	91	175	92
rect	174	93	175	94
rect	174	94	175	95
rect	174	95	175	96
rect	174	96	175	97
rect	174	97	175	98
rect	174	98	175	99
rect	174	99	175	100
rect	174	100	175	101
rect	174	101	175	102
rect	174	102	175	103
rect	174	103	175	104
rect	174	104	175	105
rect	174	105	175	106
rect	174	106	175	107
rect	174	107	175	108
rect	174	109	175	110
rect	174	110	175	111
rect	174	111	175	112
rect	174	112	175	113
rect	174	113	175	114
rect	174	114	175	115
rect	174	115	175	116
rect	174	116	175	117
rect	174	117	175	118
rect	174	118	175	119
rect	174	119	175	120
rect	174	120	175	121
rect	174	122	175	123
rect	174	123	175	124
rect	174	124	175	125
rect	174	125	175	126
rect	174	126	175	127
rect	174	127	175	128
rect	174	128	175	129
rect	174	129	175	130
rect	174	130	175	131
rect	174	131	175	132
rect	174	132	175	133
rect	174	133	175	134
rect	174	134	175	135
rect	174	135	175	136
rect	174	136	175	137
rect	174	138	175	139
rect	174	139	175	140
rect	174	140	175	141
rect	174	141	175	142
rect	174	142	175	143
rect	174	143	175	144
rect	174	144	175	145
rect	174	145	175	146
rect	174	146	175	147
rect	174	147	175	148
rect	174	148	175	149
rect	174	149	175	150
rect	174	150	175	151
rect	174	151	175	152
rect	174	152	175	153
rect	174	153	175	154
rect	174	154	175	155
rect	174	155	175	156
rect	174	156	175	157
rect	174	157	175	158
rect	174	158	175	159
rect	174	160	175	161
rect	174	161	175	162
rect	174	162	175	163
rect	174	163	175	164
rect	174	164	175	165
rect	174	165	175	166
rect	174	166	175	167
rect	174	167	175	168
rect	174	168	175	169
rect	174	169	175	170
rect	174	170	175	171
rect	174	171	175	172
rect	174	173	175	174
rect	174	174	175	175
rect	174	175	175	176
rect	174	176	175	177
rect	174	177	175	178
rect	174	178	175	179
rect	174	179	175	180
rect	174	180	175	181
rect	174	181	175	182
rect	174	182	175	183
rect	174	183	175	184
rect	174	184	175	185
rect	174	186	175	187
rect	174	187	175	188
rect	174	188	175	189
rect	174	189	175	190
rect	174	190	175	191
rect	174	191	175	192
rect	175	0	176	1
rect	175	1	176	2
rect	175	2	176	3
rect	175	3	176	4
rect	175	4	176	5
rect	175	5	176	6
rect	175	6	176	7
rect	175	7	176	8
rect	175	8	176	9
rect	175	9	176	10
rect	175	10	176	11
rect	175	11	176	12
rect	175	12	176	13
rect	175	13	176	14
rect	175	14	176	15
rect	175	15	176	16
rect	175	18	176	19
rect	175	21	176	22
rect	175	24	176	25
rect	175	25	176	26
rect	175	28	176	29
rect	175	29	176	30
rect	175	30	176	31
rect	175	31	176	32
rect	175	32	176	33
rect	175	33	176	34
rect	175	34	176	35
rect	175	35	176	36
rect	175	36	176	37
rect	175	37	176	38
rect	175	38	176	39
rect	175	39	176	40
rect	175	40	176	41
rect	175	41	176	42
rect	175	42	176	43
rect	175	43	176	44
rect	175	44	176	45
rect	175	45	176	46
rect	175	46	176	47
rect	175	47	176	48
rect	175	48	176	49
rect	175	49	176	50
rect	175	50	176	51
rect	175	51	176	52
rect	175	52	176	53
rect	175	55	176	56
rect	175	56	176	57
rect	175	57	176	58
rect	175	60	176	61
rect	175	61	176	62
rect	175	62	176	63
rect	175	63	176	64
rect	175	65	176	66
rect	175	66	176	67
rect	175	67	176	68
rect	175	68	176	69
rect	175	69	176	70
rect	175	70	176	71
rect	175	71	176	72
rect	175	74	176	75
rect	175	75	176	76
rect	175	76	176	77
rect	175	77	176	78
rect	175	78	176	79
rect	175	79	176	80
rect	175	80	176	81
rect	175	81	176	82
rect	175	82	176	83
rect	175	85	176	86
rect	175	86	176	87
rect	175	87	176	88
rect	175	88	176	89
rect	175	89	176	90
rect	175	90	176	91
rect	175	91	176	92
rect	175	93	176	94
rect	175	94	176	95
rect	175	95	176	96
rect	175	96	176	97
rect	175	97	176	98
rect	175	98	176	99
rect	175	99	176	100
rect	175	100	176	101
rect	175	101	176	102
rect	175	102	176	103
rect	175	103	176	104
rect	175	104	176	105
rect	175	105	176	106
rect	175	106	176	107
rect	175	107	176	108
rect	175	109	176	110
rect	175	110	176	111
rect	175	111	176	112
rect	175	112	176	113
rect	175	113	176	114
rect	175	114	176	115
rect	175	115	176	116
rect	175	116	176	117
rect	175	117	176	118
rect	175	118	176	119
rect	175	119	176	120
rect	175	120	176	121
rect	175	122	176	123
rect	175	123	176	124
rect	175	124	176	125
rect	175	125	176	126
rect	175	126	176	127
rect	175	127	176	128
rect	175	128	176	129
rect	175	129	176	130
rect	175	130	176	131
rect	175	131	176	132
rect	175	132	176	133
rect	175	133	176	134
rect	175	134	176	135
rect	175	135	176	136
rect	175	136	176	137
rect	175	138	176	139
rect	175	139	176	140
rect	175	140	176	141
rect	175	141	176	142
rect	175	142	176	143
rect	175	143	176	144
rect	175	144	176	145
rect	175	145	176	146
rect	175	146	176	147
rect	175	147	176	148
rect	175	148	176	149
rect	175	149	176	150
rect	175	150	176	151
rect	175	151	176	152
rect	175	152	176	153
rect	175	153	176	154
rect	175	154	176	155
rect	175	155	176	156
rect	175	156	176	157
rect	175	157	176	158
rect	175	158	176	159
rect	175	160	176	161
rect	175	161	176	162
rect	175	162	176	163
rect	175	163	176	164
rect	175	164	176	165
rect	175	165	176	166
rect	175	166	176	167
rect	175	167	176	168
rect	175	168	176	169
rect	175	169	176	170
rect	175	170	176	171
rect	175	171	176	172
rect	175	173	176	174
rect	175	174	176	175
rect	175	175	176	176
rect	175	176	176	177
rect	175	177	176	178
rect	175	178	176	179
rect	175	179	176	180
rect	175	180	176	181
rect	175	181	176	182
rect	175	182	176	183
rect	175	183	176	184
rect	175	184	176	185
rect	175	186	176	187
rect	175	187	176	188
rect	175	188	176	189
rect	175	189	176	190
rect	175	190	176	191
rect	175	191	176	192
rect	176	0	177	1
rect	176	1	177	2
rect	176	2	177	3
rect	176	3	177	4
rect	176	4	177	5
rect	176	5	177	6
rect	176	6	177	7
rect	176	7	177	8
rect	176	8	177	9
rect	176	9	177	10
rect	176	10	177	11
rect	176	11	177	12
rect	176	12	177	13
rect	176	13	177	14
rect	176	14	177	15
rect	176	15	177	16
rect	176	16	177	17
rect	176	18	177	19
rect	176	19	177	20
rect	176	21	177	22
rect	176	22	177	23
rect	176	24	177	25
rect	176	25	177	26
rect	176	28	177	29
rect	176	29	177	30
rect	176	30	177	31
rect	176	31	177	32
rect	176	32	177	33
rect	176	33	177	34
rect	176	34	177	35
rect	176	35	177	36
rect	176	36	177	37
rect	176	37	177	38
rect	176	38	177	39
rect	176	39	177	40
rect	176	40	177	41
rect	176	41	177	42
rect	176	42	177	43
rect	176	43	177	44
rect	176	44	177	45
rect	176	45	177	46
rect	176	46	177	47
rect	176	47	177	48
rect	176	48	177	49
rect	176	49	177	50
rect	176	50	177	51
rect	176	51	177	52
rect	176	52	177	53
rect	176	53	177	54
rect	176	55	177	56
rect	176	56	177	57
rect	176	57	177	58
rect	176	59	177	60
rect	176	60	177	61
rect	176	61	177	62
rect	176	62	177	63
rect	176	63	177	64
rect	176	65	177	66
rect	176	66	177	67
rect	176	67	177	68
rect	176	68	177	69
rect	176	69	177	70
rect	176	70	177	71
rect	176	71	177	72
rect	176	72	177	73
rect	176	74	177	75
rect	176	75	177	76
rect	176	76	177	77
rect	176	77	177	78
rect	176	78	177	79
rect	176	79	177	80
rect	176	80	177	81
rect	176	81	177	82
rect	176	82	177	83
rect	176	84	177	85
rect	176	85	177	86
rect	176	86	177	87
rect	176	87	177	88
rect	176	88	177	89
rect	176	89	177	90
rect	176	90	177	91
rect	176	91	177	92
rect	176	93	177	94
rect	176	94	177	95
rect	176	95	177	96
rect	176	96	177	97
rect	176	97	177	98
rect	176	98	177	99
rect	176	99	177	100
rect	176	100	177	101
rect	176	101	177	102
rect	176	102	177	103
rect	176	103	177	104
rect	176	104	177	105
rect	176	105	177	106
rect	176	106	177	107
rect	176	107	177	108
rect	176	109	177	110
rect	176	110	177	111
rect	176	111	177	112
rect	176	112	177	113
rect	176	113	177	114
rect	176	114	177	115
rect	176	115	177	116
rect	176	116	177	117
rect	176	117	177	118
rect	176	118	177	119
rect	176	119	177	120
rect	176	120	177	121
rect	176	122	177	123
rect	176	123	177	124
rect	176	124	177	125
rect	176	125	177	126
rect	176	126	177	127
rect	176	127	177	128
rect	176	128	177	129
rect	176	129	177	130
rect	176	130	177	131
rect	176	131	177	132
rect	176	132	177	133
rect	176	133	177	134
rect	176	134	177	135
rect	176	135	177	136
rect	176	136	177	137
rect	176	138	177	139
rect	176	139	177	140
rect	176	140	177	141
rect	176	141	177	142
rect	176	142	177	143
rect	176	143	177	144
rect	176	144	177	145
rect	176	145	177	146
rect	176	146	177	147
rect	176	147	177	148
rect	176	148	177	149
rect	176	149	177	150
rect	176	150	177	151
rect	176	151	177	152
rect	176	152	177	153
rect	176	153	177	154
rect	176	154	177	155
rect	176	155	177	156
rect	176	156	177	157
rect	176	157	177	158
rect	176	158	177	159
rect	176	160	177	161
rect	176	161	177	162
rect	176	162	177	163
rect	176	163	177	164
rect	176	164	177	165
rect	176	165	177	166
rect	176	166	177	167
rect	176	167	177	168
rect	176	168	177	169
rect	176	169	177	170
rect	176	170	177	171
rect	176	171	177	172
rect	176	173	177	174
rect	176	174	177	175
rect	176	175	177	176
rect	176	176	177	177
rect	176	177	177	178
rect	176	178	177	179
rect	176	179	177	180
rect	176	180	177	181
rect	176	181	177	182
rect	176	182	177	183
rect	176	183	177	184
rect	176	184	177	185
rect	176	186	177	187
rect	176	187	177	188
rect	176	188	177	189
rect	176	189	177	190
rect	176	190	177	191
rect	176	191	177	192
rect	220	0	221	1
rect	220	1	221	2
rect	220	2	221	3
rect	220	3	221	4
rect	220	4	221	5
rect	220	5	221	6
rect	220	7	221	8
rect	220	8	221	9
rect	220	9	221	10
rect	220	10	221	11
rect	220	11	221	12
rect	220	12	221	13
rect	220	13	221	14
rect	220	14	221	15
rect	220	15	221	16
rect	220	16	221	17
rect	220	17	221	18
rect	220	18	221	19
rect	220	19	221	20
rect	220	20	221	21
rect	220	21	221	22
rect	220	22	221	23
rect	220	24	221	25
rect	220	25	221	26
rect	220	27	221	28
rect	220	28	221	29
rect	220	29	221	30
rect	220	30	221	31
rect	220	32	221	33
rect	220	33	221	34
rect	220	34	221	35
rect	220	35	221	36
rect	220	36	221	37
rect	220	37	221	38
rect	220	38	221	39
rect	220	39	221	40
rect	220	40	221	41
rect	220	41	221	42
rect	220	42	221	43
rect	220	43	221	44
rect	220	44	221	45
rect	220	45	221	46
rect	220	46	221	47
rect	220	47	221	48
rect	220	48	221	49
rect	220	49	221	50
rect	220	50	221	51
rect	220	51	221	52
rect	220	52	221	53
rect	220	53	221	54
rect	220	54	221	55
rect	220	55	221	56
rect	220	57	221	58
rect	220	58	221	59
rect	220	59	221	60
rect	220	60	221	61
rect	220	61	221	62
rect	220	62	221	63
rect	220	63	221	64
rect	220	64	221	65
rect	220	65	221	66
rect	220	66	221	67
rect	220	67	221	68
rect	220	68	221	69
rect	220	69	221	70
rect	220	70	221	71
rect	220	71	221	72
rect	220	72	221	73
rect	220	73	221	74
rect	220	74	221	75
rect	220	75	221	76
rect	220	76	221	77
rect	220	77	221	78
rect	220	78	221	79
rect	220	79	221	80
rect	220	80	221	81
rect	220	82	221	83
rect	220	83	221	84
rect	220	84	221	85
rect	220	85	221	86
rect	220	86	221	87
rect	220	87	221	88
rect	220	88	221	89
rect	220	89	221	90
rect	220	90	221	91
rect	220	91	221	92
rect	220	92	221	93
rect	220	93	221	94
rect	220	94	221	95
rect	220	95	221	96
rect	220	96	221	97
rect	220	98	221	99
rect	220	99	221	100
rect	220	100	221	101
rect	220	101	221	102
rect	220	102	221	103
rect	220	103	221	104
rect	220	104	221	105
rect	220	105	221	106
rect	220	106	221	107
rect	220	107	221	108
rect	220	108	221	109
rect	220	109	221	110
rect	220	111	221	112
rect	220	112	221	113
rect	220	113	221	114
rect	220	114	221	115
rect	220	115	221	116
rect	220	116	221	117
rect	220	117	221	118
rect	220	118	221	119
rect	220	119	221	120
rect	220	120	221	121
rect	220	121	221	122
rect	220	122	221	123
rect	220	123	221	124
rect	220	124	221	125
rect	220	125	221	126
rect	220	126	221	127
rect	220	127	221	128
rect	220	128	221	129
rect	220	130	221	131
rect	220	131	221	132
rect	220	132	221	133
rect	220	133	221	134
rect	220	134	221	135
rect	220	135	221	136
rect	220	136	221	137
rect	220	137	221	138
rect	220	138	221	139
rect	220	139	221	140
rect	220	140	221	141
rect	220	141	221	142
rect	220	142	221	143
rect	220	143	221	144
rect	220	144	221	145
rect	220	145	221	146
rect	220	146	221	147
rect	220	147	221	148
rect	220	149	221	150
rect	220	150	221	151
rect	220	151	221	152
rect	220	152	221	153
rect	220	153	221	154
rect	220	154	221	155
rect	220	155	221	156
rect	220	156	221	157
rect	220	157	221	158
rect	220	158	221	159
rect	220	159	221	160
rect	220	160	221	161
rect	220	161	221	162
rect	220	162	221	163
rect	220	163	221	164
rect	220	165	221	166
rect	220	166	221	167
rect	220	167	221	168
rect	220	168	221	169
rect	220	169	221	170
rect	220	170	221	171
rect	221	0	222	1
rect	221	1	222	2
rect	221	2	222	3
rect	221	3	222	4
rect	221	4	222	5
rect	221	5	222	6
rect	221	7	222	8
rect	221	8	222	9
rect	221	9	222	10
rect	221	10	222	11
rect	221	11	222	12
rect	221	12	222	13
rect	221	13	222	14
rect	221	14	222	15
rect	221	15	222	16
rect	221	16	222	17
rect	221	17	222	18
rect	221	18	222	19
rect	221	19	222	20
rect	221	20	222	21
rect	221	21	222	22
rect	221	22	222	23
rect	221	24	222	25
rect	221	25	222	26
rect	221	27	222	28
rect	221	28	222	29
rect	221	29	222	30
rect	221	30	222	31
rect	221	32	222	33
rect	221	33	222	34
rect	221	34	222	35
rect	221	35	222	36
rect	221	36	222	37
rect	221	37	222	38
rect	221	38	222	39
rect	221	39	222	40
rect	221	40	222	41
rect	221	41	222	42
rect	221	42	222	43
rect	221	43	222	44
rect	221	44	222	45
rect	221	45	222	46
rect	221	46	222	47
rect	221	47	222	48
rect	221	48	222	49
rect	221	49	222	50
rect	221	50	222	51
rect	221	51	222	52
rect	221	52	222	53
rect	221	53	222	54
rect	221	54	222	55
rect	221	55	222	56
rect	221	57	222	58
rect	221	58	222	59
rect	221	59	222	60
rect	221	60	222	61
rect	221	61	222	62
rect	221	62	222	63
rect	221	63	222	64
rect	221	64	222	65
rect	221	65	222	66
rect	221	66	222	67
rect	221	67	222	68
rect	221	68	222	69
rect	221	69	222	70
rect	221	70	222	71
rect	221	71	222	72
rect	221	72	222	73
rect	221	73	222	74
rect	221	74	222	75
rect	221	75	222	76
rect	221	76	222	77
rect	221	77	222	78
rect	221	78	222	79
rect	221	79	222	80
rect	221	80	222	81
rect	221	82	222	83
rect	221	83	222	84
rect	221	84	222	85
rect	221	85	222	86
rect	221	86	222	87
rect	221	87	222	88
rect	221	88	222	89
rect	221	89	222	90
rect	221	90	222	91
rect	221	91	222	92
rect	221	92	222	93
rect	221	93	222	94
rect	221	94	222	95
rect	221	95	222	96
rect	221	96	222	97
rect	221	98	222	99
rect	221	99	222	100
rect	221	100	222	101
rect	221	101	222	102
rect	221	102	222	103
rect	221	103	222	104
rect	221	104	222	105
rect	221	105	222	106
rect	221	106	222	107
rect	221	107	222	108
rect	221	108	222	109
rect	221	109	222	110
rect	221	111	222	112
rect	221	112	222	113
rect	221	113	222	114
rect	221	114	222	115
rect	221	115	222	116
rect	221	116	222	117
rect	221	117	222	118
rect	221	118	222	119
rect	221	119	222	120
rect	221	120	222	121
rect	221	121	222	122
rect	221	122	222	123
rect	221	123	222	124
rect	221	124	222	125
rect	221	125	222	126
rect	221	126	222	127
rect	221	127	222	128
rect	221	128	222	129
rect	221	130	222	131
rect	221	131	222	132
rect	221	132	222	133
rect	221	133	222	134
rect	221	134	222	135
rect	221	135	222	136
rect	221	136	222	137
rect	221	137	222	138
rect	221	138	222	139
rect	221	139	222	140
rect	221	140	222	141
rect	221	141	222	142
rect	221	142	222	143
rect	221	143	222	144
rect	221	144	222	145
rect	221	145	222	146
rect	221	146	222	147
rect	221	147	222	148
rect	221	149	222	150
rect	221	150	222	151
rect	221	151	222	152
rect	221	152	222	153
rect	221	153	222	154
rect	221	154	222	155
rect	221	155	222	156
rect	221	156	222	157
rect	221	157	222	158
rect	221	158	222	159
rect	221	159	222	160
rect	221	160	222	161
rect	221	161	222	162
rect	221	162	222	163
rect	221	163	222	164
rect	221	165	222	166
rect	221	166	222	167
rect	221	167	222	168
rect	221	168	222	169
rect	221	169	222	170
rect	221	170	222	171
rect	222	0	223	1
rect	222	1	223	2
rect	222	2	223	3
rect	222	3	223	4
rect	222	4	223	5
rect	222	5	223	6
rect	222	7	223	8
rect	222	8	223	9
rect	222	9	223	10
rect	222	10	223	11
rect	222	11	223	12
rect	222	12	223	13
rect	222	13	223	14
rect	222	14	223	15
rect	222	15	223	16
rect	222	16	223	17
rect	222	17	223	18
rect	222	18	223	19
rect	222	19	223	20
rect	222	20	223	21
rect	222	21	223	22
rect	222	22	223	23
rect	222	24	223	25
rect	222	25	223	26
rect	222	27	223	28
rect	222	28	223	29
rect	222	29	223	30
rect	222	30	223	31
rect	222	32	223	33
rect	222	33	223	34
rect	222	34	223	35
rect	222	35	223	36
rect	222	36	223	37
rect	222	37	223	38
rect	222	38	223	39
rect	222	39	223	40
rect	222	40	223	41
rect	222	41	223	42
rect	222	42	223	43
rect	222	43	223	44
rect	222	44	223	45
rect	222	45	223	46
rect	222	46	223	47
rect	222	47	223	48
rect	222	48	223	49
rect	222	49	223	50
rect	222	50	223	51
rect	222	51	223	52
rect	222	52	223	53
rect	222	53	223	54
rect	222	54	223	55
rect	222	55	223	56
rect	222	57	223	58
rect	222	58	223	59
rect	222	59	223	60
rect	222	60	223	61
rect	222	61	223	62
rect	222	62	223	63
rect	222	63	223	64
rect	222	64	223	65
rect	222	65	223	66
rect	222	66	223	67
rect	222	67	223	68
rect	222	68	223	69
rect	222	69	223	70
rect	222	70	223	71
rect	222	71	223	72
rect	222	72	223	73
rect	222	73	223	74
rect	222	74	223	75
rect	222	75	223	76
rect	222	76	223	77
rect	222	77	223	78
rect	222	78	223	79
rect	222	79	223	80
rect	222	80	223	81
rect	222	82	223	83
rect	222	83	223	84
rect	222	84	223	85
rect	222	85	223	86
rect	222	86	223	87
rect	222	87	223	88
rect	222	88	223	89
rect	222	89	223	90
rect	222	90	223	91
rect	222	91	223	92
rect	222	92	223	93
rect	222	93	223	94
rect	222	94	223	95
rect	222	95	223	96
rect	222	96	223	97
rect	222	98	223	99
rect	222	99	223	100
rect	222	100	223	101
rect	222	101	223	102
rect	222	102	223	103
rect	222	103	223	104
rect	222	104	223	105
rect	222	105	223	106
rect	222	106	223	107
rect	222	107	223	108
rect	222	108	223	109
rect	222	109	223	110
rect	222	111	223	112
rect	222	112	223	113
rect	222	113	223	114
rect	222	114	223	115
rect	222	115	223	116
rect	222	116	223	117
rect	222	117	223	118
rect	222	118	223	119
rect	222	119	223	120
rect	222	120	223	121
rect	222	121	223	122
rect	222	122	223	123
rect	222	123	223	124
rect	222	124	223	125
rect	222	125	223	126
rect	222	126	223	127
rect	222	127	223	128
rect	222	128	223	129
rect	222	130	223	131
rect	222	131	223	132
rect	222	132	223	133
rect	222	133	223	134
rect	222	134	223	135
rect	222	135	223	136
rect	222	136	223	137
rect	222	137	223	138
rect	222	138	223	139
rect	222	139	223	140
rect	222	140	223	141
rect	222	141	223	142
rect	222	142	223	143
rect	222	143	223	144
rect	222	144	223	145
rect	222	145	223	146
rect	222	146	223	147
rect	222	147	223	148
rect	222	149	223	150
rect	222	150	223	151
rect	222	151	223	152
rect	222	152	223	153
rect	222	153	223	154
rect	222	154	223	155
rect	222	155	223	156
rect	222	156	223	157
rect	222	157	223	158
rect	222	158	223	159
rect	222	159	223	160
rect	222	160	223	161
rect	222	161	223	162
rect	222	162	223	163
rect	222	163	223	164
rect	222	165	223	166
rect	222	166	223	167
rect	222	167	223	168
rect	222	168	223	169
rect	222	169	223	170
rect	222	170	223	171
rect	223	0	224	1
rect	223	1	224	2
rect	223	2	224	3
rect	223	3	224	4
rect	223	4	224	5
rect	223	5	224	6
rect	223	7	224	8
rect	223	8	224	9
rect	223	9	224	10
rect	223	10	224	11
rect	223	11	224	12
rect	223	12	224	13
rect	223	13	224	14
rect	223	14	224	15
rect	223	15	224	16
rect	223	16	224	17
rect	223	17	224	18
rect	223	18	224	19
rect	223	19	224	20
rect	223	20	224	21
rect	223	21	224	22
rect	223	22	224	23
rect	223	24	224	25
rect	223	25	224	26
rect	223	27	224	28
rect	223	28	224	29
rect	223	29	224	30
rect	223	30	224	31
rect	223	32	224	33
rect	223	33	224	34
rect	223	34	224	35
rect	223	35	224	36
rect	223	36	224	37
rect	223	37	224	38
rect	223	38	224	39
rect	223	39	224	40
rect	223	40	224	41
rect	223	41	224	42
rect	223	42	224	43
rect	223	43	224	44
rect	223	44	224	45
rect	223	45	224	46
rect	223	46	224	47
rect	223	47	224	48
rect	223	48	224	49
rect	223	49	224	50
rect	223	50	224	51
rect	223	51	224	52
rect	223	52	224	53
rect	223	53	224	54
rect	223	54	224	55
rect	223	55	224	56
rect	223	57	224	58
rect	223	58	224	59
rect	223	59	224	60
rect	223	60	224	61
rect	223	61	224	62
rect	223	62	224	63
rect	223	63	224	64
rect	223	64	224	65
rect	223	65	224	66
rect	223	66	224	67
rect	223	67	224	68
rect	223	68	224	69
rect	223	69	224	70
rect	223	70	224	71
rect	223	71	224	72
rect	223	72	224	73
rect	223	73	224	74
rect	223	74	224	75
rect	223	75	224	76
rect	223	76	224	77
rect	223	77	224	78
rect	223	78	224	79
rect	223	79	224	80
rect	223	80	224	81
rect	223	82	224	83
rect	223	83	224	84
rect	223	84	224	85
rect	223	85	224	86
rect	223	86	224	87
rect	223	87	224	88
rect	223	88	224	89
rect	223	89	224	90
rect	223	90	224	91
rect	223	91	224	92
rect	223	92	224	93
rect	223	93	224	94
rect	223	94	224	95
rect	223	95	224	96
rect	223	96	224	97
rect	223	98	224	99
rect	223	99	224	100
rect	223	100	224	101
rect	223	101	224	102
rect	223	102	224	103
rect	223	103	224	104
rect	223	104	224	105
rect	223	105	224	106
rect	223	106	224	107
rect	223	107	224	108
rect	223	108	224	109
rect	223	109	224	110
rect	223	111	224	112
rect	223	112	224	113
rect	223	113	224	114
rect	223	114	224	115
rect	223	115	224	116
rect	223	116	224	117
rect	223	117	224	118
rect	223	118	224	119
rect	223	119	224	120
rect	223	120	224	121
rect	223	121	224	122
rect	223	122	224	123
rect	223	123	224	124
rect	223	124	224	125
rect	223	125	224	126
rect	223	126	224	127
rect	223	127	224	128
rect	223	128	224	129
rect	223	130	224	131
rect	223	131	224	132
rect	223	132	224	133
rect	223	133	224	134
rect	223	134	224	135
rect	223	135	224	136
rect	223	136	224	137
rect	223	137	224	138
rect	223	138	224	139
rect	223	139	224	140
rect	223	140	224	141
rect	223	141	224	142
rect	223	142	224	143
rect	223	143	224	144
rect	223	144	224	145
rect	223	145	224	146
rect	223	146	224	147
rect	223	147	224	148
rect	223	149	224	150
rect	223	150	224	151
rect	223	151	224	152
rect	223	152	224	153
rect	223	153	224	154
rect	223	154	224	155
rect	223	155	224	156
rect	223	156	224	157
rect	223	157	224	158
rect	223	158	224	159
rect	223	159	224	160
rect	223	160	224	161
rect	223	161	224	162
rect	223	162	224	163
rect	223	163	224	164
rect	223	165	224	166
rect	223	166	224	167
rect	223	167	224	168
rect	223	168	224	169
rect	223	169	224	170
rect	223	170	224	171
rect	224	0	225	1
rect	224	1	225	2
rect	224	2	225	3
rect	224	3	225	4
rect	224	4	225	5
rect	224	5	225	6
rect	224	7	225	8
rect	224	8	225	9
rect	224	9	225	10
rect	224	10	225	11
rect	224	11	225	12
rect	224	12	225	13
rect	224	13	225	14
rect	224	14	225	15
rect	224	15	225	16
rect	224	16	225	17
rect	224	17	225	18
rect	224	18	225	19
rect	224	19	225	20
rect	224	20	225	21
rect	224	21	225	22
rect	224	22	225	23
rect	224	24	225	25
rect	224	25	225	26
rect	224	27	225	28
rect	224	28	225	29
rect	224	29	225	30
rect	224	30	225	31
rect	224	32	225	33
rect	224	33	225	34
rect	224	34	225	35
rect	224	35	225	36
rect	224	36	225	37
rect	224	37	225	38
rect	224	38	225	39
rect	224	39	225	40
rect	224	40	225	41
rect	224	41	225	42
rect	224	42	225	43
rect	224	43	225	44
rect	224	44	225	45
rect	224	45	225	46
rect	224	46	225	47
rect	224	47	225	48
rect	224	48	225	49
rect	224	49	225	50
rect	224	50	225	51
rect	224	51	225	52
rect	224	52	225	53
rect	224	53	225	54
rect	224	54	225	55
rect	224	55	225	56
rect	224	57	225	58
rect	224	58	225	59
rect	224	59	225	60
rect	224	60	225	61
rect	224	61	225	62
rect	224	62	225	63
rect	224	63	225	64
rect	224	64	225	65
rect	224	65	225	66
rect	224	66	225	67
rect	224	67	225	68
rect	224	68	225	69
rect	224	69	225	70
rect	224	70	225	71
rect	224	71	225	72
rect	224	72	225	73
rect	224	73	225	74
rect	224	74	225	75
rect	224	75	225	76
rect	224	76	225	77
rect	224	77	225	78
rect	224	78	225	79
rect	224	79	225	80
rect	224	80	225	81
rect	224	82	225	83
rect	224	83	225	84
rect	224	84	225	85
rect	224	85	225	86
rect	224	86	225	87
rect	224	87	225	88
rect	224	88	225	89
rect	224	89	225	90
rect	224	90	225	91
rect	224	91	225	92
rect	224	92	225	93
rect	224	93	225	94
rect	224	94	225	95
rect	224	95	225	96
rect	224	96	225	97
rect	224	98	225	99
rect	224	99	225	100
rect	224	100	225	101
rect	224	101	225	102
rect	224	102	225	103
rect	224	103	225	104
rect	224	104	225	105
rect	224	105	225	106
rect	224	106	225	107
rect	224	107	225	108
rect	224	108	225	109
rect	224	109	225	110
rect	224	111	225	112
rect	224	112	225	113
rect	224	113	225	114
rect	224	114	225	115
rect	224	115	225	116
rect	224	116	225	117
rect	224	117	225	118
rect	224	118	225	119
rect	224	119	225	120
rect	224	120	225	121
rect	224	121	225	122
rect	224	122	225	123
rect	224	123	225	124
rect	224	124	225	125
rect	224	125	225	126
rect	224	126	225	127
rect	224	127	225	128
rect	224	128	225	129
rect	224	130	225	131
rect	224	131	225	132
rect	224	132	225	133
rect	224	133	225	134
rect	224	134	225	135
rect	224	135	225	136
rect	224	136	225	137
rect	224	137	225	138
rect	224	138	225	139
rect	224	139	225	140
rect	224	140	225	141
rect	224	141	225	142
rect	224	142	225	143
rect	224	143	225	144
rect	224	144	225	145
rect	224	145	225	146
rect	224	146	225	147
rect	224	147	225	148
rect	224	149	225	150
rect	224	150	225	151
rect	224	151	225	152
rect	224	152	225	153
rect	224	153	225	154
rect	224	154	225	155
rect	224	155	225	156
rect	224	156	225	157
rect	224	157	225	158
rect	224	158	225	159
rect	224	159	225	160
rect	224	160	225	161
rect	224	161	225	162
rect	224	162	225	163
rect	224	163	225	164
rect	224	165	225	166
rect	224	166	225	167
rect	224	167	225	168
rect	224	168	225	169
rect	224	169	225	170
rect	224	170	225	171
rect	225	0	226	1
rect	225	1	226	2
rect	225	2	226	3
rect	225	3	226	4
rect	225	4	226	5
rect	225	5	226	6
rect	225	7	226	8
rect	225	8	226	9
rect	225	9	226	10
rect	225	10	226	11
rect	225	11	226	12
rect	225	12	226	13
rect	225	13	226	14
rect	225	14	226	15
rect	225	15	226	16
rect	225	16	226	17
rect	225	17	226	18
rect	225	18	226	19
rect	225	19	226	20
rect	225	20	226	21
rect	225	21	226	22
rect	225	22	226	23
rect	225	24	226	25
rect	225	25	226	26
rect	225	27	226	28
rect	225	28	226	29
rect	225	29	226	30
rect	225	30	226	31
rect	225	32	226	33
rect	225	33	226	34
rect	225	34	226	35
rect	225	35	226	36
rect	225	36	226	37
rect	225	37	226	38
rect	225	38	226	39
rect	225	39	226	40
rect	225	40	226	41
rect	225	41	226	42
rect	225	42	226	43
rect	225	43	226	44
rect	225	44	226	45
rect	225	45	226	46
rect	225	46	226	47
rect	225	47	226	48
rect	225	48	226	49
rect	225	49	226	50
rect	225	50	226	51
rect	225	51	226	52
rect	225	52	226	53
rect	225	53	226	54
rect	225	54	226	55
rect	225	55	226	56
rect	225	57	226	58
rect	225	58	226	59
rect	225	59	226	60
rect	225	60	226	61
rect	225	61	226	62
rect	225	62	226	63
rect	225	63	226	64
rect	225	64	226	65
rect	225	65	226	66
rect	225	66	226	67
rect	225	67	226	68
rect	225	68	226	69
rect	225	69	226	70
rect	225	70	226	71
rect	225	71	226	72
rect	225	72	226	73
rect	225	73	226	74
rect	225	74	226	75
rect	225	75	226	76
rect	225	76	226	77
rect	225	77	226	78
rect	225	78	226	79
rect	225	79	226	80
rect	225	80	226	81
rect	225	82	226	83
rect	225	83	226	84
rect	225	84	226	85
rect	225	85	226	86
rect	225	86	226	87
rect	225	87	226	88
rect	225	88	226	89
rect	225	89	226	90
rect	225	90	226	91
rect	225	91	226	92
rect	225	92	226	93
rect	225	93	226	94
rect	225	94	226	95
rect	225	95	226	96
rect	225	96	226	97
rect	225	98	226	99
rect	225	99	226	100
rect	225	100	226	101
rect	225	101	226	102
rect	225	102	226	103
rect	225	103	226	104
rect	225	104	226	105
rect	225	105	226	106
rect	225	106	226	107
rect	225	107	226	108
rect	225	108	226	109
rect	225	109	226	110
rect	225	111	226	112
rect	225	112	226	113
rect	225	113	226	114
rect	225	114	226	115
rect	225	115	226	116
rect	225	116	226	117
rect	225	117	226	118
rect	225	118	226	119
rect	225	119	226	120
rect	225	120	226	121
rect	225	121	226	122
rect	225	122	226	123
rect	225	123	226	124
rect	225	124	226	125
rect	225	125	226	126
rect	225	126	226	127
rect	225	127	226	128
rect	225	128	226	129
rect	225	130	226	131
rect	225	131	226	132
rect	225	132	226	133
rect	225	133	226	134
rect	225	134	226	135
rect	225	135	226	136
rect	225	136	226	137
rect	225	137	226	138
rect	225	138	226	139
rect	225	139	226	140
rect	225	140	226	141
rect	225	141	226	142
rect	225	142	226	143
rect	225	143	226	144
rect	225	144	226	145
rect	225	145	226	146
rect	225	146	226	147
rect	225	147	226	148
rect	225	149	226	150
rect	225	150	226	151
rect	225	151	226	152
rect	225	152	226	153
rect	225	153	226	154
rect	225	154	226	155
rect	225	155	226	156
rect	225	156	226	157
rect	225	157	226	158
rect	225	158	226	159
rect	225	159	226	160
rect	225	160	226	161
rect	225	161	226	162
rect	225	162	226	163
rect	225	163	226	164
rect	225	165	226	166
rect	225	166	226	167
rect	225	167	226	168
rect	225	168	226	169
rect	225	169	226	170
rect	225	170	226	171
rect	261	0	262	1
rect	261	1	262	2
rect	261	2	262	3
rect	261	3	262	4
rect	261	4	262	5
rect	261	5	262	6
rect	261	6	262	7
rect	261	7	262	8
rect	261	8	262	9
rect	261	10	262	11
rect	261	11	262	12
rect	261	12	262	13
rect	261	13	262	14
rect	261	14	262	15
rect	261	15	262	16
rect	261	16	262	17
rect	261	17	262	18
rect	261	18	262	19
rect	261	19	262	20
rect	261	20	262	21
rect	261	21	262	22
rect	261	22	262	23
rect	261	23	262	24
rect	261	24	262	25
rect	261	25	262	26
rect	261	26	262	27
rect	261	27	262	28
rect	261	29	262	30
rect	261	30	262	31
rect	261	31	262	32
rect	261	32	262	33
rect	261	33	262	34
rect	261	34	262	35
rect	261	35	262	36
rect	261	36	262	37
rect	261	37	262	38
rect	261	38	262	39
rect	261	39	262	40
rect	261	40	262	41
rect	261	41	262	42
rect	261	42	262	43
rect	261	43	262	44
rect	261	44	262	45
rect	261	45	262	46
rect	261	46	262	47
rect	261	47	262	48
rect	261	48	262	49
rect	261	49	262	50
rect	261	50	262	51
rect	261	51	262	52
rect	261	52	262	53
rect	261	53	262	54
rect	261	54	262	55
rect	261	55	262	56
rect	261	56	262	57
rect	261	57	262	58
rect	261	58	262	59
rect	261	59	262	60
rect	261	60	262	61
rect	261	61	262	62
rect	261	63	262	64
rect	261	64	262	65
rect	261	65	262	66
rect	261	66	262	67
rect	261	67	262	68
rect	261	68	262	69
rect	261	69	262	70
rect	261	70	262	71
rect	261	71	262	72
rect	261	72	262	73
rect	261	73	262	74
rect	261	74	262	75
rect	261	75	262	76
rect	261	76	262	77
rect	261	77	262	78
rect	261	79	262	80
rect	261	80	262	81
rect	261	81	262	82
rect	261	82	262	83
rect	261	83	262	84
rect	261	84	262	85
rect	261	85	262	86
rect	261	86	262	87
rect	261	87	262	88
rect	261	88	262	89
rect	261	89	262	90
rect	261	90	262	91
rect	261	92	262	93
rect	261	93	262	94
rect	261	94	262	95
rect	261	95	262	96
rect	261	96	262	97
rect	261	97	262	98
rect	261	98	262	99
rect	261	99	262	100
rect	261	100	262	101
rect	261	101	262	102
rect	261	102	262	103
rect	261	103	262	104
rect	261	105	262	106
rect	261	106	262	107
rect	261	107	262	108
rect	261	108	262	109
rect	261	109	262	110
rect	261	110	262	111
rect	261	111	262	112
rect	261	112	262	113
rect	261	113	262	114
rect	261	115	262	116
rect	261	116	262	117
rect	261	117	262	118
rect	261	118	262	119
rect	261	119	262	120
rect	261	120	262	121
rect	261	122	262	123
rect	261	123	262	124
rect	261	124	262	125
rect	261	125	262	126
rect	261	126	262	127
rect	261	127	262	128
rect	261	128	262	129
rect	261	129	262	130
rect	261	130	262	131
rect	261	132	262	133
rect	261	133	262	134
rect	261	134	262	135
rect	261	135	262	136
rect	261	136	262	137
rect	261	137	262	138
rect	261	138	262	139
rect	261	139	262	140
rect	261	140	262	141
rect	262	0	263	1
rect	262	1	263	2
rect	262	2	263	3
rect	262	3	263	4
rect	262	4	263	5
rect	262	5	263	6
rect	262	6	263	7
rect	262	7	263	8
rect	262	8	263	9
rect	262	10	263	11
rect	262	11	263	12
rect	262	12	263	13
rect	262	13	263	14
rect	262	14	263	15
rect	262	15	263	16
rect	262	16	263	17
rect	262	17	263	18
rect	262	18	263	19
rect	262	19	263	20
rect	262	20	263	21
rect	262	21	263	22
rect	262	22	263	23
rect	262	23	263	24
rect	262	24	263	25
rect	262	25	263	26
rect	262	26	263	27
rect	262	27	263	28
rect	262	29	263	30
rect	262	30	263	31
rect	262	31	263	32
rect	262	32	263	33
rect	262	33	263	34
rect	262	34	263	35
rect	262	35	263	36
rect	262	36	263	37
rect	262	37	263	38
rect	262	38	263	39
rect	262	39	263	40
rect	262	40	263	41
rect	262	41	263	42
rect	262	42	263	43
rect	262	43	263	44
rect	262	44	263	45
rect	262	45	263	46
rect	262	46	263	47
rect	262	47	263	48
rect	262	48	263	49
rect	262	49	263	50
rect	262	50	263	51
rect	262	51	263	52
rect	262	52	263	53
rect	262	53	263	54
rect	262	54	263	55
rect	262	55	263	56
rect	262	56	263	57
rect	262	57	263	58
rect	262	58	263	59
rect	262	59	263	60
rect	262	60	263	61
rect	262	61	263	62
rect	262	63	263	64
rect	262	64	263	65
rect	262	65	263	66
rect	262	66	263	67
rect	262	67	263	68
rect	262	68	263	69
rect	262	69	263	70
rect	262	70	263	71
rect	262	71	263	72
rect	262	72	263	73
rect	262	73	263	74
rect	262	74	263	75
rect	262	75	263	76
rect	262	76	263	77
rect	262	77	263	78
rect	262	79	263	80
rect	262	80	263	81
rect	262	81	263	82
rect	262	82	263	83
rect	262	83	263	84
rect	262	84	263	85
rect	262	85	263	86
rect	262	86	263	87
rect	262	87	263	88
rect	262	88	263	89
rect	262	89	263	90
rect	262	90	263	91
rect	262	92	263	93
rect	262	93	263	94
rect	262	94	263	95
rect	262	95	263	96
rect	262	96	263	97
rect	262	97	263	98
rect	262	98	263	99
rect	262	99	263	100
rect	262	100	263	101
rect	262	101	263	102
rect	262	102	263	103
rect	262	103	263	104
rect	262	105	263	106
rect	262	106	263	107
rect	262	107	263	108
rect	262	108	263	109
rect	262	109	263	110
rect	262	110	263	111
rect	262	111	263	112
rect	262	112	263	113
rect	262	113	263	114
rect	262	115	263	116
rect	262	116	263	117
rect	262	117	263	118
rect	262	118	263	119
rect	262	119	263	120
rect	262	120	263	121
rect	262	122	263	123
rect	262	123	263	124
rect	262	124	263	125
rect	262	125	263	126
rect	262	126	263	127
rect	262	127	263	128
rect	262	128	263	129
rect	262	129	263	130
rect	262	130	263	131
rect	262	132	263	133
rect	262	133	263	134
rect	262	134	263	135
rect	262	135	263	136
rect	262	136	263	137
rect	262	137	263	138
rect	262	138	263	139
rect	262	139	263	140
rect	262	140	263	141
rect	263	0	264	1
rect	263	1	264	2
rect	263	2	264	3
rect	263	3	264	4
rect	263	4	264	5
rect	263	5	264	6
rect	263	6	264	7
rect	263	7	264	8
rect	263	8	264	9
rect	263	10	264	11
rect	263	11	264	12
rect	263	12	264	13
rect	263	13	264	14
rect	263	14	264	15
rect	263	15	264	16
rect	263	16	264	17
rect	263	17	264	18
rect	263	18	264	19
rect	263	19	264	20
rect	263	20	264	21
rect	263	21	264	22
rect	263	22	264	23
rect	263	23	264	24
rect	263	24	264	25
rect	263	25	264	26
rect	263	26	264	27
rect	263	27	264	28
rect	263	29	264	30
rect	263	30	264	31
rect	263	31	264	32
rect	263	32	264	33
rect	263	33	264	34
rect	263	34	264	35
rect	263	35	264	36
rect	263	36	264	37
rect	263	37	264	38
rect	263	38	264	39
rect	263	39	264	40
rect	263	40	264	41
rect	263	41	264	42
rect	263	42	264	43
rect	263	43	264	44
rect	263	44	264	45
rect	263	45	264	46
rect	263	46	264	47
rect	263	47	264	48
rect	263	48	264	49
rect	263	49	264	50
rect	263	50	264	51
rect	263	51	264	52
rect	263	52	264	53
rect	263	53	264	54
rect	263	54	264	55
rect	263	55	264	56
rect	263	56	264	57
rect	263	57	264	58
rect	263	58	264	59
rect	263	59	264	60
rect	263	60	264	61
rect	263	61	264	62
rect	263	63	264	64
rect	263	64	264	65
rect	263	65	264	66
rect	263	66	264	67
rect	263	67	264	68
rect	263	68	264	69
rect	263	69	264	70
rect	263	70	264	71
rect	263	71	264	72
rect	263	72	264	73
rect	263	73	264	74
rect	263	74	264	75
rect	263	75	264	76
rect	263	76	264	77
rect	263	77	264	78
rect	263	79	264	80
rect	263	80	264	81
rect	263	81	264	82
rect	263	82	264	83
rect	263	83	264	84
rect	263	84	264	85
rect	263	85	264	86
rect	263	86	264	87
rect	263	87	264	88
rect	263	88	264	89
rect	263	89	264	90
rect	263	90	264	91
rect	263	92	264	93
rect	263	93	264	94
rect	263	94	264	95
rect	263	95	264	96
rect	263	96	264	97
rect	263	97	264	98
rect	263	98	264	99
rect	263	99	264	100
rect	263	100	264	101
rect	263	101	264	102
rect	263	102	264	103
rect	263	103	264	104
rect	263	105	264	106
rect	263	106	264	107
rect	263	107	264	108
rect	263	108	264	109
rect	263	109	264	110
rect	263	110	264	111
rect	263	111	264	112
rect	263	112	264	113
rect	263	113	264	114
rect	263	115	264	116
rect	263	116	264	117
rect	263	117	264	118
rect	263	118	264	119
rect	263	119	264	120
rect	263	120	264	121
rect	263	122	264	123
rect	263	123	264	124
rect	263	124	264	125
rect	263	125	264	126
rect	263	126	264	127
rect	263	127	264	128
rect	263	128	264	129
rect	263	129	264	130
rect	263	130	264	131
rect	263	132	264	133
rect	263	133	264	134
rect	263	134	264	135
rect	263	135	264	136
rect	263	136	264	137
rect	263	137	264	138
rect	263	138	264	139
rect	263	139	264	140
rect	263	140	264	141
rect	264	0	265	1
rect	264	1	265	2
rect	264	2	265	3
rect	264	3	265	4
rect	264	4	265	5
rect	264	5	265	6
rect	264	6	265	7
rect	264	7	265	8
rect	264	8	265	9
rect	264	10	265	11
rect	264	11	265	12
rect	264	12	265	13
rect	264	13	265	14
rect	264	14	265	15
rect	264	15	265	16
rect	264	16	265	17
rect	264	17	265	18
rect	264	18	265	19
rect	264	19	265	20
rect	264	20	265	21
rect	264	21	265	22
rect	264	22	265	23
rect	264	23	265	24
rect	264	24	265	25
rect	264	25	265	26
rect	264	26	265	27
rect	264	27	265	28
rect	264	29	265	30
rect	264	30	265	31
rect	264	31	265	32
rect	264	32	265	33
rect	264	33	265	34
rect	264	34	265	35
rect	264	35	265	36
rect	264	36	265	37
rect	264	37	265	38
rect	264	38	265	39
rect	264	39	265	40
rect	264	40	265	41
rect	264	41	265	42
rect	264	42	265	43
rect	264	43	265	44
rect	264	44	265	45
rect	264	45	265	46
rect	264	46	265	47
rect	264	47	265	48
rect	264	48	265	49
rect	264	49	265	50
rect	264	50	265	51
rect	264	51	265	52
rect	264	52	265	53
rect	264	53	265	54
rect	264	54	265	55
rect	264	55	265	56
rect	264	56	265	57
rect	264	57	265	58
rect	264	58	265	59
rect	264	59	265	60
rect	264	60	265	61
rect	264	61	265	62
rect	264	63	265	64
rect	264	64	265	65
rect	264	65	265	66
rect	264	66	265	67
rect	264	67	265	68
rect	264	68	265	69
rect	264	69	265	70
rect	264	70	265	71
rect	264	71	265	72
rect	264	72	265	73
rect	264	73	265	74
rect	264	74	265	75
rect	264	75	265	76
rect	264	76	265	77
rect	264	77	265	78
rect	264	79	265	80
rect	264	80	265	81
rect	264	81	265	82
rect	264	82	265	83
rect	264	83	265	84
rect	264	84	265	85
rect	264	85	265	86
rect	264	86	265	87
rect	264	87	265	88
rect	264	88	265	89
rect	264	89	265	90
rect	264	90	265	91
rect	264	92	265	93
rect	264	93	265	94
rect	264	94	265	95
rect	264	95	265	96
rect	264	96	265	97
rect	264	97	265	98
rect	264	98	265	99
rect	264	99	265	100
rect	264	100	265	101
rect	264	101	265	102
rect	264	102	265	103
rect	264	103	265	104
rect	264	105	265	106
rect	264	106	265	107
rect	264	107	265	108
rect	264	108	265	109
rect	264	109	265	110
rect	264	110	265	111
rect	264	111	265	112
rect	264	112	265	113
rect	264	113	265	114
rect	264	115	265	116
rect	264	116	265	117
rect	264	117	265	118
rect	264	118	265	119
rect	264	119	265	120
rect	264	120	265	121
rect	264	122	265	123
rect	264	123	265	124
rect	264	124	265	125
rect	264	125	265	126
rect	264	126	265	127
rect	264	127	265	128
rect	264	128	265	129
rect	264	129	265	130
rect	264	130	265	131
rect	264	132	265	133
rect	264	133	265	134
rect	264	134	265	135
rect	264	135	265	136
rect	264	136	265	137
rect	264	137	265	138
rect	264	138	265	139
rect	264	139	265	140
rect	264	140	265	141
rect	265	0	266	1
rect	265	1	266	2
rect	265	2	266	3
rect	265	3	266	4
rect	265	4	266	5
rect	265	5	266	6
rect	265	6	266	7
rect	265	7	266	8
rect	265	8	266	9
rect	265	10	266	11
rect	265	11	266	12
rect	265	12	266	13
rect	265	13	266	14
rect	265	14	266	15
rect	265	15	266	16
rect	265	16	266	17
rect	265	17	266	18
rect	265	18	266	19
rect	265	19	266	20
rect	265	20	266	21
rect	265	21	266	22
rect	265	22	266	23
rect	265	23	266	24
rect	265	24	266	25
rect	265	25	266	26
rect	265	26	266	27
rect	265	27	266	28
rect	265	29	266	30
rect	265	30	266	31
rect	265	31	266	32
rect	265	32	266	33
rect	265	33	266	34
rect	265	34	266	35
rect	265	35	266	36
rect	265	36	266	37
rect	265	37	266	38
rect	265	38	266	39
rect	265	39	266	40
rect	265	40	266	41
rect	265	41	266	42
rect	265	42	266	43
rect	265	43	266	44
rect	265	44	266	45
rect	265	45	266	46
rect	265	46	266	47
rect	265	47	266	48
rect	265	48	266	49
rect	265	49	266	50
rect	265	50	266	51
rect	265	51	266	52
rect	265	52	266	53
rect	265	53	266	54
rect	265	54	266	55
rect	265	55	266	56
rect	265	56	266	57
rect	265	57	266	58
rect	265	58	266	59
rect	265	59	266	60
rect	265	60	266	61
rect	265	61	266	62
rect	265	63	266	64
rect	265	64	266	65
rect	265	65	266	66
rect	265	66	266	67
rect	265	67	266	68
rect	265	68	266	69
rect	265	69	266	70
rect	265	70	266	71
rect	265	71	266	72
rect	265	72	266	73
rect	265	73	266	74
rect	265	74	266	75
rect	265	75	266	76
rect	265	76	266	77
rect	265	77	266	78
rect	265	79	266	80
rect	265	80	266	81
rect	265	81	266	82
rect	265	82	266	83
rect	265	83	266	84
rect	265	84	266	85
rect	265	85	266	86
rect	265	86	266	87
rect	265	87	266	88
rect	265	88	266	89
rect	265	89	266	90
rect	265	90	266	91
rect	265	92	266	93
rect	265	93	266	94
rect	265	94	266	95
rect	265	95	266	96
rect	265	96	266	97
rect	265	97	266	98
rect	265	98	266	99
rect	265	99	266	100
rect	265	100	266	101
rect	265	101	266	102
rect	265	102	266	103
rect	265	103	266	104
rect	265	105	266	106
rect	265	106	266	107
rect	265	107	266	108
rect	265	108	266	109
rect	265	109	266	110
rect	265	110	266	111
rect	265	111	266	112
rect	265	112	266	113
rect	265	113	266	114
rect	265	115	266	116
rect	265	116	266	117
rect	265	117	266	118
rect	265	118	266	119
rect	265	119	266	120
rect	265	120	266	121
rect	265	122	266	123
rect	265	123	266	124
rect	265	124	266	125
rect	265	125	266	126
rect	265	126	266	127
rect	265	127	266	128
rect	265	128	266	129
rect	265	129	266	130
rect	265	130	266	131
rect	265	132	266	133
rect	265	133	266	134
rect	265	134	266	135
rect	265	135	266	136
rect	265	136	266	137
rect	265	137	266	138
rect	265	138	266	139
rect	265	139	266	140
rect	265	140	266	141
rect	266	0	267	1
rect	266	1	267	2
rect	266	2	267	3
rect	266	3	267	4
rect	266	4	267	5
rect	266	5	267	6
rect	266	6	267	7
rect	266	7	267	8
rect	266	8	267	9
rect	266	10	267	11
rect	266	11	267	12
rect	266	12	267	13
rect	266	13	267	14
rect	266	14	267	15
rect	266	15	267	16
rect	266	16	267	17
rect	266	17	267	18
rect	266	18	267	19
rect	266	19	267	20
rect	266	20	267	21
rect	266	21	267	22
rect	266	22	267	23
rect	266	23	267	24
rect	266	24	267	25
rect	266	25	267	26
rect	266	26	267	27
rect	266	27	267	28
rect	266	29	267	30
rect	266	30	267	31
rect	266	31	267	32
rect	266	32	267	33
rect	266	33	267	34
rect	266	34	267	35
rect	266	35	267	36
rect	266	36	267	37
rect	266	37	267	38
rect	266	38	267	39
rect	266	39	267	40
rect	266	40	267	41
rect	266	41	267	42
rect	266	42	267	43
rect	266	43	267	44
rect	266	44	267	45
rect	266	45	267	46
rect	266	46	267	47
rect	266	47	267	48
rect	266	48	267	49
rect	266	49	267	50
rect	266	50	267	51
rect	266	51	267	52
rect	266	52	267	53
rect	266	53	267	54
rect	266	54	267	55
rect	266	55	267	56
rect	266	56	267	57
rect	266	57	267	58
rect	266	58	267	59
rect	266	59	267	60
rect	266	60	267	61
rect	266	61	267	62
rect	266	63	267	64
rect	266	64	267	65
rect	266	65	267	66
rect	266	66	267	67
rect	266	67	267	68
rect	266	68	267	69
rect	266	69	267	70
rect	266	70	267	71
rect	266	71	267	72
rect	266	72	267	73
rect	266	73	267	74
rect	266	74	267	75
rect	266	75	267	76
rect	266	76	267	77
rect	266	77	267	78
rect	266	79	267	80
rect	266	80	267	81
rect	266	81	267	82
rect	266	82	267	83
rect	266	83	267	84
rect	266	84	267	85
rect	266	85	267	86
rect	266	86	267	87
rect	266	87	267	88
rect	266	88	267	89
rect	266	89	267	90
rect	266	90	267	91
rect	266	92	267	93
rect	266	93	267	94
rect	266	94	267	95
rect	266	95	267	96
rect	266	96	267	97
rect	266	97	267	98
rect	266	98	267	99
rect	266	99	267	100
rect	266	100	267	101
rect	266	101	267	102
rect	266	102	267	103
rect	266	103	267	104
rect	266	105	267	106
rect	266	106	267	107
rect	266	107	267	108
rect	266	108	267	109
rect	266	109	267	110
rect	266	110	267	111
rect	266	111	267	112
rect	266	112	267	113
rect	266	113	267	114
rect	266	115	267	116
rect	266	116	267	117
rect	266	117	267	118
rect	266	118	267	119
rect	266	119	267	120
rect	266	120	267	121
rect	266	122	267	123
rect	266	123	267	124
rect	266	124	267	125
rect	266	125	267	126
rect	266	126	267	127
rect	266	127	267	128
rect	266	128	267	129
rect	266	129	267	130
rect	266	130	267	131
rect	266	132	267	133
rect	266	133	267	134
rect	266	134	267	135
rect	266	135	267	136
rect	266	136	267	137
rect	266	137	267	138
rect	266	138	267	139
rect	266	139	267	140
rect	266	140	267	141
rect	284	0	285	1
rect	284	1	285	2
rect	284	2	285	3
rect	284	3	285	4
rect	284	4	285	5
rect	284	5	285	6
rect	284	7	285	8
rect	284	8	285	9
rect	284	9	285	10
rect	284	10	285	11
rect	284	11	285	12
rect	284	12	285	13
rect	284	13	285	14
rect	284	14	285	15
rect	284	15	285	16
rect	284	17	285	18
rect	284	18	285	19
rect	284	19	285	20
rect	284	20	285	21
rect	284	21	285	22
rect	284	22	285	23
rect	284	24	285	25
rect	284	25	285	26
rect	284	26	285	27
rect	284	27	285	28
rect	284	28	285	29
rect	284	29	285	30
rect	284	31	285	32
rect	284	32	285	33
rect	284	33	285	34
rect	284	34	285	35
rect	284	35	285	36
rect	284	36	285	37
rect	284	38	285	39
rect	284	39	285	40
rect	284	40	285	41
rect	284	41	285	42
rect	284	42	285	43
rect	284	43	285	44
rect	284	44	285	45
rect	284	45	285	46
rect	284	46	285	47
rect	284	48	285	49
rect	284	49	285	50
rect	284	50	285	51
rect	284	51	285	52
rect	284	52	285	53
rect	284	53	285	54
rect	284	54	285	55
rect	284	55	285	56
rect	284	56	285	57
rect	284	58	285	59
rect	284	59	285	60
rect	284	60	285	61
rect	284	61	285	62
rect	284	62	285	63
rect	284	63	285	64
rect	284	65	285	66
rect	284	66	285	67
rect	284	67	285	68
rect	284	68	285	69
rect	284	69	285	70
rect	284	70	285	71
rect	284	72	285	73
rect	284	73	285	74
rect	284	74	285	75
rect	284	75	285	76
rect	284	76	285	77
rect	284	77	285	78
rect	285	0	286	1
rect	285	1	286	2
rect	285	2	286	3
rect	285	3	286	4
rect	285	4	286	5
rect	285	5	286	6
rect	285	7	286	8
rect	285	8	286	9
rect	285	9	286	10
rect	285	10	286	11
rect	285	11	286	12
rect	285	12	286	13
rect	285	13	286	14
rect	285	14	286	15
rect	285	15	286	16
rect	285	17	286	18
rect	285	18	286	19
rect	285	19	286	20
rect	285	20	286	21
rect	285	21	286	22
rect	285	22	286	23
rect	285	24	286	25
rect	285	25	286	26
rect	285	26	286	27
rect	285	27	286	28
rect	285	28	286	29
rect	285	29	286	30
rect	285	31	286	32
rect	285	32	286	33
rect	285	33	286	34
rect	285	34	286	35
rect	285	35	286	36
rect	285	36	286	37
rect	285	38	286	39
rect	285	39	286	40
rect	285	40	286	41
rect	285	41	286	42
rect	285	42	286	43
rect	285	43	286	44
rect	285	44	286	45
rect	285	45	286	46
rect	285	46	286	47
rect	285	48	286	49
rect	285	49	286	50
rect	285	50	286	51
rect	285	51	286	52
rect	285	52	286	53
rect	285	53	286	54
rect	285	54	286	55
rect	285	55	286	56
rect	285	56	286	57
rect	285	58	286	59
rect	285	59	286	60
rect	285	60	286	61
rect	285	61	286	62
rect	285	62	286	63
rect	285	63	286	64
rect	285	65	286	66
rect	285	66	286	67
rect	285	67	286	68
rect	285	68	286	69
rect	285	69	286	70
rect	285	70	286	71
rect	285	72	286	73
rect	285	73	286	74
rect	285	74	286	75
rect	285	75	286	76
rect	285	76	286	77
rect	285	77	286	78
rect	286	0	287	1
rect	286	1	287	2
rect	286	2	287	3
rect	286	3	287	4
rect	286	4	287	5
rect	286	5	287	6
rect	286	7	287	8
rect	286	8	287	9
rect	286	9	287	10
rect	286	10	287	11
rect	286	11	287	12
rect	286	12	287	13
rect	286	13	287	14
rect	286	14	287	15
rect	286	15	287	16
rect	286	17	287	18
rect	286	18	287	19
rect	286	19	287	20
rect	286	20	287	21
rect	286	21	287	22
rect	286	22	287	23
rect	286	24	287	25
rect	286	25	287	26
rect	286	26	287	27
rect	286	27	287	28
rect	286	28	287	29
rect	286	29	287	30
rect	286	31	287	32
rect	286	32	287	33
rect	286	33	287	34
rect	286	34	287	35
rect	286	35	287	36
rect	286	36	287	37
rect	286	38	287	39
rect	286	39	287	40
rect	286	40	287	41
rect	286	41	287	42
rect	286	42	287	43
rect	286	43	287	44
rect	286	44	287	45
rect	286	45	287	46
rect	286	46	287	47
rect	286	48	287	49
rect	286	49	287	50
rect	286	50	287	51
rect	286	51	287	52
rect	286	52	287	53
rect	286	53	287	54
rect	286	54	287	55
rect	286	55	287	56
rect	286	56	287	57
rect	286	58	287	59
rect	286	59	287	60
rect	286	60	287	61
rect	286	61	287	62
rect	286	62	287	63
rect	286	63	287	64
rect	286	65	287	66
rect	286	66	287	67
rect	286	67	287	68
rect	286	68	287	69
rect	286	69	287	70
rect	286	70	287	71
rect	286	72	287	73
rect	286	73	287	74
rect	286	74	287	75
rect	286	75	287	76
rect	286	76	287	77
rect	286	77	287	78
rect	287	0	288	1
rect	287	1	288	2
rect	287	2	288	3
rect	287	3	288	4
rect	287	4	288	5
rect	287	5	288	6
rect	287	7	288	8
rect	287	8	288	9
rect	287	9	288	10
rect	287	10	288	11
rect	287	11	288	12
rect	287	12	288	13
rect	287	13	288	14
rect	287	14	288	15
rect	287	15	288	16
rect	287	17	288	18
rect	287	18	288	19
rect	287	19	288	20
rect	287	20	288	21
rect	287	21	288	22
rect	287	22	288	23
rect	287	24	288	25
rect	287	25	288	26
rect	287	26	288	27
rect	287	27	288	28
rect	287	28	288	29
rect	287	29	288	30
rect	287	31	288	32
rect	287	32	288	33
rect	287	33	288	34
rect	287	34	288	35
rect	287	35	288	36
rect	287	36	288	37
rect	287	38	288	39
rect	287	39	288	40
rect	287	40	288	41
rect	287	41	288	42
rect	287	42	288	43
rect	287	43	288	44
rect	287	44	288	45
rect	287	45	288	46
rect	287	46	288	47
rect	287	48	288	49
rect	287	49	288	50
rect	287	50	288	51
rect	287	51	288	52
rect	287	52	288	53
rect	287	53	288	54
rect	287	54	288	55
rect	287	55	288	56
rect	287	56	288	57
rect	287	58	288	59
rect	287	59	288	60
rect	287	60	288	61
rect	287	61	288	62
rect	287	62	288	63
rect	287	63	288	64
rect	287	65	288	66
rect	287	66	288	67
rect	287	67	288	68
rect	287	68	288	69
rect	287	69	288	70
rect	287	70	288	71
rect	287	72	288	73
rect	287	73	288	74
rect	287	74	288	75
rect	287	75	288	76
rect	287	76	288	77
rect	287	77	288	78
rect	288	0	289	1
rect	288	1	289	2
rect	288	2	289	3
rect	288	3	289	4
rect	288	4	289	5
rect	288	5	289	6
rect	288	7	289	8
rect	288	8	289	9
rect	288	9	289	10
rect	288	10	289	11
rect	288	11	289	12
rect	288	12	289	13
rect	288	13	289	14
rect	288	14	289	15
rect	288	15	289	16
rect	288	17	289	18
rect	288	18	289	19
rect	288	19	289	20
rect	288	20	289	21
rect	288	21	289	22
rect	288	22	289	23
rect	288	24	289	25
rect	288	25	289	26
rect	288	26	289	27
rect	288	27	289	28
rect	288	28	289	29
rect	288	29	289	30
rect	288	31	289	32
rect	288	32	289	33
rect	288	33	289	34
rect	288	34	289	35
rect	288	35	289	36
rect	288	36	289	37
rect	288	38	289	39
rect	288	39	289	40
rect	288	40	289	41
rect	288	41	289	42
rect	288	42	289	43
rect	288	43	289	44
rect	288	44	289	45
rect	288	45	289	46
rect	288	46	289	47
rect	288	48	289	49
rect	288	49	289	50
rect	288	50	289	51
rect	288	51	289	52
rect	288	52	289	53
rect	288	53	289	54
rect	288	54	289	55
rect	288	55	289	56
rect	288	56	289	57
rect	288	58	289	59
rect	288	59	289	60
rect	288	60	289	61
rect	288	61	289	62
rect	288	62	289	63
rect	288	63	289	64
rect	288	65	289	66
rect	288	66	289	67
rect	288	67	289	68
rect	288	68	289	69
rect	288	69	289	70
rect	288	70	289	71
rect	288	72	289	73
rect	288	73	289	74
rect	288	74	289	75
rect	288	75	289	76
rect	288	76	289	77
rect	288	77	289	78
rect	289	0	290	1
rect	289	1	290	2
rect	289	2	290	3
rect	289	3	290	4
rect	289	4	290	5
rect	289	5	290	6
rect	289	7	290	8
rect	289	8	290	9
rect	289	9	290	10
rect	289	10	290	11
rect	289	11	290	12
rect	289	12	290	13
rect	289	13	290	14
rect	289	14	290	15
rect	289	15	290	16
rect	289	17	290	18
rect	289	18	290	19
rect	289	19	290	20
rect	289	20	290	21
rect	289	21	290	22
rect	289	22	290	23
rect	289	24	290	25
rect	289	25	290	26
rect	289	26	290	27
rect	289	27	290	28
rect	289	28	290	29
rect	289	29	290	30
rect	289	31	290	32
rect	289	32	290	33
rect	289	33	290	34
rect	289	34	290	35
rect	289	35	290	36
rect	289	36	290	37
rect	289	38	290	39
rect	289	39	290	40
rect	289	40	290	41
rect	289	41	290	42
rect	289	42	290	43
rect	289	43	290	44
rect	289	44	290	45
rect	289	45	290	46
rect	289	46	290	47
rect	289	48	290	49
rect	289	49	290	50
rect	289	50	290	51
rect	289	51	290	52
rect	289	52	290	53
rect	289	53	290	54
rect	289	54	290	55
rect	289	55	290	56
rect	289	56	290	57
rect	289	58	290	59
rect	289	59	290	60
rect	289	60	290	61
rect	289	61	290	62
rect	289	62	290	63
rect	289	63	290	64
rect	289	65	290	66
rect	289	66	290	67
rect	289	67	290	68
rect	289	68	290	69
rect	289	69	290	70
rect	289	70	290	71
rect	289	72	290	73
rect	289	73	290	74
rect	289	74	290	75
rect	289	75	290	76
rect	289	76	290	77
rect	289	77	290	78
<< metal1 >>
rect	0	41	1	42
rect	0	42	1	43
rect	0	43	1	44
rect	0	44	1	45
rect	0	45	1	46
rect	2	38	3	39
rect	2	39	3	40
rect	2	41	3	42
rect	2	42	3	43
rect	2	64	3	65
rect	2	65	3	66
rect	2	66	3	67
rect	2	67	3	68
rect	2	68	3	69
rect	2	69	3	70
rect	2	70	3	71
rect	2	71	3	72
rect	2	72	3	73
rect	2	84	3	85
rect	2	85	3	86
rect	2	86	3	87
rect	2	91	3	92
rect	2	92	3	93
rect	4	5	5	6
rect	4	6	5	7
rect	4	7	5	8
rect	4	8	5	9
rect	4	9	5	10
rect	4	34	5	35
rect	4	35	5	36
rect	4	36	5	37
rect	4	38	5	39
rect	4	39	5	40
rect	4	41	5	42
rect	4	42	5	43
rect	4	44	5	45
rect	4	45	5	46
rect	4	47	5	48
rect	4	48	5	49
rect	4	49	5	50
rect	4	61	5	62
rect	4	62	5	63
rect	4	64	5	65
rect	4	65	5	66
rect	4	78	5	79
rect	4	79	5	80
rect	4	80	5	81
rect	4	81	5	82
rect	4	82	5	83
rect	4	84	5	85
rect	4	85	5	86
rect	4	86	5	87
rect	4	88	5	89
rect	4	89	5	90
rect	4	91	5	92
rect	4	92	5	93
rect	4	94	5	95
rect	4	95	5	96
rect	4	96	5	97
rect	4	97	5	98
rect	4	98	5	99
rect	4	99	5	100
rect	4	100	5	101
rect	4	101	5	102
rect	4	102	5	103
rect	6	2	7	3
rect	6	3	7	4
rect	6	5	7	6
rect	6	6	7	7
rect	6	18	7	19
rect	6	19	7	20
rect	6	24	7	25
rect	6	25	7	26
rect	6	26	7	27
rect	6	27	7	28
rect	6	28	7	29
rect	6	29	7	30
rect	6	30	7	31
rect	6	31	7	32
rect	6	32	7	33
rect	6	34	7	35
rect	6	35	7	36
rect	6	36	7	37
rect	6	38	7	39
rect	6	39	7	40
rect	6	41	7	42
rect	6	42	7	43
rect	6	44	7	45
rect	6	45	7	46
rect	6	47	7	48
rect	6	48	7	49
rect	6	49	7	50
rect	6	51	7	52
rect	6	52	7	53
rect	6	53	7	54
rect	6	54	7	55
rect	6	55	7	56
rect	6	56	7	57
rect	6	57	7	58
rect	6	58	7	59
rect	6	59	7	60
rect	6	61	7	62
rect	6	62	7	63
rect	6	64	7	65
rect	6	65	7	66
rect	6	67	7	68
rect	6	68	7	69
rect	6	69	7	70
rect	6	70	7	71
rect	6	71	7	72
rect	6	72	7	73
rect	6	74	7	75
rect	6	75	7	76
rect	6	76	7	77
rect	6	78	7	79
rect	6	79	7	80
rect	6	80	7	81
rect	6	81	7	82
rect	6	82	7	83
rect	6	84	7	85
rect	6	85	7	86
rect	6	86	7	87
rect	6	88	7	89
rect	6	89	7	90
rect	6	91	7	92
rect	6	92	7	93
rect	6	94	7	95
rect	6	95	7	96
rect	6	96	7	97
rect	15	51	16	52
rect	15	52	16	53
rect	15	55	16	56
rect	15	56	16	57
rect	15	57	16	58
rect	15	60	16	61
rect	15	61	16	62
rect	15	62	16	63
rect	15	64	16	65
rect	15	65	16	66
rect	15	67	16	68
rect	15	68	16	69
rect	15	69	16	70
rect	15	70	16	71
rect	17	44	18	45
rect	17	45	18	46
rect	17	47	18	48
rect	17	48	18	49
rect	17	49	18	50
rect	17	50	18	51
rect	17	51	18	52
rect	17	52	18	53
rect	17	78	18	79
rect	17	79	18	80
rect	17	82	18	83
rect	17	85	18	86
rect	17	86	18	87
rect	17	88	18	89
rect	17	89	18	90
rect	17	90	18	91
rect	17	91	18	92
rect	17	92	18	93
rect	17	94	18	95
rect	17	95	18	96
rect	17	96	18	97
rect	17	97	18	98
rect	17	98	18	99
rect	17	99	18	100
rect	17	101	18	102
rect	17	102	18	103
rect	17	104	18	105
rect	17	105	18	106
rect	17	106	18	107
rect	17	107	18	108
rect	17	108	18	109
rect	17	109	18	110
rect	17	110	18	111
rect	17	111	18	112
rect	17	112	18	113
rect	17	113	18	114
rect	17	114	18	115
rect	19	8	20	9
rect	19	9	20	10
rect	19	11	20	12
rect	19	12	20	13
rect	19	13	20	14
rect	19	15	20	16
rect	19	40	20	41
rect	19	41	20	42
rect	19	42	20	43
rect	19	43	20	44
rect	19	44	20	45
rect	19	45	20	46
rect	19	47	20	48
rect	19	48	20	49
rect	19	49	20	50
rect	19	50	20	51
rect	19	51	20	52
rect	19	52	20	53
rect	19	56	20	57
rect	19	57	20	58
rect	19	60	20	61
rect	19	61	20	62
rect	19	62	20	63
rect	19	64	20	65
rect	19	65	20	66
rect	19	67	20	68
rect	19	68	20	69
rect	19	69	20	70
rect	19	70	20	71
rect	19	76	20	77
rect	19	94	20	95
rect	19	95	20	96
rect	19	96	20	97
rect	19	97	20	98
rect	19	98	20	99
rect	19	99	20	100
rect	19	101	20	102
rect	19	102	20	103
rect	19	104	20	105
rect	19	105	20	106
rect	19	106	20	107
rect	19	107	20	108
rect	19	108	20	109
rect	19	109	20	110
rect	19	110	20	111
rect	19	111	20	112
rect	21	18	22	19
rect	21	21	22	22
rect	21	30	22	31
rect	21	31	22	32
rect	21	32	22	33
rect	21	38	22	39
rect	21	40	22	41
rect	21	41	22	42
rect	21	42	22	43
rect	21	43	22	44
rect	21	44	22	45
rect	21	45	22	46
rect	21	47	22	48
rect	21	48	22	49
rect	21	49	22	50
rect	21	50	22	51
rect	21	51	22	52
rect	21	94	22	95
rect	21	95	22	96
rect	21	96	22	97
rect	21	97	22	98
rect	21	98	22	99
rect	21	99	22	100
rect	21	101	22	102
rect	21	102	22	103
rect	21	104	22	105
rect	21	105	22	106
rect	21	106	22	107
rect	21	107	22	108
rect	21	108	22	109
rect	21	109	22	110
rect	21	110	22	111
rect	21	111	22	112
rect	21	113	22	114
rect	21	114	22	115
rect	21	116	22	117
rect	21	117	22	118
rect	21	118	22	119
rect	21	119	22	120
rect	21	120	22	121
rect	21	121	22	122
rect	21	122	22	123
rect	21	123	22	124
rect	21	124	22	125
rect	21	125	22	126
rect	21	126	22	127
rect	21	127	22	128
rect	21	128	22	129
rect	21	129	22	130
rect	21	130	22	131
rect	21	131	22	132
rect	21	132	22	133
rect	21	133	22	134
rect	21	134	22	135
rect	21	135	22	136
rect	21	136	22	137
rect	21	137	22	138
rect	21	138	22	139
rect	23	11	24	12
rect	23	12	24	13
rect	23	13	24	14
rect	23	21	24	22
rect	23	28	24	29
rect	23	30	24	31
rect	23	31	24	32
rect	23	32	24	33
rect	23	33	24	34
rect	23	36	24	37
rect	23	37	24	38
rect	23	38	24	39
rect	23	40	24	41
rect	23	41	24	42
rect	23	47	24	48
rect	23	48	24	49
rect	23	49	24	50
rect	23	50	24	51
rect	23	51	24	52
rect	23	56	24	57
rect	23	57	24	58
rect	23	62	24	63
rect	23	69	24	70
rect	23	70	24	71
rect	23	85	24	86
rect	23	86	24	87
rect	23	88	24	89
rect	23	89	24	90
rect	23	90	24	91
rect	23	91	24	92
rect	23	92	24	93
rect	23	94	24	95
rect	23	95	24	96
rect	23	104	24	105
rect	23	105	24	106
rect	23	106	24	107
rect	23	107	24	108
rect	23	108	24	109
rect	23	109	24	110
rect	23	110	24	111
rect	23	111	24	112
rect	23	113	24	114
rect	23	114	24	115
rect	23	116	24	117
rect	23	117	24	118
rect	23	118	24	119
rect	23	119	24	120
rect	23	120	24	121
rect	23	121	24	122
rect	23	122	24	123
rect	23	123	24	124
rect	23	124	24	125
rect	23	125	24	126
rect	23	126	24	127
rect	23	127	24	128
rect	23	128	24	129
rect	23	129	24	130
rect	23	130	24	131
rect	23	131	24	132
rect	23	132	24	133
rect	23	133	24	134
rect	23	134	24	135
rect	23	135	24	136
rect	23	136	24	137
rect	23	137	24	138
rect	23	138	24	139
rect	23	140	24	141
rect	23	141	24	142
rect	25	15	26	16
rect	25	18	26	19
rect	25	21	26	22
rect	25	24	26	25
rect	25	27	26	28
rect	25	28	26	29
rect	25	30	26	31
rect	25	31	26	32
rect	25	32	26	33
rect	25	33	26	34
rect	25	36	26	37
rect	25	37	26	38
rect	25	38	26	39
rect	25	40	26	41
rect	25	41	26	42
rect	25	43	26	44
rect	25	44	26	45
rect	25	45	26	46
rect	25	46	26	47
rect	25	47	26	48
rect	25	48	26	49
rect	25	49	26	50
rect	25	50	26	51
rect	25	51	26	52
rect	25	56	26	57
rect	25	57	26	58
rect	25	60	26	61
rect	25	62	26	63
rect	25	63	26	64
rect	25	64	26	65
rect	25	65	26	66
rect	25	67	26	68
rect	25	69	26	70
rect	25	70	26	71
rect	25	76	26	77
rect	25	78	26	79
rect	25	79	26	80
rect	25	82	26	83
rect	25	85	26	86
rect	25	86	26	87
rect	25	88	26	89
rect	25	89	26	90
rect	25	90	26	91
rect	25	91	26	92
rect	25	92	26	93
rect	25	94	26	95
rect	25	95	26	96
rect	25	97	26	98
rect	25	98	26	99
rect	25	100	26	101
rect	25	101	26	102
rect	27	2	28	3
rect	27	3	28	4
rect	27	12	28	13
rect	27	13	28	14
rect	27	15	28	16
rect	27	18	28	19
rect	27	27	28	28
rect	27	28	28	29
rect	27	30	28	31
rect	27	31	28	32
rect	27	32	28	33
rect	27	33	28	34
rect	27	36	28	37
rect	27	37	28	38
rect	27	38	28	39
rect	27	40	28	41
rect	27	41	28	42
rect	27	43	28	44
rect	27	44	28	45
rect	27	45	28	46
rect	27	46	28	47
rect	27	47	28	48
rect	27	48	28	49
rect	27	65	28	66
rect	27	82	28	83
rect	27	88	28	89
rect	27	89	28	90
rect	27	90	28	91
rect	27	91	28	92
rect	27	92	28	93
rect	27	94	28	95
rect	27	95	28	96
rect	27	97	28	98
rect	27	98	28	99
rect	27	100	28	101
rect	27	101	28	102
rect	27	103	28	104
rect	27	104	28	105
rect	27	105	28	106
rect	27	106	28	107
rect	27	107	28	108
rect	27	108	28	109
rect	27	109	28	110
rect	27	110	28	111
rect	27	111	28	112
rect	27	113	28	114
rect	27	114	28	115
rect	27	116	28	117
rect	27	117	28	118
rect	27	118	28	119
rect	27	119	28	120
rect	27	120	28	121
rect	27	121	28	122
rect	27	122	28	123
rect	27	123	28	124
rect	27	124	28	125
rect	27	125	28	126
rect	27	126	28	127
rect	27	127	28	128
rect	27	128	28	129
rect	27	129	28	130
rect	27	130	28	131
rect	27	131	28	132
rect	29	5	30	6
rect	29	6	30	7
rect	29	8	30	9
rect	29	9	30	10
rect	29	10	30	11
rect	29	12	30	13
rect	29	13	30	14
rect	29	15	30	16
rect	29	18	30	19
rect	29	21	30	22
rect	29	24	30	25
rect	29	27	30	28
rect	29	28	30	29
rect	29	30	30	31
rect	29	31	30	32
rect	29	37	30	38
rect	29	38	30	39
rect	29	40	30	41
rect	29	41	30	42
rect	29	43	30	44
rect	29	44	30	45
rect	29	45	30	46
rect	29	46	30	47
rect	29	47	30	48
rect	29	48	30	49
rect	29	50	30	51
rect	29	51	30	52
rect	29	56	30	57
rect	29	57	30	58
rect	29	60	30	61
rect	29	62	30	63
rect	29	63	30	64
rect	29	65	30	66
rect	29	66	30	67
rect	29	67	30	68
rect	29	69	30	70
rect	29	70	30	71
rect	29	76	30	77
rect	29	78	30	79
rect	29	79	30	80
rect	29	88	30	89
rect	29	89	30	90
rect	29	90	30	91
rect	29	91	30	92
rect	29	92	30	93
rect	29	94	30	95
rect	29	95	30	96
rect	29	97	30	98
rect	29	98	30	99
rect	29	100	30	101
rect	29	101	30	102
rect	29	103	30	104
rect	29	104	30	105
rect	29	105	30	106
rect	29	106	30	107
rect	29	107	30	108
rect	29	108	30	109
rect	29	109	30	110
rect	29	110	30	111
rect	29	111	30	112
rect	29	113	30	114
rect	29	114	30	115
rect	29	116	30	117
rect	29	117	30	118
rect	29	118	30	119
rect	29	119	30	120
rect	29	120	30	121
rect	29	121	30	122
rect	29	122	30	123
rect	29	123	30	124
rect	29	124	30	125
rect	29	125	30	126
rect	38	60	39	61
rect	38	62	39	63
rect	38	63	39	64
rect	38	65	39	66
rect	38	66	39	67
rect	38	67	39	68
rect	38	69	39	70
rect	40	60	41	61
rect	40	62	41	63
rect	40	63	41	64
rect	40	65	41	66
rect	40	66	41	67
rect	40	67	41	68
rect	42	56	43	57
rect	42	57	43	58
rect	42	60	43	61
rect	42	62	43	63
rect	42	63	43	64
rect	42	65	43	66
rect	42	66	43	67
rect	42	91	43	92
rect	42	92	43	93
rect	42	103	43	104
rect	42	104	43	105
rect	42	105	43	106
rect	42	106	43	107
rect	42	107	43	108
rect	44	11	45	12
rect	44	12	45	13
rect	44	13	45	14
rect	44	15	45	16
rect	44	18	45	19
rect	44	21	45	22
rect	44	24	45	25
rect	44	27	45	28
rect	44	28	45	29
rect	44	46	45	47
rect	44	47	45	48
rect	44	48	45	49
rect	44	49	45	50
rect	44	50	45	51
rect	44	51	45	52
rect	44	55	45	56
rect	44	56	45	57
rect	44	57	45	58
rect	44	60	45	61
rect	44	78	45	79
rect	44	79	45	80
rect	44	82	45	83
rect	44	85	45	86
rect	44	86	45	87
rect	44	87	45	88
rect	44	88	45	89
rect	44	100	45	101
rect	44	101	45	102
rect	44	102	45	103
rect	44	103	45	104
rect	44	104	45	105
rect	46	8	47	9
rect	46	9	47	10
rect	46	11	47	12
rect	46	12	47	13
rect	46	13	47	14
rect	46	15	47	16
rect	46	18	47	19
rect	46	21	47	22
rect	46	24	47	25
rect	46	27	47	28
rect	46	28	47	29
rect	46	55	47	56
rect	46	56	47	57
rect	46	57	47	58
rect	46	60	47	61
rect	46	65	47	66
rect	46	66	47	67
rect	46	68	47	69
rect	46	69	47	70
rect	46	71	47	72
rect	46	82	47	83
rect	46	85	47	86
rect	46	86	47	87
rect	46	87	47	88
rect	46	88	47	89
rect	46	90	47	91
rect	46	91	47	92
rect	46	97	47	98
rect	46	98	47	99
rect	46	99	47	100
rect	46	100	47	101
rect	46	101	47	102
rect	46	102	47	103
rect	46	103	47	104
rect	46	104	47	105
rect	46	106	47	107
rect	46	107	47	108
rect	46	109	47	110
rect	46	110	47	111
rect	46	111	47	112
rect	46	113	47	114
rect	46	114	47	115
rect	46	116	47	117
rect	46	117	47	118
rect	46	118	47	119
rect	46	119	47	120
rect	46	120	47	121
rect	46	121	47	122
rect	46	138	47	139
rect	46	139	47	140
rect	46	140	47	141
rect	46	141	47	142
rect	46	148	47	149
rect	46	149	47	150
rect	46	150	47	151
rect	46	151	47	152
rect	46	152	47	153
rect	46	153	47	154
rect	46	154	47	155
rect	46	155	47	156
rect	46	156	47	157
rect	48	8	49	9
rect	48	9	49	10
rect	48	11	49	12
rect	48	12	49	13
rect	48	13	49	14
rect	48	15	49	16
rect	48	18	49	19
rect	48	21	49	22
rect	48	24	49	25
rect	48	40	49	41
rect	48	41	49	42
rect	48	43	49	44
rect	48	44	49	45
rect	48	46	49	47
rect	48	47	49	48
rect	48	48	49	49
rect	48	49	49	50
rect	48	50	49	51
rect	48	51	49	52
rect	48	52	49	53
rect	48	55	49	56
rect	48	56	49	57
rect	48	57	49	58
rect	48	60	49	61
rect	48	62	49	63
rect	48	63	49	64
rect	48	64	49	65
rect	48	65	49	66
rect	48	66	49	67
rect	48	68	49	69
rect	48	69	49	70
rect	48	71	49	72
rect	48	77	49	78
rect	48	78	49	79
rect	48	79	49	80
rect	48	82	49	83
rect	48	85	49	86
rect	48	86	49	87
rect	48	87	49	88
rect	48	88	49	89
rect	48	90	49	91
rect	48	91	49	92
rect	48	93	49	94
rect	48	94	49	95
rect	48	95	49	96
rect	48	96	49	97
rect	48	97	49	98
rect	48	98	49	99
rect	48	99	49	100
rect	48	100	49	101
rect	48	101	49	102
rect	48	102	49	103
rect	48	103	49	104
rect	48	104	49	105
rect	48	106	49	107
rect	48	107	49	108
rect	48	109	49	110
rect	48	110	49	111
rect	48	111	49	112
rect	48	113	49	114
rect	48	114	49	115
rect	48	116	49	117
rect	48	117	49	118
rect	48	118	49	119
rect	48	119	49	120
rect	48	120	49	121
rect	48	121	49	122
rect	48	122	49	123
rect	48	123	49	124
rect	48	124	49	125
rect	48	125	49	126
rect	48	126	49	127
rect	48	127	49	128
rect	48	128	49	129
rect	48	130	49	131
rect	48	131	49	132
rect	48	133	49	134
rect	48	134	49	135
rect	48	135	49	136
rect	48	136	49	137
rect	48	138	49	139
rect	48	139	49	140
rect	48	140	49	141
rect	48	141	49	142
rect	48	142	49	143
rect	48	143	49	144
rect	48	144	49	145
rect	48	145	49	146
rect	48	146	49	147
rect	48	148	49	149
rect	48	149	49	150
rect	48	150	49	151
rect	48	151	49	152
rect	48	152	49	153
rect	48	153	49	154
rect	48	154	49	155
rect	48	155	49	156
rect	48	156	49	157
rect	48	158	49	159
rect	48	159	49	160
rect	48	160	49	161
rect	48	161	49	162
rect	48	162	49	163
rect	48	163	49	164
rect	48	164	49	165
rect	48	165	49	166
rect	50	24	51	25
rect	50	33	51	34
rect	50	36	51	37
rect	50	37	51	38
rect	50	38	51	39
rect	50	43	51	44
rect	50	44	51	45
rect	50	46	51	47
rect	50	47	51	48
rect	50	48	51	49
rect	50	49	51	50
rect	50	50	51	51
rect	50	51	51	52
rect	50	52	51	53
rect	50	55	51	56
rect	50	56	51	57
rect	50	57	51	58
rect	50	60	51	61
rect	50	62	51	63
rect	50	63	51	64
rect	50	77	51	78
rect	50	78	51	79
rect	50	79	51	80
rect	50	82	51	83
rect	50	85	51	86
rect	50	86	51	87
rect	50	87	51	88
rect	50	88	51	89
rect	50	90	51	91
rect	50	91	51	92
rect	50	93	51	94
rect	50	94	51	95
rect	50	95	51	96
rect	50	96	51	97
rect	50	97	51	98
rect	50	98	51	99
rect	50	99	51	100
rect	50	100	51	101
rect	50	101	51	102
rect	50	113	51	114
rect	50	114	51	115
rect	50	116	51	117
rect	50	117	51	118
rect	50	118	51	119
rect	50	119	51	120
rect	50	120	51	121
rect	50	121	51	122
rect	50	122	51	123
rect	50	123	51	124
rect	50	133	51	134
rect	50	134	51	135
rect	50	135	51	136
rect	50	136	51	137
rect	50	138	51	139
rect	50	139	51	140
rect	50	140	51	141
rect	50	141	51	142
rect	50	142	51	143
rect	50	143	51	144
rect	50	144	51	145
rect	50	145	51	146
rect	50	146	51	147
rect	50	148	51	149
rect	50	149	51	150
rect	50	150	51	151
rect	50	151	51	152
rect	50	152	51	153
rect	50	153	51	154
rect	50	154	51	155
rect	50	155	51	156
rect	50	156	51	157
rect	50	158	51	159
rect	50	159	51	160
rect	52	15	53	16
rect	52	21	53	22
rect	52	36	53	37
rect	52	37	53	38
rect	52	38	53	39
rect	52	40	53	41
rect	52	41	53	42
rect	52	50	53	51
rect	52	51	53	52
rect	52	52	53	53
rect	52	77	53	78
rect	52	78	53	79
rect	52	79	53	80
rect	52	82	53	83
rect	52	87	53	88
rect	52	88	53	89
rect	52	90	53	91
rect	52	91	53	92
rect	52	93	53	94
rect	52	94	53	95
rect	52	95	53	96
rect	52	100	53	101
rect	52	101	53	102
rect	52	103	53	104
rect	52	104	53	105
rect	52	106	53	107
rect	52	107	53	108
rect	52	109	53	110
rect	52	110	53	111
rect	52	111	53	112
rect	52	112	53	113
rect	52	113	53	114
rect	52	114	53	115
rect	52	116	53	117
rect	52	117	53	118
rect	52	118	53	119
rect	52	119	53	120
rect	52	120	53	121
rect	52	121	53	122
rect	52	122	53	123
rect	52	123	53	124
rect	52	125	53	126
rect	52	126	53	127
rect	52	127	53	128
rect	52	128	53	129
rect	52	130	53	131
rect	52	131	53	132
rect	52	132	53	133
rect	52	133	53	134
rect	52	134	53	135
rect	52	135	53	136
rect	52	136	53	137
rect	52	138	53	139
rect	52	139	53	140
rect	52	140	53	141
rect	52	141	53	142
rect	52	142	53	143
rect	52	143	53	144
rect	52	144	53	145
rect	52	145	53	146
rect	52	146	53	147
rect	52	148	53	149
rect	52	149	53	150
rect	52	150	53	151
rect	52	151	53	152
rect	52	152	53	153
rect	52	153	53	154
rect	52	154	53	155
rect	52	155	53	156
rect	52	156	53	157
rect	52	158	53	159
rect	52	159	53	160
rect	52	161	53	162
rect	52	162	53	163
rect	54	5	55	6
rect	54	6	55	7
rect	54	8	55	9
rect	54	9	55	10
rect	54	11	55	12
rect	54	12	55	13
rect	54	21	55	22
rect	54	24	55	25
rect	54	27	55	28
rect	54	28	55	29
rect	54	30	55	31
rect	54	31	55	32
rect	54	32	55	33
rect	54	36	55	37
rect	54	37	55	38
rect	54	38	55	39
rect	54	40	55	41
rect	54	41	55	42
rect	54	43	55	44
rect	54	44	55	45
rect	54	46	55	47
rect	54	47	55	48
rect	54	48	55	49
rect	54	50	55	51
rect	54	51	55	52
rect	54	52	55	53
rect	54	56	55	57
rect	54	57	55	58
rect	54	60	55	61
rect	54	62	55	63
rect	54	63	55	64
rect	54	65	55	66
rect	54	66	55	67
rect	54	68	55	69
rect	54	69	55	70
rect	54	71	55	72
rect	54	77	55	78
rect	54	78	55	79
rect	54	79	55	80
rect	54	82	55	83
rect	54	85	55	86
rect	54	87	55	88
rect	54	88	55	89
rect	54	90	55	91
rect	54	91	55	92
rect	54	93	55	94
rect	54	94	55	95
rect	54	95	55	96
rect	54	97	55	98
rect	54	98	55	99
rect	54	100	55	101
rect	54	101	55	102
rect	54	103	55	104
rect	54	104	55	105
rect	54	106	55	107
rect	54	107	55	108
rect	54	109	55	110
rect	54	110	55	111
rect	54	116	55	117
rect	54	117	55	118
rect	54	118	55	119
rect	54	119	55	120
rect	54	120	55	121
rect	54	130	55	131
rect	54	131	55	132
rect	54	132	55	133
rect	54	133	55	134
rect	54	142	55	143
rect	54	143	55	144
rect	54	144	55	145
rect	54	145	55	146
rect	54	146	55	147
rect	54	148	55	149
rect	54	149	55	150
rect	63	167	64	168
rect	63	168	64	169
rect	63	169	64	170
rect	63	170	64	171
rect	63	171	64	172
rect	63	172	64	173
rect	63	173	64	174
rect	63	174	64	175
rect	63	175	64	176
rect	63	176	64	177
rect	63	177	64	178
rect	65	116	66	117
rect	65	117	66	118
rect	65	118	66	119
rect	65	119	66	120
rect	65	120	66	121
rect	65	122	66	123
rect	65	123	66	124
rect	65	125	66	126
rect	65	126	66	127
rect	65	127	66	128
rect	65	129	66	130
rect	65	130	66	131
rect	65	131	66	132
rect	65	132	66	133
rect	65	133	66	134
rect	65	135	66	136
rect	65	136	66	137
rect	65	138	66	139
rect	65	139	66	140
rect	65	140	66	141
rect	65	141	66	142
rect	65	142	66	143
rect	65	143	66	144
rect	65	144	66	145
rect	65	145	66	146
rect	65	146	66	147
rect	65	148	66	149
rect	65	149	66	150
rect	65	151	66	152
rect	65	152	66	153
rect	65	153	66	154
rect	65	155	66	156
rect	65	156	66	157
rect	65	157	66	158
rect	65	158	66	159
rect	65	159	66	160
rect	65	161	66	162
rect	65	162	66	163
rect	65	164	66	165
rect	65	165	66	166
rect	67	112	68	113
rect	67	113	68	114
rect	67	114	68	115
rect	69	109	70	110
rect	69	110	70	111
rect	69	111	70	112
rect	69	155	70	156
rect	69	156	70	157
rect	69	157	70	158
rect	69	158	70	159
rect	69	159	70	160
rect	69	161	70	162
rect	69	162	70	163
rect	69	164	70	165
rect	69	165	70	166
rect	69	167	70	168
rect	69	168	70	169
rect	69	169	70	170
rect	69	170	70	171
rect	69	171	70	172
rect	69	172	70	173
rect	69	173	70	174
rect	69	174	70	175
rect	69	175	70	176
rect	69	176	70	177
rect	69	177	70	178
rect	69	179	70	180
rect	69	180	70	181
rect	69	181	70	182
rect	69	182	70	183
rect	69	183	70	184
rect	69	184	70	185
rect	69	185	70	186
rect	69	186	70	187
rect	69	187	70	188
rect	69	188	70	189
rect	69	189	70	190
rect	69	190	70	191
rect	69	191	70	192
rect	69	192	70	193
rect	69	193	70	194
rect	69	194	70	195
rect	69	195	70	196
rect	69	196	70	197
rect	69	197	70	198
rect	69	198	70	199
rect	69	199	70	200
rect	69	200	70	201
rect	69	201	70	202
rect	69	202	70	203
rect	69	203	70	204
rect	69	204	70	205
rect	69	205	70	206
rect	69	206	70	207
rect	69	207	70	208
rect	71	62	72	63
rect	71	63	72	64
rect	71	65	72	66
rect	71	66	72	67
rect	71	68	72	69
rect	71	69	72	70
rect	71	71	72	72
rect	71	77	72	78
rect	71	78	72	79
rect	71	79	72	80
rect	71	82	72	83
rect	71	106	72	107
rect	71	107	72	108
rect	71	108	72	109
rect	71	135	72	136
rect	71	136	72	137
rect	71	138	72	139
rect	71	139	72	140
rect	71	140	72	141
rect	71	141	72	142
rect	71	142	72	143
rect	71	143	72	144
rect	71	144	72	145
rect	71	145	72	146
rect	71	146	72	147
rect	71	148	72	149
rect	71	149	72	150
rect	71	151	72	152
rect	71	152	72	153
rect	73	77	74	78
rect	73	78	74	79
rect	73	79	74	80
rect	73	82	74	83
rect	73	103	74	104
rect	73	104	74	105
rect	73	105	74	106
rect	73	106	74	107
rect	73	107	74	108
rect	73	108	74	109
rect	73	110	74	111
rect	73	111	74	112
rect	73	113	74	114
rect	73	114	74	115
rect	73	116	74	117
rect	73	117	74	118
rect	73	118	74	119
rect	73	119	74	120
rect	73	120	74	121
rect	73	122	74	123
rect	73	123	74	124
rect	73	125	74	126
rect	73	126	74	127
rect	73	127	74	128
rect	73	129	74	130
rect	73	130	74	131
rect	73	131	74	132
rect	73	132	74	133
rect	73	133	74	134
rect	75	76	76	77
rect	75	77	76	78
rect	75	78	76	79
rect	75	79	76	80
rect	75	93	76	94
rect	75	94	76	95
rect	75	95	76	96
rect	75	96	76	97
rect	75	97	76	98
rect	75	98	76	99
rect	75	99	76	100
rect	75	100	76	101
rect	75	101	76	102
rect	75	102	76	103
rect	75	103	76	104
rect	75	104	76	105
rect	75	105	76	106
rect	75	125	76	126
rect	75	126	76	127
rect	75	127	76	128
rect	75	129	76	130
rect	75	130	76	131
rect	75	131	76	132
rect	75	132	76	133
rect	75	133	76	134
rect	75	135	76	136
rect	75	136	76	137
rect	75	138	76	139
rect	75	139	76	140
rect	75	148	76	149
rect	75	149	76	150
rect	75	151	76	152
rect	75	152	76	153
rect	75	154	76	155
rect	75	155	76	156
rect	77	71	78	72
rect	77	76	78	77
rect	77	90	78	91
rect	77	91	78	92
rect	77	92	78	93
rect	77	93	78	94
rect	77	94	78	95
rect	77	95	78	96
rect	77	96	78	97
rect	77	97	78	98
rect	77	98	78	99
rect	77	99	78	100
rect	77	100	78	101
rect	77	101	78	102
rect	77	102	78	103
rect	77	126	78	127
rect	77	127	78	128
rect	77	129	78	130
rect	77	130	78	131
rect	77	131	78	132
rect	77	132	78	133
rect	77	133	78	134
rect	77	135	78	136
rect	77	136	78	137
rect	77	138	78	139
rect	77	139	78	140
rect	77	141	78	142
rect	77	142	78	143
rect	77	143	78	144
rect	77	144	78	145
rect	77	145	78	146
rect	77	146	78	147
rect	79	68	80	69
rect	79	69	80	70
rect	79	70	80	71
rect	79	71	80	72
rect	79	87	80	88
rect	79	88	80	89
rect	79	89	80	90
rect	79	90	80	91
rect	79	91	80	92
rect	79	92	80	93
rect	79	98	80	99
rect	79	99	80	100
rect	79	100	80	101
rect	79	101	80	102
rect	79	102	80	103
rect	79	104	80	105
rect	79	105	80	106
rect	79	107	80	108
rect	79	108	80	109
rect	79	110	80	111
rect	79	111	80	112
rect	79	113	80	114
rect	79	114	80	115
rect	79	116	80	117
rect	79	117	80	118
rect	79	118	80	119
rect	79	119	80	120
rect	79	120	80	121
rect	79	122	80	123
rect	79	123	80	124
rect	79	124	80	125
rect	79	126	80	127
rect	79	127	80	128
rect	79	129	80	130
rect	79	130	80	131
rect	79	131	80	132
rect	79	132	80	133
rect	79	133	80	134
rect	79	135	80	136
rect	79	136	80	137
rect	79	138	80	139
rect	79	139	80	140
rect	79	141	80	142
rect	79	142	80	143
rect	79	143	80	144
rect	79	144	80	145
rect	79	145	80	146
rect	79	146	80	147
rect	79	148	80	149
rect	79	149	80	150
rect	79	151	80	152
rect	79	152	80	153
rect	79	154	80	155
rect	79	155	80	156
rect	79	157	80	158
rect	79	158	80	159
rect	79	159	80	160
rect	79	161	80	162
rect	79	162	80	163
rect	79	164	80	165
rect	79	165	80	166
rect	79	167	80	168
rect	79	168	80	169
rect	81	18	82	19
rect	81	21	82	22
rect	81	24	82	25
rect	81	27	82	28
rect	81	28	82	29
rect	81	43	82	44
rect	81	44	82	45
rect	81	46	82	47
rect	81	47	82	48
rect	81	48	82	49
rect	81	50	82	51
rect	81	51	82	52
rect	81	65	82	66
rect	81	66	82	67
rect	81	67	82	68
rect	81	76	82	77
rect	81	78	82	79
rect	81	79	82	80
rect	81	82	82	83
rect	81	85	82	86
rect	81	86	82	87
rect	81	87	82	88
rect	81	88	82	89
rect	81	89	82	90
rect	81	90	82	91
rect	81	91	82	92
rect	81	92	82	93
rect	81	94	82	95
rect	81	95	82	96
rect	81	96	82	97
rect	81	98	82	99
rect	81	99	82	100
rect	81	100	82	101
rect	81	101	82	102
rect	81	102	82	103
rect	81	104	82	105
rect	81	105	82	106
rect	81	107	82	108
rect	81	108	82	109
rect	81	110	82	111
rect	81	111	82	112
rect	81	113	82	114
rect	81	114	82	115
rect	81	116	82	117
rect	81	117	82	118
rect	81	118	82	119
rect	81	119	82	120
rect	81	120	82	121
rect	81	122	82	123
rect	81	123	82	124
rect	81	124	82	125
rect	81	126	82	127
rect	81	127	82	128
rect	83	27	84	28
rect	83	28	84	29
rect	83	40	84	41
rect	83	41	84	42
rect	83	42	84	43
rect	83	43	84	44
rect	83	44	84	45
rect	83	46	84	47
rect	83	47	84	48
rect	83	48	84	49
rect	83	60	84	61
rect	83	61	84	62
rect	83	62	84	63
rect	83	63	84	64
rect	83	64	84	65
rect	83	65	84	66
rect	83	66	84	67
rect	83	67	84	68
rect	83	69	84	70
rect	83	70	84	71
rect	83	76	84	77
rect	83	78	84	79
rect	83	79	84	80
rect	83	82	84	83
rect	83	85	84	86
rect	83	86	84	87
rect	83	87	84	88
rect	83	88	84	89
rect	83	89	84	90
rect	83	90	84	91
rect	83	91	84	92
rect	83	92	84	93
rect	83	94	84	95
rect	83	95	84	96
rect	83	96	84	97
rect	83	98	84	99
rect	83	99	84	100
rect	83	122	84	123
rect	83	123	84	124
rect	83	124	84	125
rect	83	126	84	127
rect	83	127	84	128
rect	83	164	84	165
rect	83	165	84	166
rect	83	167	84	168
rect	83	168	84	169
rect	83	170	84	171
rect	83	171	84	172
rect	85	2	86	3
rect	85	3	86	4
rect	85	4	86	5
rect	85	5	86	6
rect	85	6	86	7
rect	85	8	86	9
rect	85	9	86	10
rect	85	14	86	15
rect	85	15	86	16
rect	85	18	86	19
rect	85	21	86	22
rect	85	24	86	25
rect	85	37	86	38
rect	85	38	86	39
rect	85	43	86	44
rect	85	44	86	45
rect	85	56	86	57
rect	85	57	86	58
rect	85	60	86	61
rect	85	61	86	62
rect	85	66	86	67
rect	85	67	86	68
rect	85	69	86	70
rect	85	70	86	71
rect	85	76	86	77
rect	85	78	86	79
rect	85	79	86	80
rect	85	82	86	83
rect	85	85	86	86
rect	85	86	86	87
rect	85	87	86	88
rect	85	88	86	89
rect	85	89	86	90
rect	85	90	86	91
rect	85	91	86	92
rect	85	92	86	93
rect	85	94	86	95
rect	85	95	86	96
rect	85	96	86	97
rect	85	98	86	99
rect	85	99	86	100
rect	85	101	86	102
rect	85	102	86	103
rect	85	104	86	105
rect	85	105	86	106
rect	85	107	86	108
rect	85	108	86	109
rect	85	110	86	111
rect	85	111	86	112
rect	85	113	86	114
rect	85	114	86	115
rect	85	116	86	117
rect	85	117	86	118
rect	85	118	86	119
rect	85	119	86	120
rect	85	120	86	121
rect	85	121	86	122
rect	85	122	86	123
rect	85	123	86	124
rect	85	124	86	125
rect	85	126	86	127
rect	85	127	86	128
rect	85	129	86	130
rect	85	130	86	131
rect	85	131	86	132
rect	85	132	86	133
rect	85	133	86	134
rect	85	135	86	136
rect	85	136	86	137
rect	85	138	86	139
rect	85	139	86	140
rect	85	141	86	142
rect	85	142	86	143
rect	85	143	86	144
rect	85	144	86	145
rect	85	145	86	146
rect	85	146	86	147
rect	85	148	86	149
rect	85	149	86	150
rect	85	151	86	152
rect	85	152	86	153
rect	85	154	86	155
rect	85	155	86	156
rect	85	157	86	158
rect	85	158	86	159
rect	85	159	86	160
rect	85	161	86	162
rect	85	162	86	163
rect	87	5	88	6
rect	87	6	88	7
rect	87	12	88	13
rect	87	13	88	14
rect	87	37	88	38
rect	87	38	88	39
rect	87	40	88	41
rect	87	41	88	42
rect	87	43	88	44
rect	87	44	88	45
rect	87	45	88	46
rect	87	46	88	47
rect	87	47	88	48
rect	87	48	88	49
rect	87	49	88	50
rect	87	50	88	51
rect	87	51	88	52
rect	87	55	88	56
rect	87	56	88	57
rect	87	57	88	58
rect	87	60	88	61
rect	87	61	88	62
rect	87	63	88	64
rect	87	64	88	65
rect	87	66	88	67
rect	87	67	88	68
rect	87	69	88	70
rect	87	70	88	71
rect	87	76	88	77
rect	87	78	88	79
rect	87	79	88	80
rect	87	82	88	83
rect	87	85	88	86
rect	87	86	88	87
rect	87	87	88	88
rect	87	88	88	89
rect	87	89	88	90
rect	87	90	88	91
rect	87	91	88	92
rect	87	92	88	93
rect	87	94	88	95
rect	87	95	88	96
rect	87	96	88	97
rect	87	98	88	99
rect	87	99	88	100
rect	87	101	88	102
rect	87	102	88	103
rect	87	104	88	105
rect	87	105	88	106
rect	87	107	88	108
rect	87	108	88	109
rect	87	110	88	111
rect	87	111	88	112
rect	87	113	88	114
rect	87	114	88	115
rect	87	116	88	117
rect	87	117	88	118
rect	87	118	88	119
rect	87	119	88	120
rect	87	120	88	121
rect	87	121	88	122
rect	87	122	88	123
rect	87	123	88	124
rect	87	124	88	125
rect	87	126	88	127
rect	87	127	88	128
rect	87	129	88	130
rect	87	130	88	131
rect	87	161	88	162
rect	87	162	88	163
rect	87	164	88	165
rect	87	165	88	166
rect	87	167	88	168
rect	87	168	88	169
rect	87	170	88	171
rect	87	171	88	172
rect	87	173	88	174
rect	87	174	88	175
rect	102	40	103	41
rect	102	41	103	42
rect	102	43	103	44
rect	102	44	103	45
rect	102	45	103	46
rect	102	46	103	47
rect	102	47	103	48
rect	102	48	103	49
rect	102	49	103	50
rect	102	50	103	51
rect	102	51	103	52
rect	102	55	103	56
rect	102	56	103	57
rect	102	57	103	58
rect	102	60	103	61
rect	102	61	103	62
rect	102	63	103	64
rect	102	64	103	65
rect	102	66	103	67
rect	102	67	103	68
rect	102	69	103	70
rect	102	70	103	71
rect	102	74	103	75
rect	102	76	103	77
rect	102	78	103	79
rect	102	79	103	80
rect	102	80	103	81
rect	102	82	103	83
rect	102	85	103	86
rect	102	86	103	87
rect	102	88	103	89
rect	102	89	103	90
rect	102	91	103	92
rect	102	92	103	93
rect	102	94	103	95
rect	102	95	103	96
rect	102	96	103	97
rect	102	98	103	99
rect	102	99	103	100
rect	102	123	103	124
rect	102	124	103	125
rect	102	126	103	127
rect	102	127	103	128
rect	104	39	105	40
rect	104	40	105	41
rect	104	41	105	42
rect	104	43	105	44
rect	104	44	105	45
rect	104	45	105	46
rect	104	46	105	47
rect	104	47	105	48
rect	104	48	105	49
rect	104	49	105	50
rect	104	50	105	51
rect	104	51	105	52
rect	104	55	105	56
rect	104	56	105	57
rect	104	57	105	58
rect	104	60	105	61
rect	104	61	105	62
rect	104	63	105	64
rect	104	64	105	65
rect	104	66	105	67
rect	104	67	105	68
rect	104	69	105	70
rect	104	70	105	71
rect	104	74	105	75
rect	104	76	105	77
rect	104	78	105	79
rect	104	79	105	80
rect	104	80	105	81
rect	104	82	105	83
rect	104	85	105	86
rect	104	86	105	87
rect	104	91	105	92
rect	104	92	105	93
rect	104	94	105	95
rect	104	95	105	96
rect	104	96	105	97
rect	104	98	105	99
rect	104	99	105	100
rect	104	110	105	111
rect	104	111	105	112
rect	104	113	105	114
rect	104	114	105	115
rect	104	116	105	117
rect	104	117	105	118
rect	104	118	105	119
rect	104	120	105	121
rect	104	121	105	122
rect	104	122	105	123
rect	104	123	105	124
rect	104	124	105	125
rect	104	126	105	127
rect	104	127	105	128
rect	104	128	105	129
rect	106	48	107	49
rect	106	49	107	50
rect	106	50	107	51
rect	106	51	107	52
rect	106	55	107	56
rect	106	56	107	57
rect	106	57	107	58
rect	106	60	107	61
rect	106	61	107	62
rect	106	63	107	64
rect	106	64	107	65
rect	106	69	107	70
rect	106	70	107	71
rect	106	74	107	75
rect	106	76	107	77
rect	106	78	107	79
rect	106	79	107	80
rect	106	80	107	81
rect	106	82	107	83
rect	106	85	107	86
rect	106	86	107	87
rect	106	87	107	88
rect	106	111	107	112
rect	106	113	107	114
rect	106	114	107	115
rect	106	116	107	117
rect	106	117	107	118
rect	106	118	107	119
rect	106	120	107	121
rect	106	121	107	122
rect	106	122	107	123
rect	106	123	107	124
rect	106	124	107	125
rect	108	67	109	68
rect	108	68	109	69
rect	108	69	109	70
rect	108	70	109	71
rect	108	74	109	75
rect	108	76	109	77
rect	108	78	109	79
rect	108	79	109	80
rect	108	80	109	81
rect	108	82	109	83
rect	108	85	109	86
rect	108	86	109	87
rect	108	87	109	88
rect	108	89	109	90
rect	108	90	109	91
rect	108	91	109	92
rect	108	92	109	93
rect	108	127	109	128
rect	108	128	109	129
rect	108	130	109	131
rect	108	148	109	149
rect	108	149	109	150
rect	110	63	111	64
rect	110	64	111	65
rect	110	65	111	66
rect	110	67	111	68
rect	110	68	111	69
rect	110	69	111	70
rect	110	70	111	71
rect	110	74	111	75
rect	110	76	111	77
rect	110	78	111	79
rect	110	79	111	80
rect	110	80	111	81
rect	110	82	111	83
rect	110	85	111	86
rect	110	86	111	87
rect	110	87	111	88
rect	110	89	111	90
rect	110	90	111	91
rect	110	91	111	92
rect	110	92	111	93
rect	110	93	111	94
rect	110	94	111	95
rect	110	95	111	96
rect	110	96	111	97
rect	110	98	111	99
rect	110	99	111	100
rect	110	101	111	102
rect	110	102	111	103
rect	110	104	111	105
rect	110	105	111	106
rect	110	107	111	108
rect	110	108	111	109
rect	110	109	111	110
rect	110	111	111	112
rect	110	113	111	114
rect	110	114	111	115
rect	110	116	111	117
rect	110	117	111	118
rect	110	118	111	119
rect	110	120	111	121
rect	110	121	111	122
rect	110	122	111	123
rect	110	123	111	124
rect	110	124	111	125
rect	110	125	111	126
rect	110	127	111	128
rect	110	128	111	129
rect	110	130	111	131
rect	110	131	111	132
rect	110	132	111	133
rect	110	133	111	134
rect	110	135	111	136
rect	110	136	111	137
rect	110	138	111	139
rect	110	139	111	140
rect	110	141	111	142
rect	110	142	111	143
rect	110	143	111	144
rect	110	145	111	146
rect	110	146	111	147
rect	110	147	111	148
rect	110	148	111	149
rect	110	149	111	150
rect	110	150	111	151
rect	110	151	111	152
rect	110	152	111	153
rect	110	154	111	155
rect	110	155	111	156
rect	110	157	111	158
rect	110	158	111	159
rect	110	159	111	160
rect	110	161	111	162
rect	110	162	111	163
rect	110	163	111	164
rect	110	164	111	165
rect	110	165	111	166
rect	110	167	111	168
rect	110	168	111	169
rect	110	170	111	171
rect	110	171	111	172
rect	110	173	111	174
rect	110	174	111	175
rect	110	176	111	177
rect	110	177	111	178
rect	110	179	111	180
rect	110	180	111	181
rect	110	181	111	182
rect	110	182	111	183
rect	110	183	111	184
rect	110	184	111	185
rect	110	185	111	186
rect	110	186	111	187
rect	110	187	111	188
rect	110	188	111	189
rect	110	189	111	190
rect	110	190	111	191
rect	110	191	111	192
rect	110	192	111	193
rect	110	193	111	194
rect	110	194	111	195
rect	110	195	111	196
rect	112	27	113	28
rect	112	28	113	29
rect	112	30	113	31
rect	112	64	113	65
rect	112	65	113	66
rect	112	67	113	68
rect	112	68	113	69
rect	112	69	113	70
rect	112	70	113	71
rect	112	78	113	79
rect	112	79	113	80
rect	112	80	113	81
rect	112	82	113	83
rect	112	85	113	86
rect	112	86	113	87
rect	112	87	113	88
rect	112	89	113	90
rect	112	90	113	91
rect	112	91	113	92
rect	112	92	113	93
rect	112	93	113	94
rect	112	94	113	95
rect	112	95	113	96
rect	112	96	113	97
rect	112	104	113	105
rect	112	105	113	106
rect	112	107	113	108
rect	112	108	113	109
rect	112	109	113	110
rect	112	111	113	112
rect	112	113	113	114
rect	112	114	113	115
rect	112	116	113	117
rect	112	117	113	118
rect	112	118	113	119
rect	112	133	113	134
rect	112	135	113	136
rect	112	136	113	137
rect	112	138	113	139
rect	112	139	113	140
rect	112	141	113	142
rect	112	142	113	143
rect	112	143	113	144
rect	112	145	113	146
rect	112	146	113	147
rect	112	147	113	148
rect	112	148	113	149
rect	112	149	113	150
rect	112	150	113	151
rect	112	151	113	152
rect	112	152	113	153
rect	112	154	113	155
rect	112	155	113	156
rect	114	21	115	22
rect	114	24	115	25
rect	114	36	115	37
rect	114	37	115	38
rect	114	39	115	40
rect	114	40	115	41
rect	114	41	115	42
rect	114	61	115	62
rect	114	62	115	63
rect	114	64	115	65
rect	114	65	115	66
rect	114	67	115	68
rect	114	68	115	69
rect	114	69	115	70
rect	114	70	115	71
rect	114	71	115	72
rect	114	74	115	75
rect	114	76	115	77
rect	114	77	115	78
rect	114	78	115	79
rect	114	79	115	80
rect	114	80	115	81
rect	114	82	115	83
rect	114	85	115	86
rect	114	86	115	87
rect	114	87	115	88
rect	114	89	115	90
rect	114	90	115	91
rect	114	98	115	99
rect	114	99	115	100
rect	114	101	115	102
rect	114	102	115	103
rect	114	103	115	104
rect	114	104	115	105
rect	114	105	115	106
rect	114	135	115	136
rect	114	136	115	137
rect	114	138	115	139
rect	114	139	115	140
rect	114	141	115	142
rect	114	142	115	143
rect	114	143	115	144
rect	114	149	115	150
rect	114	150	115	151
rect	114	151	115	152
rect	114	152	115	153
rect	114	158	115	159
rect	114	159	115	160
rect	114	161	115	162
rect	114	162	115	163
rect	114	163	115	164
rect	114	164	115	165
rect	114	165	115	166
rect	114	167	115	168
rect	114	168	115	169
rect	114	170	115	171
rect	114	171	115	172
rect	114	173	115	174
rect	114	174	115	175
rect	116	18	117	19
rect	116	30	117	31
rect	116	32	117	33
rect	116	33	117	34
rect	116	55	117	56
rect	116	56	117	57
rect	116	61	117	62
rect	116	62	117	63
rect	116	64	117	65
rect	116	65	117	66
rect	116	67	117	68
rect	116	68	117	69
rect	116	69	117	70
rect	116	70	117	71
rect	116	71	117	72
rect	116	95	117	96
rect	116	96	117	97
rect	116	98	117	99
rect	116	99	117	100
rect	116	101	117	102
rect	116	102	117	103
rect	116	103	117	104
rect	116	136	117	137
rect	116	143	117	144
rect	116	144	117	145
rect	116	145	117	146
rect	116	146	117	147
rect	116	147	117	148
rect	116	149	117	150
rect	116	150	117	151
rect	116	173	117	174
rect	116	174	117	175
rect	116	175	117	176
rect	118	15	119	16
rect	118	18	119	19
rect	118	21	119	22
rect	118	24	119	25
rect	118	27	119	28
rect	118	55	119	56
rect	118	56	119	57
rect	118	61	119	62
rect	118	62	119	63
rect	118	64	119	65
rect	118	65	119	66
rect	118	67	119	68
rect	118	68	119	69
rect	118	69	119	70
rect	118	70	119	71
rect	118	71	119	72
rect	118	74	119	75
rect	118	76	119	77
rect	118	77	119	78
rect	118	78	119	79
rect	118	79	119	80
rect	118	80	119	81
rect	118	82	119	83
rect	118	85	119	86
rect	118	86	119	87
rect	118	87	119	88
rect	118	89	119	90
rect	118	90	119	91
rect	118	92	119	93
rect	118	93	119	94
rect	118	95	119	96
rect	118	96	119	97
rect	118	98	119	99
rect	118	99	119	100
rect	118	101	119	102
rect	118	102	119	103
rect	118	103	119	104
rect	118	105	119	106
rect	118	106	119	107
rect	118	107	119	108
rect	118	108	119	109
rect	118	109	119	110
rect	118	111	119	112
rect	118	112	119	113
rect	118	114	119	115
rect	118	115	119	116
rect	118	117	119	118
rect	118	118	119	119
rect	118	119	119	120
rect	118	139	119	140
rect	118	155	119	156
rect	118	156	119	157
rect	118	158	119	159
rect	118	159	119	160
rect	118	161	119	162
rect	118	162	119	163
rect	118	163	119	164
rect	118	164	119	165
rect	118	165	119	166
rect	118	170	119	171
rect	118	171	119	172
rect	118	172	119	173
rect	120	5	121	6
rect	120	6	121	7
rect	120	7	121	8
rect	120	8	121	9
rect	120	9	121	10
rect	120	10	121	11
rect	120	12	121	13
rect	120	13	121	14
rect	120	14	121	15
rect	120	15	121	16
rect	120	42	121	43
rect	120	43	121	44
rect	120	52	121	53
rect	120	55	121	56
rect	120	56	121	57
rect	120	61	121	62
rect	120	62	121	63
rect	120	64	121	65
rect	120	65	121	66
rect	120	67	121	68
rect	120	68	121	69
rect	120	79	121	80
rect	120	80	121	81
rect	120	82	121	83
rect	120	85	121	86
rect	120	86	121	87
rect	120	87	121	88
rect	120	89	121	90
rect	120	90	121	91
rect	120	92	121	93
rect	120	93	121	94
rect	120	95	121	96
rect	120	96	121	97
rect	120	98	121	99
rect	120	99	121	100
rect	120	101	121	102
rect	120	102	121	103
rect	120	103	121	104
rect	120	105	121	106
rect	120	106	121	107
rect	120	107	121	108
rect	120	108	121	109
rect	120	109	121	110
rect	120	111	121	112
rect	120	112	121	113
rect	120	114	121	115
rect	120	115	121	116
rect	120	117	121	118
rect	120	118	121	119
rect	120	119	121	120
rect	120	121	121	122
rect	120	122	121	123
rect	120	123	121	124
rect	120	124	121	125
rect	120	125	121	126
rect	120	127	121	128
rect	120	128	121	129
rect	120	130	121	131
rect	120	131	121	132
rect	120	133	121	134
rect	120	134	121	135
rect	120	136	121	137
rect	120	137	121	138
rect	120	139	121	140
rect	120	140	121	141
rect	120	141	121	142
rect	120	143	121	144
rect	120	144	121	145
rect	120	145	121	146
rect	120	146	121	147
rect	120	147	121	148
rect	120	149	121	150
rect	120	150	121	151
rect	120	152	121	153
rect	120	153	121	154
rect	120	155	121	156
rect	120	156	121	157
rect	120	158	121	159
rect	120	159	121	160
rect	120	165	121	166
rect	120	166	121	167
rect	120	167	121	168
rect	120	168	121	169
rect	120	169	121	170
rect	120	179	121	180
rect	120	180	121	181
rect	120	181	121	182
rect	122	2	123	3
rect	122	3	123	4
rect	122	5	123	6
rect	122	6	123	7
rect	122	12	123	13
rect	122	24	123	25
rect	122	27	123	28
rect	122	29	123	30
rect	122	30	123	31
rect	122	32	123	33
rect	122	33	123	34
rect	122	36	123	37
rect	122	37	123	38
rect	122	39	123	40
rect	122	40	123	41
rect	122	42	123	43
rect	122	43	123	44
rect	122	45	123	46
rect	122	46	123	47
rect	122	48	123	49
rect	122	49	123	50
rect	122	50	123	51
rect	122	52	123	53
rect	122	55	123	56
rect	122	56	123	57
rect	122	61	123	62
rect	122	62	123	63
rect	122	64	123	65
rect	122	65	123	66
rect	122	67	123	68
rect	122	68	123	69
rect	122	70	123	71
rect	122	71	123	72
rect	122	74	123	75
rect	122	76	123	77
rect	122	77	123	78
rect	122	79	123	80
rect	122	80	123	81
rect	122	82	123	83
rect	122	85	123	86
rect	122	86	123	87
rect	122	87	123	88
rect	122	89	123	90
rect	122	90	123	91
rect	122	92	123	93
rect	122	93	123	94
rect	122	95	123	96
rect	122	96	123	97
rect	122	98	123	99
rect	122	99	123	100
rect	122	101	123	102
rect	122	102	123	103
rect	122	103	123	104
rect	122	105	123	106
rect	122	106	123	107
rect	122	107	123	108
rect	122	108	123	109
rect	122	109	123	110
rect	122	111	123	112
rect	122	112	123	113
rect	122	114	123	115
rect	122	115	123	116
rect	122	117	123	118
rect	122	118	123	119
rect	122	119	123	120
rect	122	121	123	122
rect	122	122	123	123
rect	122	123	123	124
rect	122	124	123	125
rect	122	125	123	126
rect	122	127	123	128
rect	122	128	123	129
rect	122	130	123	131
rect	122	131	123	132
rect	122	133	123	134
rect	122	134	123	135
rect	122	136	123	137
rect	122	137	123	138
rect	122	139	123	140
rect	122	140	123	141
rect	122	141	123	142
rect	122	143	123	144
rect	122	144	123	145
rect	122	145	123	146
rect	122	146	123	147
rect	122	147	123	148
rect	122	149	123	150
rect	122	150	123	151
rect	122	152	123	153
rect	122	153	123	154
rect	122	155	123	156
rect	122	156	123	157
rect	122	158	123	159
rect	122	159	123	160
rect	122	160	123	161
rect	122	161	123	162
rect	122	162	123	163
rect	122	163	123	164
rect	122	165	123	166
rect	122	166	123	167
rect	122	167	123	168
rect	122	168	123	169
rect	122	169	123	170
rect	122	171	123	172
rect	122	172	123	173
rect	122	174	123	175
rect	122	175	123	176
rect	122	177	123	178
rect	122	178	123	179
rect	122	179	123	180
rect	122	180	123	181
rect	122	181	123	182
rect	122	183	123	184
rect	122	184	123	185
rect	122	185	123	186
rect	122	186	123	187
rect	122	187	123	188
rect	122	188	123	189
rect	122	189	123	190
rect	122	190	123	191
rect	122	191	123	192
rect	122	192	123	193
rect	124	2	125	3
rect	124	3	125	4
rect	124	5	125	6
rect	124	6	125	7
rect	124	8	125	9
rect	124	9	125	10
rect	124	24	125	25
rect	124	27	125	28
rect	124	29	125	30
rect	124	30	125	31
rect	124	32	125	33
rect	124	33	125	34
rect	124	36	125	37
rect	124	37	125	38
rect	124	39	125	40
rect	124	40	125	41
rect	124	42	125	43
rect	124	43	125	44
rect	124	45	125	46
rect	124	46	125	47
rect	124	48	125	49
rect	124	49	125	50
rect	124	50	125	51
rect	124	52	125	53
rect	124	55	125	56
rect	124	56	125	57
rect	124	61	125	62
rect	124	62	125	63
rect	124	64	125	65
rect	124	65	125	66
rect	124	67	125	68
rect	124	68	125	69
rect	124	70	125	71
rect	124	71	125	72
rect	124	74	125	75
rect	124	76	125	77
rect	124	77	125	78
rect	124	79	125	80
rect	124	80	125	81
rect	124	82	125	83
rect	124	85	125	86
rect	124	86	125	87
rect	124	87	125	88
rect	124	89	125	90
rect	124	90	125	91
rect	124	92	125	93
rect	124	93	125	94
rect	124	95	125	96
rect	124	96	125	97
rect	124	98	125	99
rect	124	99	125	100
rect	124	101	125	102
rect	124	102	125	103
rect	124	103	125	104
rect	124	105	125	106
rect	124	106	125	107
rect	124	107	125	108
rect	124	108	125	109
rect	124	109	125	110
rect	124	111	125	112
rect	124	112	125	113
rect	124	114	125	115
rect	124	115	125	116
rect	124	117	125	118
rect	124	118	125	119
rect	124	119	125	120
rect	124	121	125	122
rect	124	122	125	123
rect	124	123	125	124
rect	124	124	125	125
rect	124	125	125	126
rect	124	127	125	128
rect	124	128	125	129
rect	124	130	125	131
rect	124	131	125	132
rect	124	133	125	134
rect	124	134	125	135
rect	124	136	125	137
rect	124	137	125	138
rect	124	139	125	140
rect	124	140	125	141
rect	124	141	125	142
rect	124	143	125	144
rect	124	144	125	145
rect	124	162	125	163
rect	124	163	125	164
rect	124	165	125	166
rect	124	166	125	167
rect	124	180	125	181
rect	124	181	125	182
rect	124	183	125	184
rect	124	184	125	185
rect	124	185	125	186
rect	124	186	125	187
rect	124	187	125	188
rect	124	188	125	189
rect	124	189	125	190
rect	124	190	125	191
rect	124	191	125	192
rect	124	192	125	193
rect	124	194	125	195
rect	124	195	125	196
rect	124	197	125	198
rect	124	198	125	199
rect	124	199	125	200
rect	124	200	125	201
rect	124	201	125	202
rect	124	202	125	203
rect	124	203	125	204
rect	124	204	125	205
rect	124	205	125	206
rect	124	206	125	207
rect	124	207	125	208
rect	139	98	140	99
rect	139	99	140	100
rect	139	101	140	102
rect	139	102	140	103
rect	139	103	140	104
rect	141	61	142	62
rect	141	62	142	63
rect	141	64	142	65
rect	141	65	142	66
rect	141	67	142	68
rect	141	68	142	69
rect	141	70	142	71
rect	141	71	142	72
rect	141	74	142	75
rect	141	76	142	77
rect	141	77	142	78
rect	141	79	142	80
rect	141	80	142	81
rect	141	82	142	83
rect	141	85	142	86
rect	141	86	142	87
rect	141	87	142	88
rect	141	89	142	90
rect	141	90	142	91
rect	141	91	142	92
rect	141	92	142	93
rect	141	93	142	94
rect	141	95	142	96
rect	141	96	142	97
rect	143	57	144	58
rect	143	61	144	62
rect	143	62	144	63
rect	143	64	144	65
rect	143	65	144	66
rect	143	67	144	68
rect	143	68	144	69
rect	143	70	144	71
rect	143	71	144	72
rect	143	74	144	75
rect	143	76	144	77
rect	143	77	144	78
rect	145	79	146	80
rect	145	80	146	81
rect	145	82	146	83
rect	145	85	146	86
rect	145	86	146	87
rect	145	87	146	88
rect	147	76	148	77
rect	147	77	148	78
rect	147	79	148	80
rect	147	80	148	81
rect	147	82	148	83
rect	147	85	148	86
rect	147	86	148	87
rect	147	87	148	88
rect	147	88	148	89
rect	147	89	148	90
rect	149	74	150	75
rect	149	75	150	76
rect	149	76	150	77
rect	149	77	150	78
rect	149	79	150	80
rect	149	80	150	81
rect	149	82	150	83
rect	149	85	150	86
rect	149	86	150	87
rect	149	107	150	108
rect	149	108	150	109
rect	149	109	150	110
rect	149	111	150	112
rect	149	112	150	113
rect	149	117	150	118
rect	149	118	150	119
rect	151	64	152	65
rect	151	65	152	66
rect	151	67	152	68
rect	151	68	152	69
rect	151	70	152	71
rect	151	71	152	72
rect	151	74	152	75
rect	151	114	152	115
rect	151	115	152	116
rect	151	116	152	117
rect	151	117	152	118
rect	151	118	152	119
rect	151	120	152	121
rect	151	121	152	122
rect	151	122	152	123
rect	151	123	152	124
rect	151	124	152	125
rect	151	125	152	126
rect	151	127	152	128
rect	151	128	152	129
rect	151	130	152	131
rect	151	131	152	132
rect	151	168	152	169
rect	151	169	152	170
rect	151	171	152	172
rect	151	172	152	173
rect	151	174	152	175
rect	151	175	152	176
rect	151	177	152	178
rect	151	178	152	179
rect	151	180	152	181
rect	151	181	152	182
rect	151	183	152	184
rect	151	184	152	185
rect	151	185	152	186
rect	151	187	152	188
rect	151	188	152	189
rect	151	189	152	190
rect	151	190	152	191
rect	151	191	152	192
rect	151	192	152	193
rect	151	194	152	195
rect	151	195	152	196
rect	153	63	154	64
rect	153	64	154	65
rect	153	65	154	66
rect	153	67	154	68
rect	153	68	154	69
rect	153	70	154	71
rect	153	71	154	72
rect	153	74	154	75
rect	153	76	154	77
rect	153	77	154	78
rect	153	79	154	80
rect	153	80	154	81
rect	153	82	154	83
rect	153	101	154	102
rect	153	102	154	103
rect	153	103	154	104
rect	153	104	154	105
rect	153	105	154	106
rect	153	107	154	108
rect	153	108	154	109
rect	153	109	154	110
rect	153	111	154	112
rect	153	112	154	113
rect	153	114	154	115
rect	153	115	154	116
rect	153	168	154	169
rect	153	169	154	170
rect	153	171	154	172
rect	153	172	154	173
rect	153	174	154	175
rect	153	175	154	176
rect	153	177	154	178
rect	153	178	154	179
rect	153	180	154	181
rect	153	181	154	182
rect	155	18	156	19
rect	155	21	156	22
rect	155	24	156	25
rect	155	27	156	28
rect	155	29	156	30
rect	155	30	156	31
rect	155	32	156	33
rect	155	33	156	34
rect	155	34	156	35
rect	155	36	156	37
rect	155	37	156	38
rect	155	38	156	39
rect	155	39	156	40
rect	155	40	156	41
rect	155	55	156	56
rect	155	57	156	58
rect	155	61	156	62
rect	155	63	156	64
rect	155	64	156	65
rect	155	65	156	66
rect	155	67	156	68
rect	155	68	156	69
rect	155	70	156	71
rect	155	71	156	72
rect	155	95	156	96
rect	155	96	156	97
rect	155	98	156	99
rect	155	99	156	100
rect	155	133	156	134
rect	155	134	156	135
rect	155	146	156	147
rect	155	147	156	148
rect	155	177	156	178
rect	155	178	156	179
rect	155	180	156	181
rect	155	181	156	182
rect	155	182	156	183
rect	157	8	158	9
rect	157	9	158	10
rect	157	11	158	12
rect	157	12	158	13
rect	157	14	158	15
rect	157	15	158	16
rect	157	39	158	40
rect	157	40	158	41
rect	157	41	158	42
rect	157	42	158	43
rect	157	43	158	44
rect	157	45	158	46
rect	157	46	158	47
rect	157	51	158	52
rect	157	52	158	53
rect	157	55	158	56
rect	157	57	158	58
rect	157	61	158	62
rect	157	63	158	64
rect	157	64	158	65
rect	157	65	158	66
rect	157	67	158	68
rect	157	68	158	69
rect	157	85	158	86
rect	157	86	158	87
rect	157	88	158	89
rect	157	89	158	90
rect	157	91	158	92
rect	157	92	158	93
rect	157	93	158	94
rect	157	94	158	95
rect	157	95	158	96
rect	157	96	158	97
rect	157	98	158	99
rect	157	99	158	100
rect	157	101	158	102
rect	157	102	158	103
rect	157	103	158	104
rect	157	104	158	105
rect	157	105	158	106
rect	157	107	158	108
rect	157	108	158	109
rect	157	109	158	110
rect	157	111	158	112
rect	157	112	158	113
rect	157	114	158	115
rect	157	115	158	116
rect	157	117	158	118
rect	157	118	158	119
rect	157	120	158	121
rect	157	121	158	122
rect	157	122	158	123
rect	157	123	158	124
rect	157	124	158	125
rect	157	125	158	126
rect	157	127	158	128
rect	157	128	158	129
rect	157	130	158	131
rect	157	131	158	132
rect	157	133	158	134
rect	157	134	158	135
rect	157	135	158	136
rect	157	136	158	137
rect	157	137	158	138
rect	157	139	158	140
rect	157	140	158	141
rect	157	141	158	142
rect	157	142	158	143
rect	157	143	158	144
rect	157	144	158	145
rect	157	145	158	146
rect	157	146	158	147
rect	157	147	158	148
rect	157	148	158	149
rect	157	149	158	150
rect	157	150	158	151
rect	157	152	158	153
rect	157	153	158	154
rect	157	155	158	156
rect	157	156	158	157
rect	157	158	158	159
rect	157	159	158	160
rect	157	160	158	161
rect	157	162	158	163
rect	157	163	158	164
rect	157	165	158	166
rect	157	166	158	167
rect	157	168	158	169
rect	157	169	158	170
rect	157	171	158	172
rect	157	172	158	173
rect	157	174	158	175
rect	157	175	158	176
rect	157	176	158	177
rect	159	8	160	9
rect	159	9	160	10
rect	159	11	160	12
rect	159	12	160	13
rect	159	14	160	15
rect	159	15	160	16
rect	159	18	160	19
rect	159	32	160	33
rect	159	33	160	34
rect	159	34	160	35
rect	159	36	160	37
rect	159	37	160	38
rect	159	39	160	40
rect	159	40	160	41
rect	159	48	160	49
rect	159	49	160	50
rect	159	51	160	52
rect	159	52	160	53
rect	159	55	160	56
rect	159	57	160	58
rect	159	82	160	83
rect	159	85	160	86
rect	159	86	160	87
rect	159	88	160	89
rect	159	89	160	90
rect	159	91	160	92
rect	159	92	160	93
rect	159	93	160	94
rect	159	94	160	95
rect	159	95	160	96
rect	159	96	160	97
rect	159	98	160	99
rect	159	99	160	100
rect	159	101	160	102
rect	159	102	160	103
rect	159	103	160	104
rect	159	104	160	105
rect	159	105	160	106
rect	159	107	160	108
rect	159	108	160	109
rect	159	109	160	110
rect	159	111	160	112
rect	159	112	160	113
rect	159	114	160	115
rect	159	115	160	116
rect	159	117	160	118
rect	159	118	160	119
rect	159	120	160	121
rect	159	121	160	122
rect	159	122	160	123
rect	159	123	160	124
rect	159	124	160	125
rect	159	125	160	126
rect	159	127	160	128
rect	159	128	160	129
rect	159	130	160	131
rect	159	131	160	132
rect	159	133	160	134
rect	159	134	160	135
rect	159	135	160	136
rect	159	136	160	137
rect	159	137	160	138
rect	159	139	160	140
rect	159	140	160	141
rect	159	141	160	142
rect	159	142	160	143
rect	159	143	160	144
rect	159	144	160	145
rect	159	145	160	146
rect	159	146	160	147
rect	159	147	160	148
rect	159	148	160	149
rect	159	149	160	150
rect	159	150	160	151
rect	159	152	160	153
rect	159	153	160	154
rect	159	155	160	156
rect	159	156	160	157
rect	159	158	160	159
rect	159	159	160	160
rect	159	160	160	161
rect	161	5	162	6
rect	161	6	162	7
rect	161	8	162	9
rect	161	9	162	10
rect	161	14	162	15
rect	161	15	162	16
rect	161	18	162	19
rect	161	33	162	34
rect	161	34	162	35
rect	161	36	162	37
rect	161	37	162	38
rect	161	39	162	40
rect	161	40	162	41
rect	161	42	162	43
rect	161	43	162	44
rect	161	45	162	46
rect	161	46	162	47
rect	161	48	162	49
rect	161	49	162	50
rect	161	51	162	52
rect	161	52	162	53
rect	161	55	162	56
rect	161	57	162	58
rect	161	60	162	61
rect	161	61	162	62
rect	161	63	162	64
rect	161	64	162	65
rect	161	65	162	66
rect	161	67	162	68
rect	161	68	162	69
rect	161	69	162	70
rect	161	70	162	71
rect	161	71	162	72
rect	161	74	162	75
rect	161	76	162	77
rect	161	77	162	78
rect	161	79	162	80
rect	161	80	162	81
rect	161	81	162	82
rect	161	82	162	83
rect	161	85	162	86
rect	161	86	162	87
rect	161	88	162	89
rect	161	89	162	90
rect	161	91	162	92
rect	161	92	162	93
rect	161	93	162	94
rect	161	94	162	95
rect	161	95	162	96
rect	161	96	162	97
rect	161	98	162	99
rect	161	99	162	100
rect	161	101	162	102
rect	161	102	162	103
rect	161	136	162	137
rect	161	137	162	138
rect	161	149	162	150
rect	161	150	162	151
rect	163	11	164	12
rect	163	12	164	13
rect	163	13	164	14
rect	163	14	164	15
rect	163	15	164	16
rect	163	18	164	19
rect	163	21	164	22
rect	163	29	164	30
rect	163	30	164	31
rect	163	31	164	32
rect	163	33	164	34
rect	163	34	164	35
rect	163	36	164	37
rect	163	37	164	38
rect	163	39	164	40
rect	163	40	164	41
rect	163	42	164	43
rect	163	43	164	44
rect	163	45	164	46
rect	163	46	164	47
rect	163	48	164	49
rect	163	49	164	50
rect	163	51	164	52
rect	163	52	164	53
rect	163	60	164	61
rect	163	61	164	62
rect	163	63	164	64
rect	163	64	164	65
rect	163	65	164	66
rect	163	82	164	83
rect	163	85	164	86
rect	163	86	164	87
rect	163	88	164	89
rect	163	89	164	90
rect	163	91	164	92
rect	163	92	164	93
rect	163	93	164	94
rect	163	94	164	95
rect	163	95	164	96
rect	163	96	164	97
rect	163	98	164	99
rect	163	99	164	100
rect	163	101	164	102
rect	163	102	164	103
rect	163	104	164	105
rect	163	105	164	106
rect	163	107	164	108
rect	163	108	164	109
rect	163	109	164	110
rect	163	111	164	112
rect	163	112	164	113
rect	163	114	164	115
rect	163	115	164	116
rect	163	117	164	118
rect	163	118	164	119
rect	163	120	164	121
rect	163	121	164	122
rect	163	122	164	123
rect	163	123	164	124
rect	163	124	164	125
rect	163	125	164	126
rect	163	127	164	128
rect	163	128	164	129
rect	163	130	164	131
rect	163	131	164	132
rect	163	133	164	134
rect	163	134	164	135
rect	163	136	164	137
rect	163	137	164	138
rect	163	138	164	139
rect	163	139	164	140
rect	163	140	164	141
rect	163	141	164	142
rect	163	142	164	143
rect	163	143	164	144
rect	163	144	164	145
rect	163	145	164	146
rect	163	146	164	147
rect	163	147	164	148
rect	163	149	164	150
rect	163	150	164	151
rect	163	151	164	152
rect	163	152	164	153
rect	163	153	164	154
rect	163	155	164	156
rect	163	156	164	157
rect	163	158	164	159
rect	163	159	164	160
rect	163	160	164	161
rect	163	161	164	162
rect	163	162	164	163
rect	163	163	164	164
rect	163	165	164	166
rect	163	166	164	167
rect	163	168	164	169
rect	163	169	164	170
rect	163	171	164	172
rect	163	172	164	173
rect	163	174	164	175
rect	163	175	164	176
rect	163	176	164	177
rect	163	178	164	179
rect	163	180	164	181
rect	163	181	164	182
rect	163	182	164	183
rect	163	184	164	185
rect	163	185	164	186
rect	163	187	164	188
rect	163	188	164	189
rect	163	189	164	190
rect	163	190	164	191
rect	163	191	164	192
rect	163	192	164	193
rect	165	5	166	6
rect	165	6	166	7
rect	165	8	166	9
rect	165	9	166	10
rect	165	11	166	12
rect	165	12	166	13
rect	165	13	166	14
rect	165	14	166	15
rect	165	15	166	16
rect	165	18	166	19
rect	165	21	166	22
rect	165	24	166	25
rect	165	27	166	28
rect	165	28	166	29
rect	165	29	166	30
rect	165	30	166	31
rect	165	31	166	32
rect	165	33	166	34
rect	165	34	166	35
rect	165	36	166	37
rect	165	37	166	38
rect	165	39	166	40
rect	165	40	166	41
rect	165	42	166	43
rect	165	43	166	44
rect	165	45	166	46
rect	165	46	166	47
rect	165	48	166	49
rect	165	49	166	50
rect	165	51	166	52
rect	165	52	166	53
rect	165	55	166	56
rect	165	57	166	58
rect	165	60	166	61
rect	165	61	166	62
rect	165	63	166	64
rect	165	64	166	65
rect	165	65	166	66
rect	165	66	166	67
rect	165	67	166	68
rect	165	68	166	69
rect	165	69	166	70
rect	165	70	166	71
rect	165	71	166	72
rect	165	74	166	75
rect	165	76	166	77
rect	165	77	166	78
rect	165	79	166	80
rect	165	80	166	81
rect	165	82	166	83
rect	165	85	166	86
rect	165	86	166	87
rect	165	88	166	89
rect	165	89	166	90
rect	165	91	166	92
rect	165	92	166	93
rect	165	93	166	94
rect	165	94	166	95
rect	165	95	166	96
rect	165	96	166	97
rect	165	98	166	99
rect	165	99	166	100
rect	165	101	166	102
rect	165	102	166	103
rect	165	104	166	105
rect	165	105	166	106
rect	165	107	166	108
rect	165	108	166	109
rect	165	109	166	110
rect	165	111	166	112
rect	165	112	166	113
rect	165	114	166	115
rect	165	115	166	116
rect	165	117	166	118
rect	165	118	166	119
rect	165	120	166	121
rect	165	121	166	122
rect	165	122	166	123
rect	165	123	166	124
rect	165	124	166	125
rect	165	125	166	126
rect	165	127	166	128
rect	165	128	166	129
rect	165	130	166	131
rect	165	131	166	132
rect	165	133	166	134
rect	165	134	166	135
rect	165	136	166	137
rect	165	137	166	138
rect	165	138	166	139
rect	165	139	166	140
rect	165	140	166	141
rect	165	141	166	142
rect	165	142	166	143
rect	165	143	166	144
rect	165	144	166	145
rect	165	145	166	146
rect	165	146	166	147
rect	165	147	166	148
rect	165	149	166	150
rect	165	150	166	151
rect	165	155	166	156
rect	165	156	166	157
rect	165	158	166	159
rect	165	159	166	160
rect	165	160	166	161
rect	165	161	166	162
rect	165	162	166	163
rect	165	163	166	164
rect	165	171	166	172
rect	165	172	166	173
rect	165	174	166	175
rect	165	175	166	176
rect	165	176	166	177
rect	165	178	166	179
rect	165	180	166	181
rect	165	181	166	182
rect	165	182	166	183
rect	165	184	166	185
rect	165	185	166	186
rect	167	2	168	3
rect	167	3	168	4
rect	167	5	168	6
rect	167	6	168	7
rect	167	8	168	9
rect	167	9	168	10
rect	167	11	168	12
rect	167	12	168	13
rect	167	13	168	14
rect	167	14	168	15
rect	167	15	168	16
rect	167	18	168	19
rect	167	21	168	22
rect	167	24	168	25
rect	167	27	168	28
rect	167	28	168	29
rect	167	29	168	30
rect	167	30	168	31
rect	167	31	168	32
rect	167	33	168	34
rect	167	34	168	35
rect	167	36	168	37
rect	167	37	168	38
rect	167	39	168	40
rect	167	40	168	41
rect	167	42	168	43
rect	167	43	168	44
rect	167	45	168	46
rect	167	46	168	47
rect	167	48	168	49
rect	167	49	168	50
rect	167	51	168	52
rect	167	52	168	53
rect	167	55	168	56
rect	167	57	168	58
rect	167	60	168	61
rect	167	61	168	62
rect	167	63	168	64
rect	167	64	168	65
rect	167	65	168	66
rect	167	66	168	67
rect	167	67	168	68
rect	167	68	168	69
rect	167	69	168	70
rect	167	70	168	71
rect	167	71	168	72
rect	167	74	168	75
rect	167	76	168	77
rect	167	77	168	78
rect	167	79	168	80
rect	167	80	168	81
rect	167	82	168	83
rect	167	85	168	86
rect	167	86	168	87
rect	167	88	168	89
rect	167	89	168	90
rect	167	91	168	92
rect	167	92	168	93
rect	167	93	168	94
rect	167	94	168	95
rect	167	95	168	96
rect	167	96	168	97
rect	167	98	168	99
rect	167	99	168	100
rect	167	101	168	102
rect	167	102	168	103
rect	167	104	168	105
rect	167	105	168	106
rect	167	107	168	108
rect	167	108	168	109
rect	167	109	168	110
rect	167	127	168	128
rect	167	128	168	129
rect	167	130	168	131
rect	167	131	168	132
rect	167	133	168	134
rect	167	134	168	135
rect	167	136	168	137
rect	167	137	168	138
rect	167	138	168	139
rect	167	139	168	140
rect	167	140	168	141
rect	167	141	168	142
rect	167	142	168	143
rect	167	143	168	144
rect	167	144	168	145
rect	167	155	168	156
rect	167	156	168	157
rect	167	158	168	159
rect	167	159	168	160
rect	167	160	168	161
rect	167	161	168	162
rect	167	162	168	163
rect	167	163	168	164
rect	167	164	168	165
rect	167	165	168	166
rect	167	166	168	167
rect	167	168	168	169
rect	167	169	168	170
rect	167	170	168	171
rect	167	171	168	172
rect	167	172	168	173
rect	167	174	168	175
rect	167	175	168	176
rect	167	176	168	177
rect	167	178	168	179
rect	169	2	170	3
rect	169	3	170	4
rect	169	5	170	6
rect	169	6	170	7
rect	169	8	170	9
rect	169	9	170	10
rect	169	11	170	12
rect	169	12	170	13
rect	169	24	170	25
rect	169	27	170	28
rect	169	28	170	29
rect	169	29	170	30
rect	169	30	170	31
rect	169	31	170	32
rect	169	33	170	34
rect	169	34	170	35
rect	169	36	170	37
rect	169	37	170	38
rect	169	39	170	40
rect	169	40	170	41
rect	169	42	170	43
rect	169	43	170	44
rect	169	45	170	46
rect	169	46	170	47
rect	169	48	170	49
rect	169	49	170	50
rect	169	51	170	52
rect	169	52	170	53
rect	169	55	170	56
rect	169	57	170	58
rect	169	60	170	61
rect	169	61	170	62
rect	169	63	170	64
rect	169	64	170	65
rect	169	65	170	66
rect	169	66	170	67
rect	169	67	170	68
rect	169	68	170	69
rect	169	69	170	70
rect	169	70	170	71
rect	169	71	170	72
rect	169	74	170	75
rect	169	76	170	77
rect	169	77	170	78
rect	169	79	170	80
rect	169	80	170	81
rect	169	82	170	83
rect	169	85	170	86
rect	169	86	170	87
rect	169	88	170	89
rect	169	89	170	90
rect	169	91	170	92
rect	169	92	170	93
rect	169	93	170	94
rect	169	94	170	95
rect	169	95	170	96
rect	169	96	170	97
rect	169	98	170	99
rect	169	99	170	100
rect	169	101	170	102
rect	169	102	170	103
rect	169	104	170	105
rect	169	105	170	106
rect	169	107	170	108
rect	169	108	170	109
rect	169	109	170	110
rect	169	110	170	111
rect	169	111	170	112
rect	169	112	170	113
rect	169	114	170	115
rect	169	115	170	116
rect	169	117	170	118
rect	169	118	170	119
rect	169	120	170	121
rect	169	121	170	122
rect	169	122	170	123
rect	169	127	170	128
rect	169	128	170	129
rect	169	130	170	131
rect	169	131	170	132
rect	169	133	170	134
rect	169	134	170	135
rect	169	136	170	137
rect	169	137	170	138
rect	169	138	170	139
rect	169	139	170	140
rect	169	140	170	141
rect	169	141	170	142
rect	169	142	170	143
rect	169	143	170	144
rect	169	144	170	145
rect	169	146	170	147
rect	169	147	170	148
rect	169	149	170	150
rect	169	150	170	151
rect	169	152	170	153
rect	169	153	170	154
rect	169	155	170	156
rect	169	156	170	157
rect	169	158	170	159
rect	169	159	170	160
rect	169	160	170	161
rect	169	161	170	162
rect	169	162	170	163
rect	169	163	170	164
rect	169	164	170	165
rect	169	165	170	166
rect	169	166	170	167
rect	169	168	170	169
rect	169	169	170	170
rect	169	174	170	175
rect	169	175	170	176
rect	169	176	170	177
rect	169	178	170	179
rect	169	179	170	180
rect	194	65	195	66
rect	194	66	195	67
rect	194	67	195	68
rect	194	68	195	69
rect	194	70	195	71
rect	194	71	195	72
rect	194	72	195	73
rect	194	74	195	75
rect	196	77	197	78
rect	196	79	197	80
rect	196	80	197	81
rect	196	82	197	83
rect	196	84	197	85
rect	196	85	197	86
rect	196	86	197	87
rect	196	88	197	89
rect	196	89	197	90
rect	198	68	199	69
rect	198	70	199	71
rect	198	71	199	72
rect	198	72	199	73
rect	198	74	199	75
rect	198	75	199	76
rect	198	77	199	78
rect	198	95	199	96
rect	198	96	199	97
rect	198	97	199	98
rect	198	98	199	99
rect	198	99	199	100
rect	200	63	201	64
rect	200	65	201	66
rect	200	66	201	67
rect	200	68	201	69
rect	200	70	201	71
rect	200	71	201	72
rect	200	72	201	73
rect	200	74	201	75
rect	200	75	201	76
rect	200	77	201	78
rect	200	78	201	79
rect	200	93	201	94
rect	200	94	201	95
rect	200	95	201	96
rect	200	96	201	97
rect	200	97	201	98
rect	200	98	201	99
rect	200	99	201	100
rect	200	100	201	101
rect	200	101	201	102
rect	200	102	201	103
rect	200	104	201	105
rect	200	105	201	106
rect	202	62	203	63
rect	202	63	203	64
rect	202	65	203	66
rect	202	66	203	67
rect	202	68	203	69
rect	202	70	203	71
rect	202	71	203	72
rect	202	72	203	73
rect	202	74	203	75
rect	202	75	203	76
rect	202	77	203	78
rect	202	78	203	79
rect	202	80	203	81
rect	202	82	203	83
rect	202	84	203	85
rect	202	85	203	86
rect	202	86	203	87
rect	202	88	203	89
rect	202	89	203	90
rect	202	90	203	91
rect	202	91	203	92
rect	202	93	203	94
rect	202	94	203	95
rect	202	95	203	96
rect	202	96	203	97
rect	202	97	203	98
rect	202	98	203	99
rect	202	99	203	100
rect	202	100	203	101
rect	202	101	203	102
rect	202	102	203	103
rect	202	104	203	105
rect	202	105	203	106
rect	202	106	203	107
rect	202	107	203	108
rect	202	108	203	109
rect	202	109	203	110
rect	202	110	203	111
rect	202	111	203	112
rect	202	112	203	113
rect	202	113	203	114
rect	202	114	203	115
rect	202	115	203	116
rect	202	122	203	123
rect	202	124	203	125
rect	202	125	203	126
rect	202	126	203	127
rect	202	127	203	128
rect	202	128	203	129
rect	202	130	203	131
rect	202	131	203	132
rect	204	30	205	31
rect	204	31	205	32
rect	204	33	205	34
rect	204	34	205	35
rect	204	36	205	37
rect	204	37	205	38
rect	204	45	205	46
rect	204	46	205	47
rect	204	48	205	49
rect	204	49	205	50
rect	204	51	205	52
rect	204	52	205	53
rect	204	53	205	54
rect	204	55	205	56
rect	204	57	205	58
rect	204	59	205	60
rect	204	60	205	61
rect	204	62	205	63
rect	204	63	205	64
rect	204	65	205	66
rect	204	66	205	67
rect	204	68	205	69
rect	204	70	205	71
rect	204	71	205	72
rect	204	72	205	73
rect	204	74	205	75
rect	204	75	205	76
rect	204	77	205	78
rect	204	78	205	79
rect	204	80	205	81
rect	204	82	205	83
rect	204	84	205	85
rect	204	85	205	86
rect	204	86	205	87
rect	204	88	205	89
rect	204	89	205	90
rect	204	90	205	91
rect	204	91	205	92
rect	204	93	205	94
rect	204	94	205	95
rect	204	95	205	96
rect	204	96	205	97
rect	204	97	205	98
rect	204	98	205	99
rect	204	99	205	100
rect	204	100	205	101
rect	204	101	205	102
rect	204	102	205	103
rect	204	104	205	105
rect	204	105	205	106
rect	204	106	205	107
rect	204	107	205	108
rect	204	108	205	109
rect	204	109	205	110
rect	204	110	205	111
rect	204	111	205	112
rect	204	112	205	113
rect	204	113	205	114
rect	204	114	205	115
rect	204	115	205	116
rect	204	116	205	117
rect	204	117	205	118
rect	204	118	205	119
rect	204	120	205	121
rect	204	122	205	123
rect	204	124	205	125
rect	204	125	205	126
rect	204	126	205	127
rect	204	127	205	128
rect	204	128	205	129
rect	204	130	205	131
rect	204	146	205	147
rect	204	147	205	148
rect	204	149	205	150
rect	204	150	205	151
rect	204	152	205	153
rect	204	153	205	154
rect	204	155	205	156
rect	204	156	205	157
rect	204	158	205	159
rect	204	159	205	160
rect	204	160	205	161
rect	204	161	205	162
rect	204	162	205	163
rect	204	163	205	164
rect	206	40	207	41
rect	206	46	207	47
rect	206	48	207	49
rect	206	49	207	50
rect	206	70	207	71
rect	206	71	207	72
rect	206	72	207	73
rect	206	74	207	75
rect	206	75	207	76
rect	206	77	207	78
rect	206	78	207	79
rect	206	80	207	81
rect	206	82	207	83
rect	206	84	207	85
rect	206	85	207	86
rect	206	86	207	87
rect	206	88	207	89
rect	206	89	207	90
rect	206	90	207	91
rect	206	91	207	92
rect	206	93	207	94
rect	206	94	207	95
rect	206	95	207	96
rect	206	96	207	97
rect	206	97	207	98
rect	206	98	207	99
rect	206	106	207	107
rect	206	107	207	108
rect	206	108	207	109
rect	206	109	207	110
rect	206	110	207	111
rect	206	111	207	112
rect	206	112	207	113
rect	206	113	207	114
rect	206	114	207	115
rect	206	147	207	148
rect	206	149	207	150
rect	206	150	207	151
rect	206	152	207	153
rect	206	153	207	154
rect	206	155	207	156
rect	206	156	207	157
rect	208	33	209	34
rect	208	34	209	35
rect	208	43	209	44
rect	208	44	209	45
rect	208	46	209	47
rect	208	48	209	49
rect	208	49	209	50
rect	208	50	209	51
rect	208	51	209	52
rect	208	52	209	53
rect	208	53	209	54
rect	208	55	209	56
rect	208	57	209	58
rect	208	59	209	60
rect	208	60	209	61
rect	208	62	209	63
rect	208	63	209	64
rect	208	65	209	66
rect	208	66	209	67
rect	208	68	209	69
rect	208	69	209	70
rect	208	70	209	71
rect	208	71	209	72
rect	208	72	209	73
rect	208	74	209	75
rect	208	75	209	76
rect	208	77	209	78
rect	208	78	209	79
rect	208	80	209	81
rect	208	82	209	83
rect	208	84	209	85
rect	208	85	209	86
rect	208	86	209	87
rect	208	88	209	89
rect	208	89	209	90
rect	208	90	209	91
rect	208	91	209	92
rect	208	93	209	94
rect	208	94	209	95
rect	208	95	209	96
rect	208	96	209	97
rect	208	97	209	98
rect	208	98	209	99
rect	208	100	209	101
rect	208	101	209	102
rect	208	102	209	103
rect	208	104	209	105
rect	208	106	209	107
rect	208	107	209	108
rect	208	108	209	109
rect	208	109	209	110
rect	208	110	209	111
rect	208	111	209	112
rect	208	112	209	113
rect	208	113	209	114
rect	208	114	209	115
rect	208	116	209	117
rect	208	117	209	118
rect	208	118	209	119
rect	208	120	209	121
rect	208	122	209	123
rect	208	128	209	129
rect	208	130	209	131
rect	208	132	209	133
rect	208	133	209	134
rect	208	134	209	135
rect	208	144	209	145
rect	208	145	209	146
rect	208	147	209	148
rect	208	149	209	150
rect	208	150	209	151
rect	208	152	209	153
rect	208	153	209	154
rect	210	30	211	31
rect	210	31	211	32
rect	210	32	211	33
rect	210	33	211	34
rect	210	34	211	35
rect	210	35	211	36
rect	210	36	211	37
rect	210	37	211	38
rect	210	38	211	39
rect	210	40	211	41
rect	210	41	211	42
rect	210	43	211	44
rect	210	44	211	45
rect	210	46	211	47
rect	210	52	211	53
rect	210	53	211	54
rect	210	55	211	56
rect	210	71	211	72
rect	210	72	211	73
rect	210	74	211	75
rect	210	75	211	76
rect	210	77	211	78
rect	210	78	211	79
rect	210	80	211	81
rect	210	90	211	91
rect	210	91	211	92
rect	210	93	211	94
rect	210	94	211	95
rect	210	95	211	96
rect	210	96	211	97
rect	210	97	211	98
rect	210	98	211	99
rect	210	100	211	101
rect	210	101	211	102
rect	210	102	211	103
rect	210	109	211	110
rect	210	110	211	111
rect	210	111	211	112
rect	210	112	211	113
rect	210	113	211	114
rect	210	114	211	115
rect	210	116	211	117
rect	210	117	211	118
rect	210	118	211	119
rect	210	125	211	126
rect	210	126	211	127
rect	210	128	211	129
rect	210	130	211	131
rect	210	132	211	133
rect	210	133	211	134
rect	210	134	211	135
rect	210	135	211	136
rect	210	136	211	137
rect	210	137	211	138
rect	210	138	211	139
rect	210	139	211	140
rect	210	140	211	141
rect	210	141	211	142
rect	210	142	211	143
rect	210	144	211	145
rect	210	145	211	146
rect	210	147	211	148
rect	210	154	211	155
rect	210	155	211	156
rect	210	156	211	157
rect	210	157	211	158
rect	210	158	211	159
rect	212	5	213	6
rect	212	6	213	7
rect	212	27	213	28
rect	212	28	213	29
rect	212	30	213	31
rect	212	31	213	32
rect	212	32	213	33
rect	212	49	213	50
rect	212	50	213	51
rect	212	52	213	53
rect	212	53	213	54
rect	212	55	213	56
rect	212	56	213	57
rect	212	57	213	58
rect	212	59	213	60
rect	212	60	213	61
rect	212	62	213	63
rect	212	63	213	64
rect	212	65	213	66
rect	212	66	213	67
rect	212	68	213	69
rect	212	69	213	70
rect	212	71	213	72
rect	212	72	213	73
rect	212	74	213	75
rect	212	75	213	76
rect	212	77	213	78
rect	212	78	213	79
rect	212	80	213	81
rect	212	81	213	82
rect	212	82	213	83
rect	212	84	213	85
rect	212	85	213	86
rect	212	86	213	87
rect	212	96	213	97
rect	212	97	213	98
rect	212	98	213	99
rect	212	100	213	101
rect	212	101	213	102
rect	212	102	213	103
rect	212	103	213	104
rect	212	104	213	105
rect	212	106	213	107
rect	212	107	213	108
rect	212	109	213	110
rect	212	110	213	111
rect	212	111	213	112
rect	212	112	213	113
rect	212	113	213	114
rect	212	114	213	115
rect	212	116	213	117
rect	212	117	213	118
rect	212	118	213	119
rect	212	119	213	120
rect	212	120	213	121
rect	212	122	213	123
rect	212	123	213	124
rect	212	125	213	126
rect	212	126	213	127
rect	212	128	213	129
rect	212	130	213	131
rect	212	132	213	133
rect	212	133	213	134
rect	212	141	213	142
rect	212	142	213	143
rect	212	144	213	145
rect	212	145	213	146
rect	212	147	213	148
rect	212	148	213	149
rect	212	149	213	150
rect	212	150	213	151
rect	212	163	213	164
rect	212	164	213	165
rect	212	165	213	166
rect	212	166	213	167
rect	212	168	213	169
rect	212	169	213	170
rect	214	9	215	10
rect	214	11	215	12
rect	214	12	215	13
rect	214	14	215	15
rect	214	15	215	16
rect	214	16	215	17
rect	214	18	215	19
rect	214	19	215	20
rect	214	21	215	22
rect	214	22	215	23
rect	214	24	215	25
rect	214	25	215	26
rect	214	27	215	28
rect	214	28	215	29
rect	214	30	215	31
rect	214	31	215	32
rect	214	32	215	33
rect	214	34	215	35
rect	214	35	215	36
rect	214	36	215	37
rect	214	37	215	38
rect	214	38	215	39
rect	214	40	215	41
rect	214	41	215	42
rect	214	43	215	44
rect	214	44	215	45
rect	214	46	215	47
rect	214	47	215	48
rect	214	49	215	50
rect	214	50	215	51
rect	214	52	215	53
rect	214	53	215	54
rect	214	55	215	56
rect	214	56	215	57
rect	214	57	215	58
rect	214	59	215	60
rect	214	60	215	61
rect	214	62	215	63
rect	214	63	215	64
rect	214	65	215	66
rect	214	66	215	67
rect	214	68	215	69
rect	214	69	215	70
rect	214	71	215	72
rect	214	72	215	73
rect	214	74	215	75
rect	214	75	215	76
rect	214	77	215	78
rect	214	78	215	79
rect	214	80	215	81
rect	214	81	215	82
rect	214	82	215	83
rect	214	84	215	85
rect	214	85	215	86
rect	214	86	215	87
rect	214	87	215	88
rect	214	88	215	89
rect	214	90	215	91
rect	214	91	215	92
rect	214	93	215	94
rect	214	94	215	95
rect	214	96	215	97
rect	214	97	215	98
rect	214	98	215	99
rect	214	100	215	101
rect	214	101	215	102
rect	214	102	215	103
rect	214	103	215	104
rect	214	104	215	105
rect	214	106	215	107
rect	214	107	215	108
rect	214	109	215	110
rect	214	110	215	111
rect	214	111	215	112
rect	214	112	215	113
rect	214	113	215	114
rect	214	114	215	115
rect	214	116	215	117
rect	214	117	215	118
rect	214	118	215	119
rect	214	119	215	120
rect	214	120	215	121
rect	214	122	215	123
rect	214	123	215	124
rect	214	125	215	126
rect	214	126	215	127
rect	214	128	215	129
rect	214	130	215	131
rect	214	132	215	133
rect	214	133	215	134
rect	214	135	215	136
rect	214	136	215	137
rect	214	137	215	138
rect	214	138	215	139
rect	214	139	215	140
rect	214	141	215	142
rect	214	142	215	143
rect	214	144	215	145
rect	214	145	215	146
rect	214	147	215	148
rect	214	148	215	149
rect	214	149	215	150
rect	214	150	215	151
rect	214	151	215	152
rect	214	152	215	153
rect	214	154	215	155
rect	214	155	215	156
rect	214	156	215	157
rect	214	157	215	158
rect	214	158	215	159
rect	214	160	215	161
rect	214	161	215	162
rect	214	163	215	164
rect	214	164	215	165
rect	214	165	215	166
rect	214	166	215	167
rect	214	168	215	169
rect	216	2	217	3
rect	216	3	217	4
rect	216	5	217	6
rect	216	6	217	7
rect	216	7	217	8
rect	216	9	217	10
rect	216	11	217	12
rect	216	12	217	13
rect	216	14	217	15
rect	216	15	217	16
rect	216	16	217	17
rect	216	18	217	19
rect	216	19	217	20
rect	216	21	217	22
rect	216	22	217	23
rect	216	24	217	25
rect	216	25	217	26
rect	216	27	217	28
rect	216	28	217	29
rect	216	30	217	31
rect	216	31	217	32
rect	216	32	217	33
rect	216	34	217	35
rect	216	35	217	36
rect	216	36	217	37
rect	216	37	217	38
rect	216	38	217	39
rect	216	40	217	41
rect	216	41	217	42
rect	216	43	217	44
rect	216	44	217	45
rect	216	46	217	47
rect	216	47	217	48
rect	216	49	217	50
rect	216	50	217	51
rect	216	52	217	53
rect	216	53	217	54
rect	216	55	217	56
rect	216	56	217	57
rect	216	57	217	58
rect	216	59	217	60
rect	216	60	217	61
rect	216	62	217	63
rect	216	63	217	64
rect	216	65	217	66
rect	216	66	217	67
rect	216	68	217	69
rect	216	69	217	70
rect	216	71	217	72
rect	216	72	217	73
rect	216	74	217	75
rect	216	75	217	76
rect	216	77	217	78
rect	216	78	217	79
rect	216	80	217	81
rect	216	81	217	82
rect	216	82	217	83
rect	216	84	217	85
rect	216	85	217	86
rect	216	86	217	87
rect	216	87	217	88
rect	216	88	217	89
rect	216	90	217	91
rect	216	91	217	92
rect	216	93	217	94
rect	216	94	217	95
rect	216	96	217	97
rect	216	97	217	98
rect	216	98	217	99
rect	216	100	217	101
rect	216	101	217	102
rect	216	102	217	103
rect	216	103	217	104
rect	216	104	217	105
rect	216	106	217	107
rect	216	107	217	108
rect	216	109	217	110
rect	216	110	217	111
rect	216	111	217	112
rect	216	112	217	113
rect	216	113	217	114
rect	216	114	217	115
rect	216	116	217	117
rect	216	117	217	118
rect	216	118	217	119
rect	216	119	217	120
rect	216	120	217	121
rect	216	122	217	123
rect	216	123	217	124
rect	216	125	217	126
rect	216	126	217	127
rect	216	128	217	129
rect	216	130	217	131
rect	216	132	217	133
rect	216	133	217	134
rect	216	135	217	136
rect	216	136	217	137
rect	216	137	217	138
rect	216	138	217	139
rect	216	139	217	140
rect	216	141	217	142
rect	216	142	217	143
rect	216	144	217	145
rect	216	145	217	146
rect	216	147	217	148
rect	216	148	217	149
rect	216	149	217	150
rect	216	150	217	151
rect	216	151	217	152
rect	216	152	217	153
rect	216	154	217	155
rect	216	155	217	156
rect	216	184	217	185
rect	216	185	217	186
rect	216	186	217	187
rect	216	188	217	189
rect	216	189	217	190
rect	218	2	219	3
rect	218	3	219	4
rect	218	5	219	6
rect	218	6	219	7
rect	218	7	219	8
rect	218	9	219	10
rect	218	27	219	28
rect	218	28	219	29
rect	218	30	219	31
rect	218	31	219	32
rect	218	32	219	33
rect	218	34	219	35
rect	218	35	219	36
rect	218	36	219	37
rect	218	37	219	38
rect	218	38	219	39
rect	218	40	219	41
rect	218	41	219	42
rect	218	43	219	44
rect	218	44	219	45
rect	218	46	219	47
rect	218	47	219	48
rect	218	49	219	50
rect	218	50	219	51
rect	218	52	219	53
rect	218	53	219	54
rect	218	55	219	56
rect	218	56	219	57
rect	218	57	219	58
rect	218	59	219	60
rect	218	60	219	61
rect	218	62	219	63
rect	218	63	219	64
rect	218	65	219	66
rect	218	66	219	67
rect	218	68	219	69
rect	218	69	219	70
rect	218	71	219	72
rect	218	72	219	73
rect	218	74	219	75
rect	218	75	219	76
rect	218	77	219	78
rect	218	78	219	79
rect	218	80	219	81
rect	218	81	219	82
rect	218	82	219	83
rect	218	84	219	85
rect	218	85	219	86
rect	218	86	219	87
rect	218	87	219	88
rect	218	88	219	89
rect	218	90	219	91
rect	218	91	219	92
rect	218	93	219	94
rect	218	94	219	95
rect	218	96	219	97
rect	218	97	219	98
rect	218	98	219	99
rect	218	100	219	101
rect	218	101	219	102
rect	218	102	219	103
rect	218	103	219	104
rect	218	104	219	105
rect	218	106	219	107
rect	218	107	219	108
rect	218	109	219	110
rect	218	110	219	111
rect	218	111	219	112
rect	218	119	219	120
rect	218	120	219	121
rect	218	122	219	123
rect	218	123	219	124
rect	218	125	219	126
rect	218	126	219	127
rect	218	128	219	129
rect	218	138	219	139
rect	218	139	219	140
rect	218	141	219	142
rect	218	142	219	143
rect	218	144	219	145
rect	218	145	219	146
rect	218	147	219	148
rect	218	148	219	149
rect	218	149	219	150
rect	218	150	219	151
rect	218	151	219	152
rect	218	152	219	153
rect	218	154	219	155
rect	218	155	219	156
rect	218	157	219	158
rect	218	158	219	159
rect	218	160	219	161
rect	218	161	219	162
rect	218	163	219	164
rect	218	164	219	165
rect	218	165	219	166
rect	218	166	219	167
rect	218	181	219	182
rect	218	182	219	183
rect	218	183	219	184
rect	218	184	219	185
rect	218	185	219	186
rect	218	186	219	187
rect	233	34	234	35
rect	233	35	234	36
rect	233	36	234	37
rect	233	37	234	38
rect	233	38	234	39
rect	233	40	234	41
rect	233	41	234	42
rect	233	43	234	44
rect	233	44	234	45
rect	233	46	234	47
rect	233	47	234	48
rect	233	49	234	50
rect	233	50	234	51
rect	233	52	234	53
rect	233	53	234	54
rect	233	55	234	56
rect	233	56	234	57
rect	233	57	234	58
rect	233	59	234	60
rect	233	60	234	61
rect	233	62	234	63
rect	233	63	234	64
rect	233	65	234	66
rect	233	66	234	67
rect	233	68	234	69
rect	233	69	234	70
rect	233	71	234	72
rect	233	72	234	73
rect	233	74	234	75
rect	233	75	234	76
rect	233	77	234	78
rect	233	78	234	79
rect	233	80	234	81
rect	233	81	234	82
rect	233	82	234	83
rect	233	83	234	84
rect	233	84	234	85
rect	233	85	234	86
rect	233	87	234	88
rect	233	88	234	89
rect	233	90	234	91
rect	233	91	234	92
rect	233	93	234	94
rect	233	94	234	95
rect	233	96	234	97
rect	233	97	234	98
rect	233	98	234	99
rect	233	100	234	101
rect	233	101	234	102
rect	233	103	234	104
rect	233	104	234	105
rect	235	34	236	35
rect	235	35	236	36
rect	235	36	236	37
rect	235	37	236	38
rect	235	38	236	39
rect	235	40	236	41
rect	235	41	236	42
rect	237	43	238	44
rect	237	44	238	45
rect	237	46	238	47
rect	237	47	238	48
rect	237	49	238	50
rect	237	50	238	51
rect	237	52	238	53
rect	237	53	238	54
rect	237	55	238	56
rect	237	56	238	57
rect	237	57	238	58
rect	237	59	238	60
rect	237	60	238	61
rect	237	62	238	63
rect	237	63	238	64
rect	237	65	238	66
rect	237	66	238	67
rect	237	68	238	69
rect	237	69	238	70
rect	237	71	238	72
rect	237	72	238	73
rect	239	55	240	56
rect	239	56	240	57
rect	239	57	240	58
rect	239	74	240	75
rect	239	75	240	76
rect	239	77	240	78
rect	239	78	240	79
rect	239	80	240	81
rect	239	81	240	82
rect	239	82	240	83
rect	239	83	240	84
rect	239	84	240	85
rect	239	85	240	86
rect	241	21	242	22
rect	241	22	242	23
rect	241	24	242	25
rect	241	25	242	26
rect	241	27	242	28
rect	241	28	242	29
rect	241	30	242	31
rect	241	31	242	32
rect	241	32	242	33
rect	241	34	242	35
rect	241	35	242	36
rect	241	36	242	37
rect	241	37	242	38
rect	241	38	242	39
rect	241	40	242	41
rect	241	41	242	42
rect	241	43	242	44
rect	241	44	242	45
rect	241	46	242	47
rect	241	47	242	48
rect	241	49	242	50
rect	241	50	242	51
rect	241	52	242	53
rect	241	53	242	54
rect	241	54	242	55
rect	241	55	242	56
rect	241	56	242	57
rect	241	57	242	58
rect	241	58	242	59
rect	241	59	242	60
rect	241	60	242	61
rect	241	65	242	66
rect	241	66	242	67
rect	241	68	242	69
rect	241	69	242	70
rect	241	71	242	72
rect	241	72	242	73
rect	241	74	242	75
rect	241	75	242	76
rect	241	77	242	78
rect	241	78	242	79
rect	241	80	242	81
rect	241	81	242	82
rect	241	82	242	83
rect	243	21	244	22
rect	243	22	244	23
rect	243	24	244	25
rect	243	25	244	26
rect	243	27	244	28
rect	243	28	244	29
rect	243	30	244	31
rect	243	31	244	32
rect	243	32	244	33
rect	243	34	244	35
rect	243	35	244	36
rect	243	36	244	37
rect	243	37	244	38
rect	243	38	244	39
rect	243	40	244	41
rect	243	41	244	42
rect	243	43	244	44
rect	243	44	244	45
rect	243	46	244	47
rect	243	47	244	48
rect	243	49	244	50
rect	243	50	244	51
rect	243	55	244	56
rect	243	56	244	57
rect	243	57	244	58
rect	243	58	244	59
rect	243	59	244	60
rect	243	60	244	61
rect	243	61	244	62
rect	243	62	244	63
rect	243	63	244	64
rect	243	64	244	65
rect	243	65	244	66
rect	243	66	244	67
rect	243	68	244	69
rect	243	69	244	70
rect	243	71	244	72
rect	243	72	244	73
rect	243	74	244	75
rect	243	75	244	76
rect	243	77	244	78
rect	243	78	244	79
rect	243	80	244	81
rect	243	81	244	82
rect	243	82	244	83
rect	243	84	244	85
rect	243	85	244	86
rect	243	86	244	87
rect	243	87	244	88
rect	243	88	244	89
rect	243	90	244	91
rect	243	91	244	92
rect	243	93	244	94
rect	243	94	244	95
rect	243	96	244	97
rect	243	97	244	98
rect	243	98	244	99
rect	243	100	244	101
rect	243	101	244	102
rect	243	103	244	104
rect	243	104	244	105
rect	243	105	244	106
rect	243	106	244	107
rect	243	107	244	108
rect	243	109	244	110
rect	243	110	244	111
rect	243	111	244	112
rect	243	113	244	114
rect	243	114	244	115
rect	243	116	244	117
rect	243	117	244	118
rect	243	119	244	120
rect	243	120	244	121
rect	243	122	244	123
rect	243	123	244	124
rect	243	125	244	126
rect	243	126	244	127
rect	243	128	244	129
rect	243	129	244	130
rect	243	130	244	131
rect	243	132	244	133
rect	243	133	244	134
rect	245	52	246	53
rect	245	53	246	54
rect	245	55	246	56
rect	245	56	246	57
rect	245	57	246	58
rect	245	58	246	59
rect	245	59	246	60
rect	245	60	246	61
rect	245	61	246	62
rect	245	62	246	63
rect	245	63	246	64
rect	245	64	246	65
rect	245	65	246	66
rect	245	66	246	67
rect	245	68	246	69
rect	245	69	246	70
rect	245	71	246	72
rect	245	72	246	73
rect	245	74	246	75
rect	245	75	246	76
rect	247	40	248	41
rect	247	41	248	42
rect	247	43	248	44
rect	247	44	248	45
rect	247	46	248	47
rect	247	47	248	48
rect	247	49	248	50
rect	247	50	248	51
rect	247	52	248	53
rect	247	53	248	54
rect	247	55	248	56
rect	247	56	248	57
rect	247	57	248	58
rect	247	58	248	59
rect	247	59	248	60
rect	247	60	248	61
rect	247	61	248	62
rect	247	62	248	63
rect	247	63	248	64
rect	247	87	248	88
rect	247	88	248	89
rect	247	90	248	91
rect	247	91	248	92
rect	247	93	248	94
rect	247	94	248	95
rect	247	96	248	97
rect	247	97	248	98
rect	247	98	248	99
rect	247	100	248	101
rect	247	101	248	102
rect	247	130	248	131
rect	247	132	248	133
rect	247	133	248	134
rect	247	134	248	135
rect	247	135	248	136
rect	247	136	248	137
rect	247	138	248	139
rect	247	139	248	140
rect	247	141	248	142
rect	247	142	248	143
rect	247	144	248	145
rect	247	145	248	146
rect	247	147	248	148
rect	247	148	248	149
rect	247	149	248	150
rect	247	150	248	151
rect	247	151	248	152
rect	247	152	248	153
rect	247	153	248	154
rect	247	154	248	155
rect	247	155	248	156
rect	247	157	248	158
rect	247	158	248	159
rect	249	40	250	41
rect	249	41	250	42
rect	249	43	250	44
rect	249	44	250	45
rect	249	46	250	47
rect	249	47	250	48
rect	249	49	250	50
rect	249	50	250	51
rect	249	52	250	53
rect	249	53	250	54
rect	249	55	250	56
rect	249	56	250	57
rect	249	57	250	58
rect	249	58	250	59
rect	249	59	250	60
rect	249	60	250	61
rect	249	61	250	62
rect	249	62	250	63
rect	249	63	250	64
rect	249	65	250	66
rect	249	66	250	67
rect	249	68	250	69
rect	249	69	250	70
rect	249	77	250	78
rect	249	78	250	79
rect	249	80	250	81
rect	249	81	250	82
rect	249	82	250	83
rect	249	84	250	85
rect	249	85	250	86
rect	249	87	250	88
rect	249	88	250	89
rect	249	90	250	91
rect	249	91	250	92
rect	249	93	250	94
rect	249	94	250	95
rect	249	128	250	129
rect	249	130	250	131
rect	249	132	250	133
rect	251	8	252	9
rect	251	9	252	10
rect	251	10	252	11
rect	251	11	252	12
rect	251	12	252	13
rect	251	13	252	14
rect	251	15	252	16
rect	251	16	252	17
rect	251	37	252	38
rect	251	38	252	39
rect	251	40	252	41
rect	251	41	252	42
rect	251	43	252	44
rect	251	44	252	45
rect	251	46	252	47
rect	251	47	252	48
rect	251	49	252	50
rect	251	50	252	51
rect	251	52	252	53
rect	251	53	252	54
rect	251	55	252	56
rect	251	56	252	57
rect	251	57	252	58
rect	251	58	252	59
rect	251	59	252	60
rect	251	60	252	61
rect	251	61	252	62
rect	251	62	252	63
rect	251	63	252	64
rect	251	65	252	66
rect	251	66	252	67
rect	251	71	252	72
rect	251	72	252	73
rect	251	74	252	75
rect	251	75	252	76
rect	251	77	252	78
rect	251	78	252	79
rect	251	80	252	81
rect	251	81	252	82
rect	251	82	252	83
rect	251	84	252	85
rect	251	85	252	86
rect	251	87	252	88
rect	251	88	252	89
rect	251	90	252	91
rect	251	91	252	92
rect	251	107	252	108
rect	251	109	252	110
rect	251	110	252	111
rect	251	111	252	112
rect	251	113	252	114
rect	251	114	252	115
rect	251	116	252	117
rect	251	117	252	118
rect	251	127	252	128
rect	251	128	252	129
rect	251	130	252	131
rect	251	132	252	133
rect	251	134	252	135
rect	251	135	252	136
rect	251	136	252	137
rect	251	138	252	139
rect	251	139	252	140
rect	251	141	252	142
rect	251	142	252	143
rect	253	18	254	19
rect	253	19	254	20
rect	253	21	254	22
rect	253	22	254	23
rect	253	24	254	25
rect	253	25	254	26
rect	253	27	254	28
rect	253	28	254	29
rect	253	30	254	31
rect	253	31	254	32
rect	253	32	254	33
rect	253	34	254	35
rect	253	35	254	36
rect	253	37	254	38
rect	253	38	254	39
rect	253	40	254	41
rect	253	41	254	42
rect	253	43	254	44
rect	253	44	254	45
rect	253	46	254	47
rect	253	47	254	48
rect	253	49	254	50
rect	253	50	254	51
rect	253	52	254	53
rect	253	53	254	54
rect	253	55	254	56
rect	253	56	254	57
rect	253	57	254	58
rect	253	58	254	59
rect	253	59	254	60
rect	253	60	254	61
rect	253	61	254	62
rect	253	62	254	63
rect	253	63	254	64
rect	253	65	254	66
rect	253	66	254	67
rect	253	67	254	68
rect	253	68	254	69
rect	253	69	254	70
rect	253	71	254	72
rect	253	72	254	73
rect	253	74	254	75
rect	253	75	254	76
rect	253	77	254	78
rect	253	78	254	79
rect	253	80	254	81
rect	253	81	254	82
rect	253	82	254	83
rect	253	84	254	85
rect	253	85	254	86
rect	253	87	254	88
rect	253	88	254	89
rect	253	90	254	91
rect	253	91	254	92
rect	253	92	254	93
rect	253	93	254	94
rect	253	94	254	95
rect	253	95	254	96
rect	253	96	254	97
rect	253	97	254	98
rect	253	98	254	99
rect	253	103	254	104
rect	253	104	254	105
rect	253	105	254	106
rect	253	107	254	108
rect	253	109	254	110
rect	253	110	254	111
rect	253	111	254	112
rect	253	113	254	114
rect	253	114	254	115
rect	253	116	254	117
rect	253	117	254	118
rect	253	118	254	119
rect	253	119	254	120
rect	253	120	254	121
rect	253	122	254	123
rect	253	123	254	124
rect	253	125	254	126
rect	253	127	254	128
rect	253	128	254	129
rect	253	130	254	131
rect	253	132	254	133
rect	253	134	254	135
rect	253	135	254	136
rect	253	136	254	137
rect	253	138	254	139
rect	253	139	254	140
rect	255	68	256	69
rect	255	69	256	70
rect	255	71	256	72
rect	255	72	256	73
rect	255	74	256	75
rect	255	75	256	76
rect	255	77	256	78
rect	255	78	256	79
rect	255	80	256	81
rect	255	81	256	82
rect	255	82	256	83
rect	255	84	256	85
rect	255	85	256	86
rect	255	87	256	88
rect	255	88	256	89
rect	255	100	256	101
rect	255	101	256	102
rect	255	103	256	104
rect	255	104	256	105
rect	255	105	256	106
rect	255	107	256	108
rect	255	109	256	110
rect	255	110	256	111
rect	255	111	256	112
rect	255	113	256	114
rect	255	114	256	115
rect	255	116	256	117
rect	255	117	256	118
rect	255	118	256	119
rect	255	119	256	120
rect	255	120	256	121
rect	255	122	256	123
rect	255	123	256	124
rect	255	125	256	126
rect	255	127	256	128
rect	255	128	256	129
rect	255	130	256	131
rect	255	132	256	133
rect	255	134	256	135
rect	255	135	256	136
rect	255	136	256	137
rect	257	5	258	6
rect	257	6	258	7
rect	257	8	258	9
rect	257	9	258	10
rect	257	10	258	11
rect	257	11	258	12
rect	257	12	258	13
rect	257	13	258	14
rect	257	15	258	16
rect	257	16	258	17
rect	257	18	258	19
rect	257	19	258	20
rect	257	21	258	22
rect	257	22	258	23
rect	257	24	258	25
rect	257	25	258	26
rect	257	27	258	28
rect	257	28	258	29
rect	257	58	258	59
rect	257	59	258	60
rect	257	60	258	61
rect	257	61	258	62
rect	257	62	258	63
rect	257	63	258	64
rect	257	65	258	66
rect	257	66	258	67
rect	257	68	258	69
rect	257	69	258	70
rect	257	71	258	72
rect	257	72	258	73
rect	257	74	258	75
rect	257	75	258	76
rect	257	77	258	78
rect	257	78	258	79
rect	257	80	258	81
rect	257	81	258	82
rect	257	82	258	83
rect	257	84	258	85
rect	257	85	258	86
rect	257	87	258	88
rect	257	88	258	89
rect	257	89	258	90
rect	257	90	258	91
rect	257	91	258	92
rect	257	92	258	93
rect	257	93	258	94
rect	257	94	258	95
rect	257	95	258	96
rect	257	96	258	97
rect	257	97	258	98
rect	257	98	258	99
rect	257	100	258	101
rect	257	101	258	102
rect	257	103	258	104
rect	257	104	258	105
rect	257	105	258	106
rect	257	107	258	108
rect	257	109	258	110
rect	257	110	258	111
rect	257	111	258	112
rect	257	116	258	117
rect	257	117	258	118
rect	257	118	258	119
rect	257	119	258	120
rect	257	120	258	121
rect	257	125	258	126
rect	257	127	258	128
rect	257	128	258	129
rect	257	130	258	131
rect	257	140	258	141
rect	257	141	258	142
rect	257	142	258	143
rect	257	143	258	144
rect	257	144	258	145
rect	257	145	258	146
rect	257	157	258	158
rect	257	158	258	159
rect	257	159	258	160
rect	257	160	258	161
rect	257	161	258	162
rect	257	163	258	164
rect	257	164	258	165
rect	257	165	258	166
rect	259	15	260	16
rect	259	16	260	17
rect	259	18	260	19
rect	259	19	260	20
rect	259	21	260	22
rect	259	22	260	23
rect	259	24	260	25
rect	259	25	260	26
rect	259	27	260	28
rect	259	28	260	29
rect	259	29	260	30
rect	259	61	260	62
rect	259	62	260	63
rect	259	63	260	64
rect	259	65	260	66
rect	259	66	260	67
rect	259	68	260	69
rect	259	69	260	70
rect	259	71	260	72
rect	259	72	260	73
rect	259	74	260	75
rect	259	75	260	76
rect	259	77	260	78
rect	259	78	260	79
rect	259	90	260	91
rect	259	91	260	92
rect	259	92	260	93
rect	259	93	260	94
rect	259	94	260	95
rect	259	95	260	96
rect	259	96	260	97
rect	259	97	260	98
rect	259	98	260	99
rect	259	100	260	101
rect	259	101	260	102
rect	259	103	260	104
rect	259	104	260	105
rect	259	105	260	106
rect	259	107	260	108
rect	259	113	260	114
rect	259	114	260	115
rect	259	115	260	116
rect	259	116	260	117
rect	259	117	260	118
rect	259	118	260	119
rect	259	119	260	120
rect	259	120	260	121
rect	259	121	260	122
rect	259	122	260	123
rect	259	123	260	124
rect	259	124	260	125
rect	259	125	260	126
rect	259	127	260	128
rect	259	128	260	129
rect	259	130	260	131
rect	259	131	260	132
rect	259	132	260	133
rect	259	134	260	135
rect	259	135	260	136
rect	259	136	260	137
rect	259	137	260	138
rect	259	138	260	139
rect	259	140	260	141
rect	259	141	260	142
rect	259	142	260	143
rect	259	143	260	144
rect	259	144	260	145
rect	259	145	260	146
rect	259	146	260	147
rect	259	147	260	148
rect	259	148	260	149
rect	259	149	260	150
rect	259	150	260	151
rect	259	151	260	152
rect	259	152	260	153
rect	259	153	260	154
rect	259	154	260	155
rect	259	155	260	156
rect	259	156	260	157
rect	259	157	260	158
rect	259	158	260	159
rect	259	159	260	160
rect	259	160	260	161
rect	259	161	260	162
rect	268	29	269	30
rect	268	31	269	32
rect	268	32	269	33
rect	268	34	269	35
rect	268	35	269	36
rect	268	37	269	38
rect	268	38	269	39
rect	268	40	269	41
rect	268	41	269	42
rect	268	43	269	44
rect	268	44	269	45
rect	268	46	269	47
rect	268	47	269	48
rect	268	49	269	50
rect	268	50	269	51
rect	268	52	269	53
rect	268	53	269	54
rect	270	34	271	35
rect	270	35	271	36
rect	270	37	271	38
rect	270	38	271	39
rect	270	40	271	41
rect	270	41	271	42
rect	270	43	271	44
rect	270	44	271	45
rect	270	46	271	47
rect	270	47	271	48
rect	270	49	271	50
rect	270	50	271	51
rect	270	56	271	57
rect	270	58	271	59
rect	270	59	271	60
rect	272	53	273	54
rect	272	54	273	55
rect	272	56	273	57
rect	272	58	273	59
rect	272	59	273	60
rect	272	60	273	61
rect	272	61	273	62
rect	272	62	273	63
rect	272	63	273	64
rect	272	65	273	66
rect	272	66	273	67
rect	272	68	273	69
rect	272	69	273	70
rect	272	71	273	72
rect	272	72	273	73
rect	272	74	273	75
rect	272	75	273	76
rect	274	49	275	50
rect	274	50	275	51
rect	274	51	275	52
rect	274	53	275	54
rect	274	54	275	55
rect	274	56	275	57
rect	274	58	275	59
rect	274	59	275	60
rect	274	60	275	61
rect	274	61	275	62
rect	274	62	275	63
rect	274	63	275	64
rect	274	81	275	82
rect	274	82	275	83
rect	274	84	275	85
rect	274	85	275	86
rect	276	12	277	13
rect	276	13	277	14
rect	276	14	277	15
rect	276	15	277	16
rect	276	16	277	17
rect	276	18	277	19
rect	276	19	277	20
rect	276	50	277	51
rect	276	51	277	52
rect	276	53	277	54
rect	276	54	277	55
rect	276	56	277	57
rect	276	58	277	59
rect	276	59	277	60
rect	276	60	277	61
rect	276	61	277	62
rect	276	62	277	63
rect	276	63	277	64
rect	276	64	277	65
rect	276	65	277	66
rect	276	66	277	67
rect	276	68	277	69
rect	276	69	277	70
rect	276	71	277	72
rect	276	72	277	73
rect	276	74	277	75
rect	276	75	277	76
rect	276	76	277	77
rect	276	77	277	78
rect	276	78	277	79
rect	276	79	277	80
rect	276	80	277	81
rect	276	81	277	82
rect	276	82	277	83
rect	276	84	277	85
rect	276	85	277	86
rect	276	86	277	87
rect	276	87	277	88
rect	276	88	277	89
rect	276	90	277	91
rect	276	91	277	92
rect	276	92	277	93
rect	276	93	277	94
rect	276	94	277	95
rect	276	95	277	96
rect	276	96	277	97
rect	276	97	277	98
rect	276	98	277	99
rect	278	12	279	13
rect	278	13	279	14
rect	278	14	279	15
rect	278	15	279	16
rect	278	16	279	17
rect	278	22	279	23
rect	278	24	279	25
rect	278	26	279	27
rect	278	27	279	28
rect	278	29	279	30
rect	278	31	279	32
rect	278	32	279	33
rect	278	33	279	34
rect	278	34	279	35
rect	278	35	279	36
rect	278	37	279	38
rect	278	38	279	39
rect	278	46	279	47
rect	278	47	279	48
rect	278	48	279	49
rect	278	50	279	51
rect	278	51	279	52
rect	278	53	279	54
rect	278	54	279	55
rect	278	56	279	57
rect	278	58	279	59
rect	278	59	279	60
rect	278	60	279	61
rect	278	61	279	62
rect	278	62	279	63
rect	278	63	279	64
rect	278	64	279	65
rect	278	65	279	66
rect	278	66	279	67
rect	278	74	279	75
rect	278	75	279	76
rect	278	76	279	77
rect	278	77	279	78
rect	278	78	279	79
rect	278	79	279	80
rect	278	80	279	81
rect	278	81	279	82
rect	278	82	279	83
rect	280	19	281	20
rect	280	20	281	21
rect	280	22	281	23
rect	280	24	281	25
rect	280	26	281	27
rect	280	27	281	28
rect	280	29	281	30
rect	280	31	281	32
rect	280	32	281	33
rect	280	33	281	34
rect	280	34	281	35
rect	280	35	281	36
rect	280	40	281	41
rect	280	41	281	42
rect	280	43	281	44
rect	280	44	281	45
rect	280	45	281	46
rect	280	46	281	47
rect	280	47	281	48
rect	280	48	281	49
rect	280	50	281	51
rect	280	51	281	52
rect	280	53	281	54
rect	280	54	281	55
rect	280	56	281	57
rect	280	58	281	59
rect	280	59	281	60
rect	280	60	281	61
rect	280	61	281	62
rect	280	62	281	63
rect	280	63	281	64
rect	280	64	281	65
rect	280	65	281	66
rect	280	66	281	67
rect	280	67	281	68
rect	280	68	281	69
rect	280	69	281	70
rect	280	74	281	75
rect	280	75	281	76
rect	280	76	281	77
rect	280	77	281	78
rect	280	78	281	79
rect	280	79	281	80
rect	280	80	281	81
rect	280	81	281	82
rect	280	82	281	83
rect	280	83	281	84
rect	280	84	281	85
rect	280	85	281	86
rect	280	86	281	87
rect	280	87	281	88
rect	280	88	281	89
rect	280	90	281	91
rect	280	91	281	92
rect	280	92	281	93
rect	280	93	281	94
rect	280	94	281	95
rect	280	95	281	96
rect	280	96	281	97
rect	280	97	281	98
rect	280	98	281	99
rect	280	99	281	100
rect	280	100	281	101
rect	280	101	281	102
rect	280	117	281	118
rect	280	118	281	119
rect	280	120	281	121
rect	280	121	281	122
rect	280	122	281	123
rect	280	123	281	124
rect	280	124	281	125
rect	280	125	281	126
rect	280	127	281	128
rect	280	128	281	129
rect	282	5	283	6
rect	282	6	283	7
rect	282	15	283	16
rect	282	16	283	17
rect	282	17	283	18
rect	282	19	283	20
rect	282	20	283	21
rect	282	22	283	23
rect	282	31	283	32
rect	282	32	283	33
rect	282	33	283	34
rect	282	34	283	35
rect	282	35	283	36
rect	282	36	283	37
rect	282	37	283	38
rect	282	38	283	39
rect	282	40	283	41
rect	282	41	283	42
rect	282	46	283	47
rect	282	47	283	48
rect	282	48	283	49
rect	282	50	283	51
rect	282	51	283	52
rect	282	53	283	54
rect	282	54	283	55
rect	282	56	283	57
rect	282	63	283	64
rect	282	64	283	65
rect	282	65	283	66
rect	282	66	283	67
rect	282	67	283	68
rect	282	68	283	69
rect	282	69	283	70
rect	282	70	283	71
rect	282	71	283	72
rect	282	72	283	73
rect	282	74	283	75
rect	282	75	283	76
rect	282	76	283	77
rect	282	77	283	78
rect	282	78	283	79
rect	282	79	283	80
rect	282	80	283	81
rect	282	81	283	82
rect	282	82	283	83
rect	282	83	283	84
rect	282	84	283	85
rect	282	85	283	86
rect	282	86	283	87
rect	282	87	283	88
rect	282	88	283	89
rect	282	113	283	114
rect	282	114	283	115
rect	282	115	283	116
rect	282	116	283	117
rect	282	117	283	118
rect	282	118	283	119
rect	282	127	283	128
rect	282	128	283	129
rect	282	129	283	130
rect	282	130	283	131
rect	282	131	283	132
rect	282	132	283	133
rect	282	133	283	134
rect	282	134	283	135
rect	282	135	283	136
rect	282	136	283	137
rect	282	137	283	138
rect	282	138	283	139
rect	291	12	292	13
rect	291	13	292	14
rect	291	40	292	41
rect	291	41	292	42
rect	291	42	292	43
rect	291	43	292	44
rect	291	44	292	45
rect	291	56	292	57
rect	291	57	292	58
rect	291	58	292	59
rect	293	9	294	10
rect	293	10	294	11
rect	293	11	294	12
rect	293	12	294	13
rect	293	13	294	14
rect	293	14	294	15
rect	293	15	294	16
rect	293	16	294	17
rect	293	17	294	18
rect	293	18	294	19
rect	293	19	294	20
rect	293	20	294	21
rect	293	21	294	22
rect	293	22	294	23
rect	293	23	294	24
rect	293	24	294	25
rect	293	25	294	26
rect	293	26	294	27
rect	293	27	294	28
rect	293	28	294	29
rect	293	29	294	30
rect	293	30	294	31
rect	293	31	294	32
rect	293	32	294	33
rect	293	33	294	34
rect	293	34	294	35
rect	293	35	294	36
rect	293	36	294	37
rect	293	37	294	38
rect	293	38	294	39
rect	293	39	294	40
rect	293	40	294	41
rect	293	41	294	42
rect	293	42	294	43
rect	293	43	294	44
rect	293	44	294	45
rect	293	45	294	46
rect	293	46	294	47
rect	293	47	294	48
rect	293	48	294	49
rect	293	49	294	50
rect	293	50	294	51
rect	293	51	294	52
rect	293	52	294	53
rect	293	53	294	54
rect	293	54	294	55
rect	293	55	294	56
rect	293	56	294	57
rect	293	57	294	58
rect	293	58	294	59
rect	293	59	294	60
rect	293	60	294	61
rect	293	61	294	62
rect	293	62	294	63
rect	293	63	294	64
rect	293	64	294	65
rect	293	65	294	66
rect	293	66	294	67
rect	293	67	294	68
rect	293	68	294	69
rect	293	69	294	70
rect	293	70	294	71
rect	293	71	294	72
rect	293	72	294	73
<< metal2 >>
rect	1	40	2	41
rect	1	46	2	47
rect	2	40	3	41
rect	2	46	3	47
rect	3	37	4	38
rect	3	40	4	41
rect	3	43	4	44
rect	3	46	4	47
rect	3	63	4	64
rect	3	73	4	74
rect	3	83	4	84
rect	3	87	4	88
rect	3	90	4	91
rect	3	93	4	94
rect	4	37	5	38
rect	4	40	5	41
rect	4	43	5	44
rect	4	46	5	47
rect	4	63	5	64
rect	4	73	5	74
rect	4	83	5	84
rect	4	87	5	88
rect	4	90	5	91
rect	4	93	5	94
rect	5	4	6	5
rect	5	10	6	11
rect	5	33	6	34
rect	5	37	6	38
rect	5	40	6	41
rect	5	43	6	44
rect	5	46	6	47
rect	5	50	6	51
rect	5	60	6	61
rect	5	63	6	64
rect	5	66	6	67
rect	5	73	6	74
rect	5	77	6	78
rect	5	83	6	84
rect	5	87	6	88
rect	5	90	6	91
rect	5	93	6	94
rect	5	103	6	104
rect	6	4	7	5
rect	6	10	7	11
rect	6	33	7	34
rect	6	37	7	38
rect	6	40	7	41
rect	6	43	7	44
rect	6	46	7	47
rect	6	50	7	51
rect	6	60	7	61
rect	6	63	7	64
rect	6	66	7	67
rect	6	73	7	74
rect	6	77	7	78
rect	6	83	7	84
rect	6	87	7	88
rect	6	90	7	91
rect	6	93	7	94
rect	6	103	7	104
rect	7	1	8	2
rect	7	4	8	5
rect	7	7	8	8
rect	7	10	8	11
rect	7	17	8	18
rect	7	20	8	21
rect	7	23	8	24
rect	7	33	8	34
rect	7	37	8	38
rect	7	40	8	41
rect	7	43	8	44
rect	7	46	8	47
rect	7	50	8	51
rect	7	60	8	61
rect	7	63	8	64
rect	7	66	8	67
rect	7	73	8	74
rect	7	77	8	78
rect	7	83	8	84
rect	7	87	8	88
rect	7	90	8	91
rect	7	93	8	94
rect	7	97	8	98
rect	7	103	8	104
rect	9	16	10	17
rect	9	17	10	18
rect	9	19	10	20
rect	9	20	10	21
rect	9	22	10	23
rect	9	23	10	24
rect	9	25	10	26
rect	9	26	10	27
rect	9	34	10	35
rect	9	35	10	36
rect	9	53	10	54
rect	9	54	10	55
rect	9	58	10	59
rect	9	59	10	60
rect	9	72	10	73
rect	9	73	10	74
rect	9	74	10	75
rect	9	75	10	76
rect	9	80	10	81
rect	9	81	10	82
rect	9	83	10	84
rect	9	84	10	85
rect	10	16	11	17
rect	10	17	11	18
rect	10	19	11	20
rect	10	20	11	21
rect	10	22	11	23
rect	10	23	11	24
rect	10	25	11	26
rect	10	26	11	27
rect	10	34	11	35
rect	10	35	11	36
rect	10	53	11	54
rect	10	54	11	55
rect	10	58	11	59
rect	10	59	11	60
rect	10	72	11	73
rect	10	73	11	74
rect	10	74	11	75
rect	10	75	11	76
rect	10	80	11	81
rect	10	81	11	82
rect	10	83	11	84
rect	10	84	11	85
rect	11	16	12	17
rect	11	17	12	18
rect	11	19	12	20
rect	11	20	12	21
rect	11	22	12	23
rect	11	23	12	24
rect	11	25	12	26
rect	11	26	12	27
rect	11	34	12	35
rect	11	35	12	36
rect	11	53	12	54
rect	11	54	12	55
rect	11	58	12	59
rect	11	59	12	60
rect	11	72	12	73
rect	11	73	12	74
rect	11	74	12	75
rect	11	75	12	76
rect	11	80	12	81
rect	11	81	12	82
rect	11	83	12	84
rect	11	84	12	85
rect	12	16	13	17
rect	12	17	13	18
rect	12	19	13	20
rect	12	20	13	21
rect	12	22	13	23
rect	12	23	13	24
rect	12	25	13	26
rect	12	26	13	27
rect	12	34	13	35
rect	12	35	13	36
rect	12	53	13	54
rect	12	54	13	55
rect	12	58	13	59
rect	12	59	13	60
rect	12	72	13	73
rect	12	73	13	74
rect	12	74	13	75
rect	12	75	13	76
rect	12	80	13	81
rect	12	81	13	82
rect	12	83	13	84
rect	12	84	13	85
rect	13	16	14	17
rect	13	17	14	18
rect	13	19	14	20
rect	13	20	14	21
rect	13	22	14	23
rect	13	23	14	24
rect	13	25	14	26
rect	13	26	14	27
rect	13	34	14	35
rect	13	35	14	36
rect	13	53	14	54
rect	13	54	14	55
rect	13	58	14	59
rect	13	59	14	60
rect	13	72	14	73
rect	13	73	14	74
rect	13	74	14	75
rect	13	75	14	76
rect	13	80	14	81
rect	13	81	14	82
rect	13	83	14	84
rect	13	84	14	85
rect	14	1	15	2
rect	14	4	15	5
rect	14	10	15	11
rect	14	14	15	15
rect	14	16	15	17
rect	14	17	15	18
rect	14	19	15	20
rect	14	20	15	21
rect	14	22	15	23
rect	14	23	15	24
rect	14	25	15	26
rect	14	26	15	27
rect	14	27	15	28
rect	14	33	15	34
rect	14	34	15	35
rect	14	35	15	36
rect	14	37	15	38
rect	14	43	15	44
rect	14	46	15	47
rect	14	50	15	51
rect	14	53	15	54
rect	14	54	15	55
rect	14	58	15	59
rect	14	59	15	60
rect	14	63	15	64
rect	14	66	15	67
rect	14	72	15	73
rect	14	73	15	74
rect	14	74	15	75
rect	14	75	15	76
rect	14	77	15	78
rect	14	80	15	81
rect	14	81	15	82
rect	14	83	15	84
rect	14	84	15	85
rect	14	87	15	88
rect	14	93	15	94
rect	14	100	15	101
rect	14	103	15	104
rect	15	1	16	2
rect	15	4	16	5
rect	15	10	16	11
rect	15	14	16	15
rect	15	16	16	17
rect	15	17	16	18
rect	15	19	16	20
rect	15	20	16	21
rect	15	22	16	23
rect	15	23	16	24
rect	15	25	16	26
rect	15	26	16	27
rect	15	27	16	28
rect	15	33	16	34
rect	15	34	16	35
rect	15	35	16	36
rect	15	37	16	38
rect	15	43	16	44
rect	15	46	16	47
rect	15	53	16	54
rect	15	54	16	55
rect	15	58	16	59
rect	15	59	16	60
rect	15	63	16	64
rect	15	66	16	67
rect	15	72	16	73
rect	15	73	16	74
rect	15	74	16	75
rect	15	75	16	76
rect	15	77	16	78
rect	15	80	16	81
rect	15	81	16	82
rect	15	83	16	84
rect	15	84	16	85
rect	15	87	16	88
rect	15	93	16	94
rect	15	100	16	101
rect	15	103	16	104
rect	16	1	17	2
rect	16	4	17	5
rect	16	10	17	11
rect	16	14	17	15
rect	16	16	17	17
rect	16	17	17	18
rect	16	19	17	20
rect	16	20	17	21
rect	16	22	17	23
rect	16	23	17	24
rect	16	25	17	26
rect	16	26	17	27
rect	16	27	17	28
rect	16	33	17	34
rect	16	34	17	35
rect	16	35	17	36
rect	16	37	17	38
rect	16	43	17	44
rect	16	46	17	47
rect	16	53	17	54
rect	16	54	17	55
rect	16	58	17	59
rect	16	59	17	60
rect	16	63	17	64
rect	16	66	17	67
rect	16	71	17	72
rect	16	72	17	73
rect	16	73	17	74
rect	16	74	17	75
rect	16	75	17	76
rect	16	77	17	78
rect	16	80	17	81
rect	16	81	17	82
rect	16	83	17	84
rect	16	84	17	85
rect	16	87	17	88
rect	16	93	17	94
rect	16	100	17	101
rect	16	103	17	104
rect	17	1	18	2
rect	17	4	18	5
rect	17	10	18	11
rect	17	14	18	15
rect	17	16	18	17
rect	17	17	18	18
rect	17	19	18	20
rect	17	20	18	21
rect	17	22	18	23
rect	17	23	18	24
rect	17	25	18	26
rect	17	26	18	27
rect	17	27	18	28
rect	17	33	18	34
rect	17	34	18	35
rect	17	35	18	36
rect	17	37	18	38
rect	17	46	18	47
rect	17	53	18	54
rect	17	54	18	55
rect	17	58	18	59
rect	17	59	18	60
rect	17	63	18	64
rect	17	66	18	67
rect	17	71	18	72
rect	17	72	18	73
rect	17	73	18	74
rect	17	74	18	75
rect	17	75	18	76
rect	17	80	18	81
rect	17	81	18	82
rect	17	83	18	84
rect	17	84	18	85
rect	17	87	18	88
rect	17	93	18	94
rect	17	100	18	101
rect	17	103	18	104
rect	18	1	19	2
rect	18	4	19	5
rect	18	10	19	11
rect	18	14	19	15
rect	18	16	19	17
rect	18	17	19	18
rect	18	19	19	20
rect	18	20	19	21
rect	18	22	19	23
rect	18	23	19	24
rect	18	25	19	26
rect	18	26	19	27
rect	18	27	19	28
rect	18	33	19	34
rect	18	34	19	35
rect	18	35	19	36
rect	18	37	19	38
rect	18	46	19	47
rect	18	53	19	54
rect	18	54	19	55
rect	18	55	19	56
rect	18	58	19	59
rect	18	59	19	60
rect	18	63	19	64
rect	18	66	19	67
rect	18	71	19	72
rect	18	72	19	73
rect	18	73	19	74
rect	18	74	19	75
rect	18	75	19	76
rect	18	80	19	81
rect	18	81	19	82
rect	18	83	19	84
rect	18	84	19	85
rect	18	87	19	88
rect	18	93	19	94
rect	18	100	19	101
rect	18	103	19	104
rect	18	115	19	116
rect	19	1	20	2
rect	19	4	20	5
rect	19	10	20	11
rect	19	14	20	15
rect	19	16	20	17
rect	19	19	20	20
rect	19	20	20	21
rect	19	22	20	23
rect	19	23	20	24
rect	19	25	20	26
rect	19	26	20	27
rect	19	27	20	28
rect	19	33	20	34
rect	19	34	20	35
rect	19	35	20	36
rect	19	37	20	38
rect	19	46	20	47
rect	19	53	20	54
rect	19	54	20	55
rect	19	55	20	56
rect	19	58	20	59
rect	19	59	20	60
rect	19	63	20	64
rect	19	66	20	67
rect	19	71	20	72
rect	19	72	20	73
rect	19	73	20	74
rect	19	74	20	75
rect	19	75	20	76
rect	19	80	20	81
rect	19	81	20	82
rect	19	83	20	84
rect	19	84	20	85
rect	19	87	20	88
rect	19	100	20	101
rect	19	103	20	104
rect	19	115	20	116
rect	20	1	21	2
rect	20	4	21	5
rect	20	7	21	8
rect	20	10	21	11
rect	20	14	21	15
rect	20	16	21	17
rect	20	17	21	18
rect	20	19	21	20
rect	20	20	21	21
rect	20	22	21	23
rect	20	23	21	24
rect	20	25	21	26
rect	20	26	21	27
rect	20	27	21	28
rect	20	33	21	34
rect	20	34	21	35
rect	20	35	21	36
rect	20	37	21	38
rect	20	39	21	40
rect	20	46	21	47
rect	20	53	21	54
rect	20	54	21	55
rect	20	55	21	56
rect	20	58	21	59
rect	20	59	21	60
rect	20	63	21	64
rect	20	66	21	67
rect	20	71	21	72
rect	20	72	21	73
rect	20	73	21	74
rect	20	74	21	75
rect	20	75	21	76
rect	20	77	21	78
rect	20	80	21	81
rect	20	81	21	82
rect	20	83	21	84
rect	20	84	21	85
rect	20	87	21	88
rect	20	100	21	101
rect	20	103	21	104
rect	20	112	21	113
rect	20	115	21	116
rect	21	1	22	2
rect	21	4	22	5
rect	21	7	22	8
rect	21	10	22	11
rect	21	14	22	15
rect	21	16	22	17
rect	21	17	22	18
rect	21	19	22	20
rect	21	20	22	21
rect	21	22	22	23
rect	21	23	22	24
rect	21	25	22	26
rect	21	26	22	27
rect	21	27	22	28
rect	21	34	22	35
rect	21	35	22	36
rect	21	39	22	40
rect	21	46	22	47
rect	21	53	22	54
rect	21	54	22	55
rect	21	55	22	56
rect	21	58	22	59
rect	21	59	22	60
rect	21	63	22	64
rect	21	66	22	67
rect	21	71	22	72
rect	21	72	22	73
rect	21	73	22	74
rect	21	74	22	75
rect	21	75	22	76
rect	21	77	22	78
rect	21	80	22	81
rect	21	81	22	82
rect	21	83	22	84
rect	21	84	22	85
rect	21	87	22	88
rect	21	100	22	101
rect	21	103	22	104
rect	21	112	22	113
rect	21	115	22	116
rect	22	1	23	2
rect	22	4	23	5
rect	22	7	23	8
rect	22	10	23	11
rect	22	14	23	15
rect	22	16	23	17
rect	22	17	23	18
rect	22	19	23	20
rect	22	20	23	21
rect	22	22	23	23
rect	22	23	23	24
rect	22	25	23	26
rect	22	26	23	27
rect	22	27	23	28
rect	22	29	23	30
rect	22	34	23	35
rect	22	35	23	36
rect	22	39	23	40
rect	22	46	23	47
rect	22	52	23	53
rect	22	53	23	54
rect	22	54	23	55
rect	22	55	23	56
rect	22	58	23	59
rect	22	59	23	60
rect	22	63	23	64
rect	22	66	23	67
rect	22	71	23	72
rect	22	72	23	73
rect	22	73	23	74
rect	22	74	23	75
rect	22	75	23	76
rect	22	77	23	78
rect	22	80	23	81
rect	22	81	23	82
rect	22	83	23	84
rect	22	84	23	85
rect	22	87	23	88
rect	22	93	23	94
rect	22	100	23	101
rect	22	103	23	104
rect	22	112	23	113
rect	22	115	23	116
rect	22	139	23	140
rect	23	1	24	2
rect	23	4	24	5
rect	23	7	24	8
rect	23	16	24	17
rect	23	17	24	18
rect	23	19	24	20
rect	23	20	24	21
rect	23	22	24	23
rect	23	23	24	24
rect	23	25	24	26
rect	23	26	24	27
rect	23	29	24	30
rect	23	34	24	35
rect	23	35	24	36
rect	23	39	24	40
rect	23	52	24	53
rect	23	53	24	54
rect	23	54	24	55
rect	23	55	24	56
rect	23	59	24	60
rect	23	66	24	67
rect	23	71	24	72
rect	23	72	24	73
rect	23	73	24	74
rect	23	74	24	75
rect	23	75	24	76
rect	23	77	24	78
rect	23	80	24	81
rect	23	81	24	82
rect	23	83	24	84
rect	23	84	24	85
rect	23	87	24	88
rect	23	93	24	94
rect	23	112	24	113
rect	23	115	24	116
rect	23	139	24	140
rect	24	1	25	2
rect	24	4	25	5
rect	24	7	25	8
rect	24	16	25	17
rect	24	17	25	18
rect	24	19	25	20
rect	24	20	25	21
rect	24	22	25	23
rect	24	23	25	24
rect	24	25	25	26
rect	24	26	25	27
rect	24	29	25	30
rect	24	34	25	35
rect	24	35	25	36
rect	24	39	25	40
rect	24	42	25	43
rect	24	52	25	53
rect	24	53	25	54
rect	24	54	25	55
rect	24	55	25	56
rect	24	58	25	59
rect	24	59	25	60
rect	24	61	25	62
rect	24	66	25	67
rect	24	68	25	69
rect	24	71	25	72
rect	24	72	25	73
rect	24	73	25	74
rect	24	74	25	75
rect	24	75	25	76
rect	24	77	25	78
rect	24	80	25	81
rect	24	81	25	82
rect	24	83	25	84
rect	24	84	25	85
rect	24	87	25	88
rect	24	93	25	94
rect	24	96	25	97
rect	24	99	25	100
rect	24	112	25	113
rect	24	115	25	116
rect	24	139	25	140
rect	24	142	25	143
rect	25	1	26	2
rect	25	4	26	5
rect	25	7	26	8
rect	25	16	26	17
rect	25	17	26	18
rect	25	19	26	20
rect	25	20	26	21
rect	25	22	26	23
rect	25	23	26	24
rect	25	25	26	26
rect	25	26	26	27
rect	25	29	26	30
rect	25	34	26	35
rect	25	35	26	36
rect	25	39	26	40
rect	25	42	26	43
rect	25	52	26	53
rect	25	53	26	54
rect	25	54	26	55
rect	25	55	26	56
rect	25	58	26	59
rect	25	59	26	60
rect	25	61	26	62
rect	25	66	26	67
rect	25	68	26	69
rect	25	71	26	72
rect	25	72	26	73
rect	25	73	26	74
rect	25	74	26	75
rect	25	75	26	76
rect	25	77	26	78
rect	25	80	26	81
rect	25	81	26	82
rect	25	83	26	84
rect	25	84	26	85
rect	25	87	26	88
rect	25	93	26	94
rect	25	96	26	97
rect	25	99	26	100
rect	25	112	26	113
rect	25	115	26	116
rect	25	139	26	140
rect	25	142	26	143
rect	26	1	27	2
rect	26	4	27	5
rect	26	7	27	8
rect	26	14	27	15
rect	26	16	27	17
rect	26	17	27	18
rect	26	19	27	20
rect	26	20	27	21
rect	26	22	27	23
rect	26	23	27	24
rect	26	25	27	26
rect	26	26	27	27
rect	26	29	27	30
rect	26	34	27	35
rect	26	35	27	36
rect	26	39	27	40
rect	26	42	27	43
rect	26	52	27	53
rect	26	53	27	54
rect	26	54	27	55
rect	26	55	27	56
rect	26	58	27	59
rect	26	59	27	60
rect	26	61	27	62
rect	26	66	27	67
rect	26	68	27	69
rect	26	71	27	72
rect	26	72	27	73
rect	26	73	27	74
rect	26	74	27	75
rect	26	75	27	76
rect	26	77	27	78
rect	26	80	27	81
rect	26	81	27	82
rect	26	83	27	84
rect	26	84	27	85
rect	26	87	27	88
rect	26	93	27	94
rect	26	96	27	97
rect	26	99	27	100
rect	26	102	27	103
rect	26	112	27	113
rect	26	115	27	116
rect	26	139	27	140
rect	26	142	27	143
rect	27	7	28	8
rect	27	14	28	15
rect	27	16	28	17
rect	27	17	28	18
rect	27	19	28	20
rect	27	20	28	21
rect	27	22	28	23
rect	27	23	28	24
rect	27	25	28	26
rect	27	26	28	27
rect	27	29	28	30
rect	27	34	28	35
rect	27	35	28	36
rect	27	39	28	40
rect	27	42	28	43
rect	27	52	28	53
rect	27	53	28	54
rect	27	54	28	55
rect	27	55	28	56
rect	27	58	28	59
rect	27	59	28	60
rect	27	61	28	62
rect	27	68	28	69
rect	27	71	28	72
rect	27	72	28	73
rect	27	73	28	74
rect	27	74	28	75
rect	27	75	28	76
rect	27	77	28	78
rect	27	81	28	82
rect	27	84	28	85
rect	27	93	28	94
rect	27	96	28	97
rect	27	99	28	100
rect	27	102	28	103
rect	27	112	28	113
rect	27	115	28	116
rect	27	139	28	140
rect	27	142	28	143
rect	28	7	29	8
rect	28	11	29	12
rect	28	14	29	15
rect	28	16	29	17
rect	28	17	29	18
rect	28	19	29	20
rect	28	20	29	21
rect	28	22	29	23
rect	28	23	29	24
rect	28	25	29	26
rect	28	26	29	27
rect	28	29	29	30
rect	28	34	29	35
rect	28	35	29	36
rect	28	39	29	40
rect	28	42	29	43
rect	28	49	29	50
rect	28	52	29	53
rect	28	53	29	54
rect	28	54	29	55
rect	28	55	29	56
rect	28	58	29	59
rect	28	59	29	60
rect	28	61	29	62
rect	28	64	29	65
rect	28	68	29	69
rect	28	71	29	72
rect	28	72	29	73
rect	28	73	29	74
rect	28	74	29	75
rect	28	75	29	76
rect	28	77	29	78
rect	28	80	29	81
rect	28	81	29	82
rect	28	83	29	84
rect	28	84	29	85
rect	28	93	29	94
rect	28	96	29	97
rect	28	99	29	100
rect	28	102	29	103
rect	28	112	29	113
rect	28	115	29	116
rect	28	132	29	133
rect	28	139	29	140
rect	28	142	29	143
rect	29	7	30	8
rect	29	11	30	12
rect	29	14	30	15
rect	29	16	30	17
rect	29	17	30	18
rect	29	19	30	20
rect	29	20	30	21
rect	29	22	30	23
rect	29	23	30	24
rect	29	25	30	26
rect	29	26	30	27
rect	29	29	30	30
rect	29	34	30	35
rect	29	35	30	36
rect	29	39	30	40
rect	29	42	30	43
rect	29	49	30	50
rect	29	52	30	53
rect	29	53	30	54
rect	29	54	30	55
rect	29	55	30	56
rect	29	58	30	59
rect	29	59	30	60
rect	29	61	30	62
rect	29	64	30	65
rect	29	68	30	69
rect	29	71	30	72
rect	29	72	30	73
rect	29	73	30	74
rect	29	74	30	75
rect	29	75	30	76
rect	29	77	30	78
rect	29	81	30	82
rect	29	83	30	84
rect	29	84	30	85
rect	29	93	30	94
rect	29	96	30	97
rect	29	99	30	100
rect	29	102	30	103
rect	29	112	30	113
rect	29	115	30	116
rect	29	132	30	133
rect	29	139	30	140
rect	29	142	30	143
rect	30	4	31	5
rect	30	7	31	8
rect	30	11	31	12
rect	30	14	31	15
rect	30	16	31	17
rect	30	17	31	18
rect	30	19	31	20
rect	30	20	31	21
rect	30	22	31	23
rect	30	23	31	24
rect	30	25	31	26
rect	30	26	31	27
rect	30	29	31	30
rect	30	32	31	33
rect	30	34	31	35
rect	30	35	31	36
rect	30	36	31	37
rect	30	39	31	40
rect	30	42	31	43
rect	30	49	31	50
rect	30	52	31	53
rect	30	53	31	54
rect	30	54	31	55
rect	30	55	31	56
rect	30	58	31	59
rect	30	59	31	60
rect	30	61	31	62
rect	30	64	31	65
rect	30	68	31	69
rect	30	71	31	72
rect	30	72	31	73
rect	30	73	31	74
rect	30	74	31	75
rect	30	75	31	76
rect	30	77	31	78
rect	30	80	31	81
rect	30	81	31	82
rect	30	83	31	84
rect	30	84	31	85
rect	30	87	31	88
rect	30	93	31	94
rect	30	96	31	97
rect	30	99	31	100
rect	30	102	31	103
rect	30	112	31	113
rect	30	115	31	116
rect	30	126	31	127
rect	30	132	31	133
rect	30	139	31	140
rect	30	142	31	143
rect	31	16	32	17
rect	31	17	32	18
rect	31	19	32	20
rect	31	20	32	21
rect	31	22	32	23
rect	31	23	32	24
rect	31	25	32	26
rect	31	26	32	27
rect	31	34	32	35
rect	31	35	32	36
rect	31	53	32	54
rect	31	54	32	55
rect	31	58	32	59
rect	31	59	32	60
rect	31	72	32	73
rect	31	73	32	74
rect	31	74	32	75
rect	31	75	32	76
rect	31	80	32	81
rect	31	81	32	82
rect	31	83	32	84
rect	31	84	32	85
rect	32	16	33	17
rect	32	17	33	18
rect	32	19	33	20
rect	32	20	33	21
rect	32	22	33	23
rect	32	23	33	24
rect	32	25	33	26
rect	32	26	33	27
rect	32	34	33	35
rect	32	35	33	36
rect	32	53	33	54
rect	32	54	33	55
rect	32	58	33	59
rect	32	59	33	60
rect	32	72	33	73
rect	32	73	33	74
rect	32	74	33	75
rect	32	75	33	76
rect	32	80	33	81
rect	32	81	33	82
rect	32	83	33	84
rect	32	84	33	85
rect	33	16	34	17
rect	33	17	34	18
rect	33	19	34	20
rect	33	20	34	21
rect	33	22	34	23
rect	33	23	34	24
rect	33	25	34	26
rect	33	26	34	27
rect	33	34	34	35
rect	33	35	34	36
rect	33	53	34	54
rect	33	54	34	55
rect	33	58	34	59
rect	33	59	34	60
rect	33	72	34	73
rect	33	73	34	74
rect	33	74	34	75
rect	33	75	34	76
rect	33	80	34	81
rect	33	81	34	82
rect	33	83	34	84
rect	33	84	34	85
rect	34	16	35	17
rect	34	17	35	18
rect	34	19	35	20
rect	34	20	35	21
rect	34	22	35	23
rect	34	23	35	24
rect	34	25	35	26
rect	34	26	35	27
rect	34	34	35	35
rect	34	35	35	36
rect	34	53	35	54
rect	34	54	35	55
rect	34	58	35	59
rect	34	59	35	60
rect	34	72	35	73
rect	34	73	35	74
rect	34	74	35	75
rect	34	75	35	76
rect	34	80	35	81
rect	34	81	35	82
rect	34	83	35	84
rect	34	84	35	85
rect	35	16	36	17
rect	35	17	36	18
rect	35	19	36	20
rect	35	20	36	21
rect	35	22	36	23
rect	35	23	36	24
rect	35	25	36	26
rect	35	26	36	27
rect	35	34	36	35
rect	35	35	36	36
rect	35	53	36	54
rect	35	54	36	55
rect	35	58	36	59
rect	35	59	36	60
rect	35	72	36	73
rect	35	73	36	74
rect	35	74	36	75
rect	35	75	36	76
rect	35	80	36	81
rect	35	81	36	82
rect	35	83	36	84
rect	35	84	36	85
rect	36	16	37	17
rect	36	17	37	18
rect	36	19	37	20
rect	36	20	37	21
rect	36	22	37	23
rect	36	23	37	24
rect	36	25	37	26
rect	36	26	37	27
rect	36	34	37	35
rect	36	35	37	36
rect	36	53	37	54
rect	36	54	37	55
rect	36	58	37	59
rect	36	59	37	60
rect	36	72	37	73
rect	36	73	37	74
rect	36	74	37	75
rect	36	75	37	76
rect	36	80	37	81
rect	36	81	37	82
rect	36	83	37	84
rect	36	84	37	85
rect	37	4	38	5
rect	37	7	38	8
rect	37	14	38	15
rect	37	16	38	17
rect	37	17	38	18
rect	37	19	38	20
rect	37	20	38	21
rect	37	22	38	23
rect	37	23	38	24
rect	37	25	38	26
rect	37	26	38	27
rect	37	29	38	30
rect	37	32	38	33
rect	37	34	38	35
rect	37	35	38	36
rect	37	39	38	40
rect	37	42	38	43
rect	37	52	38	53
rect	37	53	38	54
rect	37	54	38	55
rect	37	55	38	56
rect	37	58	38	59
rect	37	59	38	60
rect	37	61	38	62
rect	37	64	38	65
rect	37	68	38	69
rect	37	72	38	73
rect	37	73	38	74
rect	37	74	38	75
rect	37	75	38	76
rect	37	77	38	78
rect	37	80	38	81
rect	37	81	38	82
rect	37	83	38	84
rect	37	84	38	85
rect	37	90	38	91
rect	37	93	38	94
rect	37	96	38	97
rect	37	99	38	100
rect	37	102	38	103
rect	37	112	38	113
rect	37	115	38	116
rect	37	122	38	123
rect	37	129	38	130
rect	37	132	38	133
rect	37	142	38	143
rect	38	4	39	5
rect	38	7	39	8
rect	38	14	39	15
rect	38	16	39	17
rect	38	17	39	18
rect	38	19	39	20
rect	38	20	39	21
rect	38	22	39	23
rect	38	23	39	24
rect	38	25	39	26
rect	38	26	39	27
rect	38	29	39	30
rect	38	32	39	33
rect	38	34	39	35
rect	38	35	39	36
rect	38	39	39	40
rect	38	42	39	43
rect	38	52	39	53
rect	38	53	39	54
rect	38	54	39	55
rect	38	55	39	56
rect	38	59	39	60
rect	38	61	39	62
rect	38	64	39	65
rect	38	68	39	69
rect	38	72	39	73
rect	38	73	39	74
rect	38	74	39	75
rect	38	75	39	76
rect	38	77	39	78
rect	38	80	39	81
rect	38	81	39	82
rect	38	83	39	84
rect	38	84	39	85
rect	38	90	39	91
rect	38	93	39	94
rect	38	96	39	97
rect	38	99	39	100
rect	38	102	39	103
rect	38	112	39	113
rect	38	115	39	116
rect	38	122	39	123
rect	38	129	39	130
rect	38	132	39	133
rect	38	142	39	143
rect	39	4	40	5
rect	39	7	40	8
rect	39	14	40	15
rect	39	16	40	17
rect	39	17	40	18
rect	39	19	40	20
rect	39	20	40	21
rect	39	22	40	23
rect	39	23	40	24
rect	39	25	40	26
rect	39	26	40	27
rect	39	29	40	30
rect	39	32	40	33
rect	39	34	40	35
rect	39	35	40	36
rect	39	39	40	40
rect	39	42	40	43
rect	39	52	40	53
rect	39	53	40	54
rect	39	54	40	55
rect	39	55	40	56
rect	39	58	40	59
rect	39	59	40	60
rect	39	61	40	62
rect	39	64	40	65
rect	39	68	40	69
rect	39	70	40	71
rect	39	72	40	73
rect	39	73	40	74
rect	39	74	40	75
rect	39	75	40	76
rect	39	77	40	78
rect	39	80	40	81
rect	39	81	40	82
rect	39	83	40	84
rect	39	84	40	85
rect	39	90	40	91
rect	39	93	40	94
rect	39	96	40	97
rect	39	99	40	100
rect	39	102	40	103
rect	39	112	40	113
rect	39	115	40	116
rect	39	122	40	123
rect	39	129	40	130
rect	39	132	40	133
rect	39	142	40	143
rect	40	4	41	5
rect	40	7	41	8
rect	40	14	41	15
rect	40	16	41	17
rect	40	17	41	18
rect	40	19	41	20
rect	40	20	41	21
rect	40	22	41	23
rect	40	23	41	24
rect	40	25	41	26
rect	40	26	41	27
rect	40	29	41	30
rect	40	32	41	33
rect	40	34	41	35
rect	40	35	41	36
rect	40	39	41	40
rect	40	42	41	43
rect	40	52	41	53
rect	40	53	41	54
rect	40	54	41	55
rect	40	55	41	56
rect	40	58	41	59
rect	40	59	41	60
rect	40	61	41	62
rect	40	64	41	65
rect	40	70	41	71
rect	40	72	41	73
rect	40	73	41	74
rect	40	74	41	75
rect	40	75	41	76
rect	40	77	41	78
rect	40	80	41	81
rect	40	81	41	82
rect	40	83	41	84
rect	40	84	41	85
rect	40	90	41	91
rect	40	93	41	94
rect	40	96	41	97
rect	40	99	41	100
rect	40	102	41	103
rect	40	112	41	113
rect	40	115	41	116
rect	40	122	41	123
rect	40	129	41	130
rect	40	132	41	133
rect	40	142	41	143
rect	41	4	42	5
rect	41	7	42	8
rect	41	14	42	15
rect	41	16	42	17
rect	41	17	42	18
rect	41	19	42	20
rect	41	20	42	21
rect	41	22	42	23
rect	41	23	42	24
rect	41	25	42	26
rect	41	26	42	27
rect	41	29	42	30
rect	41	32	42	33
rect	41	34	42	35
rect	41	35	42	36
rect	41	39	42	40
rect	41	42	42	43
rect	41	52	42	53
rect	41	53	42	54
rect	41	54	42	55
rect	41	55	42	56
rect	41	58	42	59
rect	41	59	42	60
rect	41	61	42	62
rect	41	64	42	65
rect	41	70	42	71
rect	41	72	42	73
rect	41	73	42	74
rect	41	74	42	75
rect	41	75	42	76
rect	41	77	42	78
rect	41	80	42	81
rect	41	81	42	82
rect	41	83	42	84
rect	41	84	42	85
rect	41	90	42	91
rect	41	93	42	94
rect	41	96	42	97
rect	41	99	42	100
rect	41	102	42	103
rect	41	112	42	113
rect	41	115	42	116
rect	41	122	42	123
rect	41	129	42	130
rect	41	132	42	133
rect	41	142	42	143
rect	42	4	43	5
rect	42	7	43	8
rect	42	14	43	15
rect	42	16	43	17
rect	42	17	43	18
rect	42	19	43	20
rect	42	20	43	21
rect	42	22	43	23
rect	42	23	43	24
rect	42	25	43	26
rect	42	26	43	27
rect	42	29	43	30
rect	42	32	43	33
rect	42	34	43	35
rect	42	35	43	36
rect	42	39	43	40
rect	42	42	43	43
rect	42	52	43	53
rect	42	53	43	54
rect	42	54	43	55
rect	42	58	43	59
rect	42	59	43	60
rect	42	61	43	62
rect	42	64	43	65
rect	42	70	43	71
rect	42	72	43	73
rect	42	73	43	74
rect	42	74	43	75
rect	42	75	43	76
rect	42	77	43	78
rect	42	80	43	81
rect	42	81	43	82
rect	42	83	43	84
rect	42	84	43	85
rect	42	96	43	97
rect	42	99	43	100
rect	42	112	43	113
rect	42	115	43	116
rect	42	122	43	123
rect	42	129	43	130
rect	42	132	43	133
rect	42	142	43	143
rect	43	4	44	5
rect	43	7	44	8
rect	43	14	44	15
rect	43	16	44	17
rect	43	17	44	18
rect	43	19	44	20
rect	43	20	44	21
rect	43	22	44	23
rect	43	23	44	24
rect	43	25	44	26
rect	43	26	44	27
rect	43	29	44	30
rect	43	32	44	33
rect	43	34	44	35
rect	43	35	44	36
rect	43	39	44	40
rect	43	42	44	43
rect	43	52	44	53
rect	43	53	44	54
rect	43	54	44	55
rect	43	58	44	59
rect	43	59	44	60
rect	43	61	44	62
rect	43	64	44	65
rect	43	67	44	68
rect	43	70	44	71
rect	43	72	44	73
rect	43	73	44	74
rect	43	74	44	75
rect	43	75	44	76
rect	43	77	44	78
rect	43	80	44	81
rect	43	81	44	82
rect	43	83	44	84
rect	43	84	44	85
rect	43	96	44	97
rect	43	99	44	100
rect	43	108	44	109
rect	43	112	44	113
rect	43	115	44	116
rect	43	122	44	123
rect	43	129	44	130
rect	43	132	44	133
rect	43	142	44	143
rect	44	4	45	5
rect	44	7	45	8
rect	44	14	45	15
rect	44	16	45	17
rect	44	17	45	18
rect	44	19	45	20
rect	44	20	45	21
rect	44	22	45	23
rect	44	23	45	24
rect	44	25	45	26
rect	44	26	45	27
rect	44	32	45	33
rect	44	34	45	35
rect	44	35	45	36
rect	44	39	45	40
rect	44	42	45	43
rect	44	52	45	53
rect	44	53	45	54
rect	44	54	45	55
rect	44	58	45	59
rect	44	59	45	60
rect	44	64	45	65
rect	44	67	45	68
rect	44	70	45	71
rect	44	72	45	73
rect	44	73	45	74
rect	44	74	45	75
rect	44	75	45	76
rect	44	80	45	81
rect	44	81	45	82
rect	44	83	45	84
rect	44	84	45	85
rect	44	96	45	97
rect	44	108	45	109
rect	44	112	45	113
rect	44	115	45	116
rect	44	122	45	123
rect	44	129	45	130
rect	44	132	45	133
rect	44	142	45	143
rect	45	4	46	5
rect	45	7	46	8
rect	45	10	46	11
rect	45	14	46	15
rect	45	16	46	17
rect	45	17	46	18
rect	45	19	46	20
rect	45	20	46	21
rect	45	22	46	23
rect	45	23	46	24
rect	45	25	46	26
rect	45	26	46	27
rect	45	32	46	33
rect	45	34	46	35
rect	45	35	46	36
rect	45	39	46	40
rect	45	42	46	43
rect	45	45	46	46
rect	45	52	46	53
rect	45	53	46	54
rect	45	54	46	55
rect	45	58	46	59
rect	45	59	46	60
rect	45	64	46	65
rect	45	67	46	68
rect	45	70	46	71
rect	45	72	46	73
rect	45	73	46	74
rect	45	74	46	75
rect	45	75	46	76
rect	45	80	46	81
rect	45	81	46	82
rect	45	83	46	84
rect	45	84	46	85
rect	45	89	46	90
rect	45	96	46	97
rect	45	105	46	106
rect	45	108	46	109
rect	45	112	46	113
rect	45	115	46	116
rect	45	122	46	123
rect	45	129	46	130
rect	45	132	46	133
rect	45	142	46	143
rect	46	4	47	5
rect	46	10	47	11
rect	46	14	47	15
rect	46	16	47	17
rect	46	17	47	18
rect	46	19	47	20
rect	46	20	47	21
rect	46	22	47	23
rect	46	23	47	24
rect	46	25	47	26
rect	46	26	47	27
rect	46	32	47	33
rect	46	34	47	35
rect	46	35	47	36
rect	46	39	47	40
rect	46	42	47	43
rect	46	45	47	46
rect	46	53	47	54
rect	46	54	47	55
rect	46	58	47	59
rect	46	59	47	60
rect	46	67	47	68
rect	46	70	47	71
rect	46	72	47	73
rect	46	73	47	74
rect	46	74	47	75
rect	46	75	47	76
rect	46	80	47	81
rect	46	81	47	82
rect	46	83	47	84
rect	46	84	47	85
rect	46	89	47	90
rect	46	105	47	106
rect	46	108	47	109
rect	46	112	47	113
rect	46	115	47	116
rect	46	129	47	130
rect	46	132	47	133
rect	47	4	48	5
rect	47	10	48	11
rect	47	14	48	15
rect	47	16	48	17
rect	47	17	48	18
rect	47	19	48	20
rect	47	20	48	21
rect	47	22	48	23
rect	47	23	48	24
rect	47	25	48	26
rect	47	26	48	27
rect	47	29	48	30
rect	47	32	48	33
rect	47	34	48	35
rect	47	35	48	36
rect	47	39	48	40
rect	47	42	48	43
rect	47	45	48	46
rect	47	53	48	54
rect	47	54	48	55
rect	47	58	48	59
rect	47	59	48	60
rect	47	61	48	62
rect	47	67	48	68
rect	47	70	48	71
rect	47	72	48	73
rect	47	73	48	74
rect	47	74	48	75
rect	47	75	48	76
rect	47	76	48	77
rect	47	80	48	81
rect	47	81	48	82
rect	47	83	48	84
rect	47	84	48	85
rect	47	89	48	90
rect	47	92	48	93
rect	47	105	48	106
rect	47	108	48	109
rect	47	112	48	113
rect	47	115	48	116
rect	47	129	48	130
rect	47	132	48	133
rect	47	137	48	138
rect	47	147	48	148
rect	47	157	48	158
rect	48	4	49	5
rect	48	10	49	11
rect	48	14	49	15
rect	48	16	49	17
rect	48	17	49	18
rect	48	19	49	20
rect	48	20	49	21
rect	48	22	49	23
rect	48	23	49	24
rect	48	25	49	26
rect	48	26	49	27
rect	48	29	49	30
rect	48	32	49	33
rect	48	34	49	35
rect	48	35	49	36
rect	48	42	49	43
rect	48	45	49	46
rect	48	53	49	54
rect	48	54	49	55
rect	48	58	49	59
rect	48	59	49	60
rect	48	61	49	62
rect	48	67	49	68
rect	48	70	49	71
rect	48	72	49	73
rect	48	73	49	74
rect	48	74	49	75
rect	48	75	49	76
rect	48	76	49	77
rect	48	80	49	81
rect	48	81	49	82
rect	48	83	49	84
rect	48	84	49	85
rect	48	89	49	90
rect	48	92	49	93
rect	48	105	49	106
rect	48	108	49	109
rect	48	112	49	113
rect	48	115	49	116
rect	48	129	49	130
rect	48	132	49	133
rect	48	137	49	138
rect	48	147	49	148
rect	48	157	49	158
rect	49	4	50	5
rect	49	7	50	8
rect	49	10	50	11
rect	49	14	50	15
rect	49	16	50	17
rect	49	17	50	18
rect	49	19	50	20
rect	49	20	50	21
rect	49	22	50	23
rect	49	23	50	24
rect	49	25	50	26
rect	49	26	50	27
rect	49	29	50	30
rect	49	32	50	33
rect	49	34	50	35
rect	49	35	50	36
rect	49	42	50	43
rect	49	45	50	46
rect	49	53	50	54
rect	49	54	50	55
rect	49	58	50	59
rect	49	59	50	60
rect	49	61	50	62
rect	49	67	50	68
rect	49	70	50	71
rect	49	72	50	73
rect	49	73	50	74
rect	49	74	50	75
rect	49	75	50	76
rect	49	76	50	77
rect	49	80	50	81
rect	49	81	50	82
rect	49	83	50	84
rect	49	84	50	85
rect	49	89	50	90
rect	49	92	50	93
rect	49	105	50	106
rect	49	108	50	109
rect	49	112	50	113
rect	49	115	50	116
rect	49	129	50	130
rect	49	132	50	133
rect	49	137	50	138
rect	49	147	50	148
rect	49	157	50	158
rect	49	166	50	167
rect	50	4	51	5
rect	50	7	51	8
rect	50	10	51	11
rect	50	14	51	15
rect	50	16	51	17
rect	50	17	51	18
rect	50	19	51	20
rect	50	20	51	21
rect	50	22	51	23
rect	50	23	51	24
rect	50	25	51	26
rect	50	26	51	27
rect	50	29	51	30
rect	50	34	51	35
rect	50	35	51	36
rect	50	45	51	46
rect	50	53	51	54
rect	50	54	51	55
rect	50	58	51	59
rect	50	59	51	60
rect	50	61	51	62
rect	50	67	51	68
rect	50	70	51	71
rect	50	72	51	73
rect	50	73	51	74
rect	50	74	51	75
rect	50	75	51	76
rect	50	76	51	77
rect	50	80	51	81
rect	50	81	51	82
rect	50	83	51	84
rect	50	84	51	85
rect	50	89	51	90
rect	50	92	51	93
rect	50	105	51	106
rect	50	108	51	109
rect	50	115	51	116
rect	50	129	51	130
rect	50	137	51	138
rect	50	147	51	148
rect	50	157	51	158
rect	50	166	51	167
rect	51	4	52	5
rect	51	7	52	8
rect	51	10	52	11
rect	51	14	52	15
rect	51	16	52	17
rect	51	17	52	18
rect	51	19	52	20
rect	51	20	52	21
rect	51	22	52	23
rect	51	23	52	24
rect	51	25	52	26
rect	51	26	52	27
rect	51	29	52	30
rect	51	34	52	35
rect	51	35	52	36
rect	51	39	52	40
rect	51	45	52	46
rect	51	53	52	54
rect	51	54	52	55
rect	51	58	52	59
rect	51	59	52	60
rect	51	61	52	62
rect	51	64	52	65
rect	51	67	52	68
rect	51	70	52	71
rect	51	72	52	73
rect	51	73	52	74
rect	51	74	52	75
rect	51	75	52	76
rect	51	76	52	77
rect	51	80	52	81
rect	51	81	52	82
rect	51	83	52	84
rect	51	84	52	85
rect	51	89	52	90
rect	51	92	52	93
rect	51	102	52	103
rect	51	105	52	106
rect	51	108	52	109
rect	51	115	52	116
rect	51	124	52	125
rect	51	129	52	130
rect	51	137	52	138
rect	51	147	52	148
rect	51	157	52	158
rect	51	160	52	161
rect	51	166	52	167
rect	52	4	53	5
rect	52	7	53	8
rect	52	10	53	11
rect	52	16	53	17
rect	52	17	53	18
rect	52	19	53	20
rect	52	20	53	21
rect	52	22	53	23
rect	52	23	53	24
rect	52	25	53	26
rect	52	26	53	27
rect	52	29	53	30
rect	52	34	53	35
rect	52	35	53	36
rect	52	39	53	40
rect	52	45	53	46
rect	52	53	53	54
rect	52	54	53	55
rect	52	58	53	59
rect	52	59	53	60
rect	52	61	53	62
rect	52	64	53	65
rect	52	67	53	68
rect	52	70	53	71
rect	52	72	53	73
rect	52	74	53	75
rect	52	75	53	76
rect	52	76	53	77
rect	52	80	53	81
rect	52	81	53	82
rect	52	84	53	85
rect	52	89	53	90
rect	52	92	53	93
rect	52	102	53	103
rect	52	105	53	106
rect	52	108	53	109
rect	52	115	53	116
rect	52	124	53	125
rect	52	129	53	130
rect	52	137	53	138
rect	52	147	53	148
rect	52	157	53	158
rect	52	160	53	161
rect	52	166	53	167
rect	53	4	54	5
rect	53	7	54	8
rect	53	10	54	11
rect	53	16	54	17
rect	53	17	54	18
rect	53	19	54	20
rect	53	20	54	21
rect	53	22	54	23
rect	53	23	54	24
rect	53	25	54	26
rect	53	26	54	27
rect	53	29	54	30
rect	53	33	54	34
rect	53	34	54	35
rect	53	35	54	36
rect	53	39	54	40
rect	53	42	54	43
rect	53	45	54	46
rect	53	49	54	50
rect	53	53	54	54
rect	53	54	54	55
rect	53	55	54	56
rect	53	58	54	59
rect	53	59	54	60
rect	53	61	54	62
rect	53	64	54	65
rect	53	67	54	68
rect	53	70	54	71
rect	53	72	54	73
rect	53	73	54	74
rect	53	74	54	75
rect	53	75	54	76
rect	53	76	54	77
rect	53	80	54	81
rect	53	81	54	82
rect	53	83	54	84
rect	53	84	54	85
rect	53	86	54	87
rect	53	89	54	90
rect	53	92	54	93
rect	53	96	54	97
rect	53	99	54	100
rect	53	102	54	103
rect	53	105	54	106
rect	53	108	54	109
rect	53	115	54	116
rect	53	124	54	125
rect	53	129	54	130
rect	53	137	54	138
rect	53	147	54	148
rect	53	157	54	158
rect	53	160	54	161
rect	53	163	54	164
rect	53	166	54	167
rect	54	7	55	8
rect	54	10	55	11
rect	54	16	55	17
rect	54	17	55	18
rect	54	19	55	20
rect	54	22	55	23
rect	54	23	55	24
rect	54	25	55	26
rect	54	26	55	27
rect	54	29	55	30
rect	54	33	55	34
rect	54	34	55	35
rect	54	35	55	36
rect	54	39	55	40
rect	54	42	55	43
rect	54	45	55	46
rect	54	49	55	50
rect	54	53	55	54
rect	54	54	55	55
rect	54	55	55	56
rect	54	58	55	59
rect	54	59	55	60
rect	54	61	55	62
rect	54	64	55	65
rect	54	67	55	68
rect	54	70	55	71
rect	54	72	55	73
rect	54	73	55	74
rect	54	74	55	75
rect	54	75	55	76
rect	54	76	55	77
rect	54	80	55	81
rect	54	81	55	82
rect	54	83	55	84
rect	54	84	55	85
rect	54	86	55	87
rect	54	89	55	90
rect	54	92	55	93
rect	54	96	55	97
rect	54	99	55	100
rect	54	102	55	103
rect	54	105	55	106
rect	54	108	55	109
rect	54	124	55	125
rect	54	137	55	138
rect	54	147	55	148
rect	54	157	55	158
rect	54	160	55	161
rect	54	163	55	164
rect	54	166	55	167
rect	55	7	56	8
rect	55	10	56	11
rect	55	13	56	14
rect	55	16	56	17
rect	55	17	56	18
rect	55	19	56	20
rect	55	20	56	21
rect	55	22	56	23
rect	55	23	56	24
rect	55	25	56	26
rect	55	26	56	27
rect	55	29	56	30
rect	55	33	56	34
rect	55	34	56	35
rect	55	35	56	36
rect	55	39	56	40
rect	55	42	56	43
rect	55	45	56	46
rect	55	49	56	50
rect	55	53	56	54
rect	55	54	56	55
rect	55	55	56	56
rect	55	58	56	59
rect	55	59	56	60
rect	55	61	56	62
rect	55	64	56	65
rect	55	67	56	68
rect	55	70	56	71
rect	55	72	56	73
rect	55	73	56	74
rect	55	74	56	75
rect	55	75	56	76
rect	55	76	56	77
rect	55	80	56	81
rect	55	81	56	82
rect	55	83	56	84
rect	55	84	56	85
rect	55	86	56	87
rect	55	89	56	90
rect	55	92	56	93
rect	55	96	56	97
rect	55	99	56	100
rect	55	102	56	103
rect	55	105	56	106
rect	55	108	56	109
rect	55	111	56	112
rect	55	121	56	122
rect	55	124	56	125
rect	55	134	56	135
rect	55	137	56	138
rect	55	141	56	142
rect	55	147	56	148
rect	55	150	56	151
rect	55	157	56	158
rect	55	160	56	161
rect	55	163	56	164
rect	55	166	56	167
rect	56	16	57	17
rect	56	17	57	18
rect	56	19	57	20
rect	56	20	57	21
rect	56	22	57	23
rect	56	23	57	24
rect	56	25	57	26
rect	56	26	57	27
rect	56	34	57	35
rect	56	35	57	36
rect	56	53	57	54
rect	56	54	57	55
rect	56	58	57	59
rect	56	59	57	60
rect	56	72	57	73
rect	56	73	57	74
rect	56	74	57	75
rect	56	75	57	76
rect	56	80	57	81
rect	56	81	57	82
rect	56	83	57	84
rect	56	84	57	85
rect	57	16	58	17
rect	57	17	58	18
rect	57	19	58	20
rect	57	20	58	21
rect	57	22	58	23
rect	57	23	58	24
rect	57	25	58	26
rect	57	26	58	27
rect	57	34	58	35
rect	57	35	58	36
rect	57	53	58	54
rect	57	54	58	55
rect	57	58	58	59
rect	57	59	58	60
rect	57	72	58	73
rect	57	73	58	74
rect	57	74	58	75
rect	57	75	58	76
rect	57	80	58	81
rect	57	81	58	82
rect	57	83	58	84
rect	57	84	58	85
rect	58	16	59	17
rect	58	17	59	18
rect	58	19	59	20
rect	58	20	59	21
rect	58	22	59	23
rect	58	23	59	24
rect	58	25	59	26
rect	58	26	59	27
rect	58	34	59	35
rect	58	35	59	36
rect	58	53	59	54
rect	58	54	59	55
rect	58	58	59	59
rect	58	59	59	60
rect	58	72	59	73
rect	58	73	59	74
rect	58	74	59	75
rect	58	75	59	76
rect	58	80	59	81
rect	58	81	59	82
rect	58	83	59	84
rect	58	84	59	85
rect	59	16	60	17
rect	59	17	60	18
rect	59	19	60	20
rect	59	20	60	21
rect	59	22	60	23
rect	59	23	60	24
rect	59	25	60	26
rect	59	26	60	27
rect	59	34	60	35
rect	59	35	60	36
rect	59	53	60	54
rect	59	54	60	55
rect	59	58	60	59
rect	59	59	60	60
rect	59	72	60	73
rect	59	73	60	74
rect	59	74	60	75
rect	59	75	60	76
rect	59	80	60	81
rect	59	81	60	82
rect	59	83	60	84
rect	59	84	60	85
rect	60	16	61	17
rect	60	17	61	18
rect	60	19	61	20
rect	60	20	61	21
rect	60	22	61	23
rect	60	23	61	24
rect	60	25	61	26
rect	60	26	61	27
rect	60	34	61	35
rect	60	35	61	36
rect	60	53	61	54
rect	60	54	61	55
rect	60	58	61	59
rect	60	59	61	60
rect	60	72	61	73
rect	60	73	61	74
rect	60	74	61	75
rect	60	75	61	76
rect	60	80	61	81
rect	60	81	61	82
rect	60	83	61	84
rect	60	84	61	85
rect	61	16	62	17
rect	61	17	62	18
rect	61	19	62	20
rect	61	20	62	21
rect	61	22	62	23
rect	61	23	62	24
rect	61	25	62	26
rect	61	26	62	27
rect	61	34	62	35
rect	61	35	62	36
rect	61	53	62	54
rect	61	54	62	55
rect	61	58	62	59
rect	61	59	62	60
rect	61	72	62	73
rect	61	73	62	74
rect	61	74	62	75
rect	61	75	62	76
rect	61	80	62	81
rect	61	81	62	82
rect	61	83	62	84
rect	61	84	62	85
rect	62	1	63	2
rect	62	7	63	8
rect	62	10	63	11
rect	62	13	63	14
rect	62	16	63	17
rect	62	17	63	18
rect	62	19	63	20
rect	62	20	63	21
rect	62	22	63	23
rect	62	23	63	24
rect	62	25	63	26
rect	62	26	63	27
rect	62	29	63	30
rect	62	34	63	35
rect	62	35	63	36
rect	62	39	63	40
rect	62	42	63	43
rect	62	45	63	46
rect	62	49	63	50
rect	62	53	63	54
rect	62	54	63	55
rect	62	55	63	56
rect	62	58	63	59
rect	62	59	63	60
rect	62	61	63	62
rect	62	64	63	65
rect	62	67	63	68
rect	62	70	63	71
rect	62	72	63	73
rect	62	73	63	74
rect	62	74	63	75
rect	62	75	63	76
rect	62	76	63	77
rect	62	80	63	81
rect	62	81	63	82
rect	62	83	63	84
rect	62	84	63	85
rect	62	86	63	87
rect	62	89	63	90
rect	62	92	63	93
rect	62	102	63	103
rect	62	105	63	106
rect	62	108	63	109
rect	62	111	63	112
rect	62	115	63	116
rect	62	121	63	122
rect	62	124	63	125
rect	62	128	63	129
rect	62	134	63	135
rect	62	137	63	138
rect	62	147	63	148
rect	62	150	63	151
rect	62	154	63	155
rect	62	160	63	161
rect	62	163	63	164
rect	62	166	63	167
rect	63	1	64	2
rect	63	7	64	8
rect	63	10	64	11
rect	63	13	64	14
rect	63	16	64	17
rect	63	17	64	18
rect	63	19	64	20
rect	63	20	64	21
rect	63	22	64	23
rect	63	23	64	24
rect	63	25	64	26
rect	63	26	64	27
rect	63	29	64	30
rect	63	34	64	35
rect	63	35	64	36
rect	63	39	64	40
rect	63	42	64	43
rect	63	45	64	46
rect	63	49	64	50
rect	63	53	64	54
rect	63	54	64	55
rect	63	55	64	56
rect	63	58	64	59
rect	63	59	64	60
rect	63	61	64	62
rect	63	64	64	65
rect	63	67	64	68
rect	63	70	64	71
rect	63	72	64	73
rect	63	73	64	74
rect	63	74	64	75
rect	63	75	64	76
rect	63	76	64	77
rect	63	80	64	81
rect	63	81	64	82
rect	63	83	64	84
rect	63	84	64	85
rect	63	86	64	87
rect	63	89	64	90
rect	63	92	64	93
rect	63	102	64	103
rect	63	105	64	106
rect	63	108	64	109
rect	63	111	64	112
rect	63	115	64	116
rect	63	121	64	122
rect	63	124	64	125
rect	63	128	64	129
rect	63	134	64	135
rect	63	137	64	138
rect	63	147	64	148
rect	63	150	64	151
rect	63	154	64	155
rect	63	160	64	161
rect	63	163	64	164
rect	64	1	65	2
rect	64	7	65	8
rect	64	10	65	11
rect	64	13	65	14
rect	64	16	65	17
rect	64	17	65	18
rect	64	19	65	20
rect	64	20	65	21
rect	64	22	65	23
rect	64	23	65	24
rect	64	25	65	26
rect	64	26	65	27
rect	64	29	65	30
rect	64	34	65	35
rect	64	35	65	36
rect	64	39	65	40
rect	64	42	65	43
rect	64	45	65	46
rect	64	49	65	50
rect	64	53	65	54
rect	64	54	65	55
rect	64	55	65	56
rect	64	58	65	59
rect	64	59	65	60
rect	64	61	65	62
rect	64	64	65	65
rect	64	67	65	68
rect	64	70	65	71
rect	64	72	65	73
rect	64	73	65	74
rect	64	74	65	75
rect	64	75	65	76
rect	64	76	65	77
rect	64	80	65	81
rect	64	81	65	82
rect	64	83	65	84
rect	64	84	65	85
rect	64	86	65	87
rect	64	89	65	90
rect	64	92	65	93
rect	64	102	65	103
rect	64	105	65	106
rect	64	108	65	109
rect	64	111	65	112
rect	64	115	65	116
rect	64	121	65	122
rect	64	124	65	125
rect	64	128	65	129
rect	64	134	65	135
rect	64	137	65	138
rect	64	147	65	148
rect	64	150	65	151
rect	64	154	65	155
rect	64	160	65	161
rect	64	163	65	164
rect	64	178	65	179
rect	65	1	66	2
rect	65	7	66	8
rect	65	10	66	11
rect	65	13	66	14
rect	65	16	66	17
rect	65	17	66	18
rect	65	19	66	20
rect	65	20	66	21
rect	65	22	66	23
rect	65	23	66	24
rect	65	25	66	26
rect	65	26	66	27
rect	65	29	66	30
rect	65	34	66	35
rect	65	35	66	36
rect	65	39	66	40
rect	65	42	66	43
rect	65	45	66	46
rect	65	49	66	50
rect	65	53	66	54
rect	65	54	66	55
rect	65	55	66	56
rect	65	58	66	59
rect	65	59	66	60
rect	65	61	66	62
rect	65	64	66	65
rect	65	67	66	68
rect	65	70	66	71
rect	65	72	66	73
rect	65	73	66	74
rect	65	74	66	75
rect	65	75	66	76
rect	65	76	66	77
rect	65	80	66	81
rect	65	81	66	82
rect	65	83	66	84
rect	65	84	66	85
rect	65	86	66	87
rect	65	89	66	90
rect	65	92	66	93
rect	65	102	66	103
rect	65	105	66	106
rect	65	108	66	109
rect	65	111	66	112
rect	65	121	66	122
rect	65	124	66	125
rect	65	128	66	129
rect	65	134	66	135
rect	65	137	66	138
rect	65	147	66	148
rect	65	150	66	151
rect	65	154	66	155
rect	65	160	66	161
rect	65	163	66	164
rect	65	178	66	179
rect	66	1	67	2
rect	66	7	67	8
rect	66	10	67	11
rect	66	13	67	14
rect	66	16	67	17
rect	66	17	67	18
rect	66	19	67	20
rect	66	20	67	21
rect	66	22	67	23
rect	66	23	67	24
rect	66	25	67	26
rect	66	26	67	27
rect	66	29	67	30
rect	66	34	67	35
rect	66	35	67	36
rect	66	39	67	40
rect	66	42	67	43
rect	66	45	67	46
rect	66	49	67	50
rect	66	53	67	54
rect	66	54	67	55
rect	66	55	67	56
rect	66	58	67	59
rect	66	59	67	60
rect	66	61	67	62
rect	66	64	67	65
rect	66	67	67	68
rect	66	70	67	71
rect	66	72	67	73
rect	66	73	67	74
rect	66	74	67	75
rect	66	75	67	76
rect	66	76	67	77
rect	66	80	67	81
rect	66	81	67	82
rect	66	83	67	84
rect	66	84	67	85
rect	66	86	67	87
rect	66	89	67	90
rect	66	92	67	93
rect	66	102	67	103
rect	66	105	67	106
rect	66	108	67	109
rect	66	111	67	112
rect	66	121	67	122
rect	66	124	67	125
rect	66	128	67	129
rect	66	134	67	135
rect	66	137	67	138
rect	66	147	67	148
rect	66	150	67	151
rect	66	154	67	155
rect	66	160	67	161
rect	66	163	67	164
rect	66	166	67	167
rect	66	178	67	179
rect	67	1	68	2
rect	67	7	68	8
rect	67	10	68	11
rect	67	13	68	14
rect	67	16	68	17
rect	67	17	68	18
rect	67	19	68	20
rect	67	20	68	21
rect	67	22	68	23
rect	67	23	68	24
rect	67	25	68	26
rect	67	26	68	27
rect	67	29	68	30
rect	67	34	68	35
rect	67	35	68	36
rect	67	39	68	40
rect	67	42	68	43
rect	67	45	68	46
rect	67	49	68	50
rect	67	53	68	54
rect	67	54	68	55
rect	67	55	68	56
rect	67	58	68	59
rect	67	59	68	60
rect	67	61	68	62
rect	67	64	68	65
rect	67	67	68	68
rect	67	70	68	71
rect	67	72	68	73
rect	67	73	68	74
rect	67	74	68	75
rect	67	75	68	76
rect	67	76	68	77
rect	67	80	68	81
rect	67	81	68	82
rect	67	83	68	84
rect	67	84	68	85
rect	67	86	68	87
rect	67	89	68	90
rect	67	92	68	93
rect	67	102	68	103
rect	67	105	68	106
rect	67	108	68	109
rect	67	121	68	122
rect	67	124	68	125
rect	67	128	68	129
rect	67	134	68	135
rect	67	137	68	138
rect	67	147	68	148
rect	67	150	68	151
rect	67	154	68	155
rect	67	160	68	161
rect	67	163	68	164
rect	67	166	68	167
rect	67	178	68	179
rect	68	1	69	2
rect	68	7	69	8
rect	68	10	69	11
rect	68	13	69	14
rect	68	16	69	17
rect	68	17	69	18
rect	68	19	69	20
rect	68	20	69	21
rect	68	22	69	23
rect	68	23	69	24
rect	68	25	69	26
rect	68	26	69	27
rect	68	29	69	30
rect	68	34	69	35
rect	68	35	69	36
rect	68	39	69	40
rect	68	42	69	43
rect	68	45	69	46
rect	68	49	69	50
rect	68	53	69	54
rect	68	54	69	55
rect	68	55	69	56
rect	68	58	69	59
rect	68	59	69	60
rect	68	61	69	62
rect	68	64	69	65
rect	68	67	69	68
rect	68	70	69	71
rect	68	72	69	73
rect	68	73	69	74
rect	68	74	69	75
rect	68	75	69	76
rect	68	76	69	77
rect	68	80	69	81
rect	68	81	69	82
rect	68	83	69	84
rect	68	84	69	85
rect	68	86	69	87
rect	68	89	69	90
rect	68	92	69	93
rect	68	102	69	103
rect	68	105	69	106
rect	68	108	69	109
rect	68	115	69	116
rect	68	121	69	122
rect	68	124	69	125
rect	68	128	69	129
rect	68	134	69	135
rect	68	137	69	138
rect	68	147	69	148
rect	68	150	69	151
rect	68	154	69	155
rect	68	160	69	161
rect	68	163	69	164
rect	68	166	69	167
rect	68	178	69	179
rect	69	1	70	2
rect	69	7	70	8
rect	69	10	70	11
rect	69	13	70	14
rect	69	16	70	17
rect	69	17	70	18
rect	69	19	70	20
rect	69	20	70	21
rect	69	22	70	23
rect	69	23	70	24
rect	69	25	70	26
rect	69	26	70	27
rect	69	29	70	30
rect	69	34	70	35
rect	69	35	70	36
rect	69	39	70	40
rect	69	42	70	43
rect	69	45	70	46
rect	69	49	70	50
rect	69	53	70	54
rect	69	54	70	55
rect	69	55	70	56
rect	69	58	70	59
rect	69	59	70	60
rect	69	61	70	62
rect	69	64	70	65
rect	69	67	70	68
rect	69	70	70	71
rect	69	72	70	73
rect	69	73	70	74
rect	69	74	70	75
rect	69	75	70	76
rect	69	76	70	77
rect	69	80	70	81
rect	69	81	70	82
rect	69	83	70	84
rect	69	84	70	85
rect	69	86	70	87
rect	69	89	70	90
rect	69	92	70	93
rect	69	102	70	103
rect	69	105	70	106
rect	69	115	70	116
rect	69	121	70	122
rect	69	124	70	125
rect	69	128	70	129
rect	69	134	70	135
rect	69	137	70	138
rect	69	147	70	148
rect	69	150	70	151
rect	69	160	70	161
rect	69	163	70	164
rect	69	166	70	167
rect	69	178	70	179
rect	70	1	71	2
rect	70	7	71	8
rect	70	10	71	11
rect	70	13	71	14
rect	70	16	71	17
rect	70	17	71	18
rect	70	19	71	20
rect	70	20	71	21
rect	70	22	71	23
rect	70	23	71	24
rect	70	25	71	26
rect	70	26	71	27
rect	70	29	71	30
rect	70	34	71	35
rect	70	35	71	36
rect	70	39	71	40
rect	70	42	71	43
rect	70	45	71	46
rect	70	49	71	50
rect	70	53	71	54
rect	70	54	71	55
rect	70	55	71	56
rect	70	58	71	59
rect	70	59	71	60
rect	70	61	71	62
rect	70	64	71	65
rect	70	67	71	68
rect	70	70	71	71
rect	70	72	71	73
rect	70	73	71	74
rect	70	74	71	75
rect	70	75	71	76
rect	70	76	71	77
rect	70	80	71	81
rect	70	81	71	82
rect	70	83	71	84
rect	70	84	71	85
rect	70	86	71	87
rect	70	89	71	90
rect	70	92	71	93
rect	70	102	71	103
rect	70	105	71	106
rect	70	112	71	113
rect	70	115	71	116
rect	70	121	71	122
rect	70	124	71	125
rect	70	128	71	129
rect	70	134	71	135
rect	70	137	71	138
rect	70	147	71	148
rect	70	150	71	151
rect	70	160	71	161
rect	70	163	71	164
rect	70	166	71	167
rect	70	178	71	179
rect	70	208	71	209
rect	71	1	72	2
rect	71	7	72	8
rect	71	10	72	11
rect	71	13	72	14
rect	71	16	72	17
rect	71	17	72	18
rect	71	19	72	20
rect	71	20	72	21
rect	71	22	72	23
rect	71	23	72	24
rect	71	25	72	26
rect	71	26	72	27
rect	71	29	72	30
rect	71	34	72	35
rect	71	35	72	36
rect	71	39	72	40
rect	71	42	72	43
rect	71	45	72	46
rect	71	49	72	50
rect	71	53	72	54
rect	71	54	72	55
rect	71	55	72	56
rect	71	58	72	59
rect	71	59	72	60
rect	71	64	72	65
rect	71	67	72	68
rect	71	70	72	71
rect	71	72	72	73
rect	71	73	72	74
rect	71	74	72	75
rect	71	75	72	76
rect	71	76	72	77
rect	71	80	72	81
rect	71	81	72	82
rect	71	83	72	84
rect	71	84	72	85
rect	71	86	72	87
rect	71	89	72	90
rect	71	92	72	93
rect	71	102	72	103
rect	71	112	72	113
rect	71	115	72	116
rect	71	121	72	122
rect	71	124	72	125
rect	71	128	72	129
rect	71	137	72	138
rect	71	147	72	148
rect	71	150	72	151
rect	71	160	72	161
rect	71	163	72	164
rect	71	166	72	167
rect	71	178	72	179
rect	71	208	72	209
rect	72	1	73	2
rect	72	7	73	8
rect	72	10	73	11
rect	72	13	73	14
rect	72	16	73	17
rect	72	17	73	18
rect	72	19	73	20
rect	72	20	73	21
rect	72	22	73	23
rect	72	23	73	24
rect	72	25	73	26
rect	72	26	73	27
rect	72	29	73	30
rect	72	34	73	35
rect	72	35	73	36
rect	72	39	73	40
rect	72	42	73	43
rect	72	45	73	46
rect	72	49	73	50
rect	72	53	73	54
rect	72	54	73	55
rect	72	55	73	56
rect	72	58	73	59
rect	72	59	73	60
rect	72	64	73	65
rect	72	67	73	68
rect	72	70	73	71
rect	72	72	73	73
rect	72	73	73	74
rect	72	74	73	75
rect	72	75	73	76
rect	72	76	73	77
rect	72	80	73	81
rect	72	81	73	82
rect	72	83	73	84
rect	72	84	73	85
rect	72	86	73	87
rect	72	89	73	90
rect	72	92	73	93
rect	72	102	73	103
rect	72	109	73	110
rect	72	112	73	113
rect	72	115	73	116
rect	72	121	73	122
rect	72	124	73	125
rect	72	128	73	129
rect	72	137	73	138
rect	72	147	73	148
rect	72	150	73	151
rect	72	153	73	154
rect	72	160	73	161
rect	72	163	73	164
rect	72	166	73	167
rect	72	178	73	179
rect	72	208	73	209
rect	73	1	74	2
rect	73	7	74	8
rect	73	10	74	11
rect	73	13	74	14
rect	73	16	74	17
rect	73	17	74	18
rect	73	19	74	20
rect	73	20	74	21
rect	73	22	74	23
rect	73	23	74	24
rect	73	25	74	26
rect	73	26	74	27
rect	73	29	74	30
rect	73	34	74	35
rect	73	35	74	36
rect	73	39	74	40
rect	73	42	74	43
rect	73	45	74	46
rect	73	49	74	50
rect	73	53	74	54
rect	73	54	74	55
rect	73	55	74	56
rect	73	58	74	59
rect	73	59	74	60
rect	73	64	74	65
rect	73	67	74	68
rect	73	70	74	71
rect	73	72	74	73
rect	73	73	74	74
rect	73	74	74	75
rect	73	75	74	76
rect	73	80	74	81
rect	73	81	74	82
rect	73	84	74	85
rect	73	86	74	87
rect	73	89	74	90
rect	73	92	74	93
rect	73	109	74	110
rect	73	112	74	113
rect	73	115	74	116
rect	73	121	74	122
rect	73	124	74	125
rect	73	128	74	129
rect	73	137	74	138
rect	73	147	74	148
rect	73	150	74	151
rect	73	153	74	154
rect	73	160	74	161
rect	73	163	74	164
rect	73	166	74	167
rect	73	178	74	179
rect	73	208	74	209
rect	74	1	75	2
rect	74	7	75	8
rect	74	10	75	11
rect	74	13	75	14
rect	74	16	75	17
rect	74	17	75	18
rect	74	19	75	20
rect	74	20	75	21
rect	74	22	75	23
rect	74	23	75	24
rect	74	25	75	26
rect	74	26	75	27
rect	74	29	75	30
rect	74	34	75	35
rect	74	35	75	36
rect	74	39	75	40
rect	74	42	75	43
rect	74	45	75	46
rect	74	49	75	50
rect	74	53	75	54
rect	74	54	75	55
rect	74	55	75	56
rect	74	58	75	59
rect	74	59	75	60
rect	74	64	75	65
rect	74	67	75	68
rect	74	70	75	71
rect	74	72	75	73
rect	74	73	75	74
rect	74	74	75	75
rect	74	75	75	76
rect	74	80	75	81
rect	74	81	75	82
rect	74	83	75	84
rect	74	84	75	85
rect	74	86	75	87
rect	74	89	75	90
rect	74	92	75	93
rect	74	109	75	110
rect	74	112	75	113
rect	74	115	75	116
rect	74	121	75	122
rect	74	124	75	125
rect	74	128	75	129
rect	74	134	75	135
rect	74	137	75	138
rect	74	147	75	148
rect	74	150	75	151
rect	74	153	75	154
rect	74	160	75	161
rect	74	163	75	164
rect	74	166	75	167
rect	74	178	75	179
rect	74	208	75	209
rect	75	1	76	2
rect	75	7	76	8
rect	75	10	76	11
rect	75	13	76	14
rect	75	16	76	17
rect	75	17	76	18
rect	75	19	76	20
rect	75	20	76	21
rect	75	22	76	23
rect	75	23	76	24
rect	75	25	76	26
rect	75	26	76	27
rect	75	29	76	30
rect	75	34	76	35
rect	75	35	76	36
rect	75	39	76	40
rect	75	42	76	43
rect	75	45	76	46
rect	75	49	76	50
rect	75	53	76	54
rect	75	54	76	55
rect	75	55	76	56
rect	75	58	76	59
rect	75	59	76	60
rect	75	64	76	65
rect	75	67	76	68
rect	75	70	76	71
rect	75	72	76	73
rect	75	74	76	75
rect	75	75	76	76
rect	75	81	76	82
rect	75	83	76	84
rect	75	84	76	85
rect	75	86	76	87
rect	75	89	76	90
rect	75	109	76	110
rect	75	112	76	113
rect	75	115	76	116
rect	75	121	76	122
rect	75	128	76	129
rect	75	134	76	135
rect	75	137	76	138
rect	75	150	76	151
rect	75	153	76	154
rect	75	160	76	161
rect	75	163	76	164
rect	75	166	76	167
rect	75	178	76	179
rect	75	208	76	209
rect	76	1	77	2
rect	76	7	77	8
rect	76	10	77	11
rect	76	13	77	14
rect	76	16	77	17
rect	76	17	77	18
rect	76	19	77	20
rect	76	20	77	21
rect	76	22	77	23
rect	76	23	77	24
rect	76	25	77	26
rect	76	26	77	27
rect	76	29	77	30
rect	76	34	77	35
rect	76	35	77	36
rect	76	39	77	40
rect	76	42	77	43
rect	76	45	77	46
rect	76	49	77	50
rect	76	53	77	54
rect	76	54	77	55
rect	76	55	77	56
rect	76	58	77	59
rect	76	59	77	60
rect	76	64	77	65
rect	76	67	77	68
rect	76	70	77	71
rect	76	72	77	73
rect	76	73	77	74
rect	76	74	77	75
rect	76	75	77	76
rect	76	80	77	81
rect	76	81	77	82
rect	76	83	77	84
rect	76	84	77	85
rect	76	86	77	87
rect	76	89	77	90
rect	76	106	77	107
rect	76	109	77	110
rect	76	112	77	113
rect	76	115	77	116
rect	76	121	77	122
rect	76	128	77	129
rect	76	134	77	135
rect	76	137	77	138
rect	76	140	77	141
rect	76	150	77	151
rect	76	153	77	154
rect	76	156	77	157
rect	76	160	77	161
rect	76	163	77	164
rect	76	166	77	167
rect	76	178	77	179
rect	76	208	77	209
rect	77	1	78	2
rect	77	7	78	8
rect	77	10	78	11
rect	77	13	78	14
rect	77	16	78	17
rect	77	17	78	18
rect	77	19	78	20
rect	77	20	78	21
rect	77	22	78	23
rect	77	23	78	24
rect	77	25	78	26
rect	77	26	78	27
rect	77	29	78	30
rect	77	34	78	35
rect	77	35	78	36
rect	77	39	78	40
rect	77	42	78	43
rect	77	45	78	46
rect	77	49	78	50
rect	77	53	78	54
rect	77	54	78	55
rect	77	55	78	56
rect	77	58	78	59
rect	77	59	78	60
rect	77	64	78	65
rect	77	67	78	68
rect	77	72	78	73
rect	77	73	78	74
rect	77	74	78	75
rect	77	75	78	76
rect	77	80	78	81
rect	77	81	78	82
rect	77	83	78	84
rect	77	84	78	85
rect	77	86	78	87
rect	77	106	78	107
rect	77	109	78	110
rect	77	112	78	113
rect	77	115	78	116
rect	77	121	78	122
rect	77	128	78	129
rect	77	134	78	135
rect	77	137	78	138
rect	77	140	78	141
rect	77	150	78	151
rect	77	153	78	154
rect	77	156	78	157
rect	77	160	78	161
rect	77	163	78	164
rect	77	166	78	167
rect	77	178	78	179
rect	77	208	78	209
rect	78	1	79	2
rect	78	7	79	8
rect	78	10	79	11
rect	78	13	79	14
rect	78	16	79	17
rect	78	17	79	18
rect	78	19	79	20
rect	78	20	79	21
rect	78	22	79	23
rect	78	23	79	24
rect	78	25	79	26
rect	78	26	79	27
rect	78	29	79	30
rect	78	34	79	35
rect	78	35	79	36
rect	78	39	79	40
rect	78	42	79	43
rect	78	45	79	46
rect	78	49	79	50
rect	78	53	79	54
rect	78	54	79	55
rect	78	55	79	56
rect	78	58	79	59
rect	78	59	79	60
rect	78	64	79	65
rect	78	67	79	68
rect	78	72	79	73
rect	78	73	79	74
rect	78	74	79	75
rect	78	75	79	76
rect	78	77	79	78
rect	78	80	79	81
rect	78	81	79	82
rect	78	83	79	84
rect	78	84	79	85
rect	78	86	79	87
rect	78	103	79	104
rect	78	106	79	107
rect	78	109	79	110
rect	78	112	79	113
rect	78	115	79	116
rect	78	121	79	122
rect	78	125	79	126
rect	78	128	79	129
rect	78	134	79	135
rect	78	137	79	138
rect	78	140	79	141
rect	78	147	79	148
rect	78	150	79	151
rect	78	153	79	154
rect	78	156	79	157
rect	78	160	79	161
rect	78	163	79	164
rect	78	166	79	167
rect	78	178	79	179
rect	78	208	79	209
rect	79	1	80	2
rect	79	7	80	8
rect	79	10	80	11
rect	79	13	80	14
rect	79	16	80	17
rect	79	17	80	18
rect	79	19	80	20
rect	79	20	80	21
rect	79	22	80	23
rect	79	23	80	24
rect	79	25	80	26
rect	79	26	80	27
rect	79	29	80	30
rect	79	34	80	35
rect	79	35	80	36
rect	79	39	80	40
rect	79	42	80	43
rect	79	45	80	46
rect	79	49	80	50
rect	79	53	80	54
rect	79	54	80	55
rect	79	55	80	56
rect	79	58	80	59
rect	79	59	80	60
rect	79	64	80	65
rect	79	72	80	73
rect	79	73	80	74
rect	79	74	80	75
rect	79	75	80	76
rect	79	77	80	78
rect	79	80	80	81
rect	79	81	80	82
rect	79	83	80	84
rect	79	84	80	85
rect	79	103	80	104
rect	79	106	80	107
rect	79	109	80	110
rect	79	112	80	113
rect	79	115	80	116
rect	79	121	80	122
rect	79	125	80	126
rect	79	128	80	129
rect	79	134	80	135
rect	79	137	80	138
rect	79	140	80	141
rect	79	147	80	148
rect	79	150	80	151
rect	79	153	80	154
rect	79	156	80	157
rect	79	160	80	161
rect	79	163	80	164
rect	79	166	80	167
rect	79	178	80	179
rect	79	208	80	209
rect	80	1	81	2
rect	80	7	81	8
rect	80	10	81	11
rect	80	13	81	14
rect	80	16	81	17
rect	80	17	81	18
rect	80	19	81	20
rect	80	20	81	21
rect	80	22	81	23
rect	80	23	81	24
rect	80	25	81	26
rect	80	26	81	27
rect	80	29	81	30
rect	80	34	81	35
rect	80	35	81	36
rect	80	39	81	40
rect	80	42	81	43
rect	80	45	81	46
rect	80	49	81	50
rect	80	53	81	54
rect	80	54	81	55
rect	80	55	81	56
rect	80	58	81	59
rect	80	59	81	60
rect	80	64	81	65
rect	80	72	81	73
rect	80	73	81	74
rect	80	74	81	75
rect	80	75	81	76
rect	80	77	81	78
rect	80	80	81	81
rect	80	81	81	82
rect	80	83	81	84
rect	80	84	81	85
rect	80	93	81	94
rect	80	97	81	98
rect	80	103	81	104
rect	80	106	81	107
rect	80	109	81	110
rect	80	112	81	113
rect	80	115	81	116
rect	80	121	81	122
rect	80	125	81	126
rect	80	128	81	129
rect	80	134	81	135
rect	80	137	81	138
rect	80	140	81	141
rect	80	147	81	148
rect	80	150	81	151
rect	80	153	81	154
rect	80	156	81	157
rect	80	160	81	161
rect	80	163	81	164
rect	80	166	81	167
rect	80	169	81	170
rect	80	178	81	179
rect	80	208	81	209
rect	81	1	82	2
rect	81	7	82	8
rect	81	10	82	11
rect	81	13	82	14
rect	81	16	82	17
rect	81	19	82	20
rect	81	20	82	21
rect	81	22	82	23
rect	81	23	82	24
rect	81	25	82	26
rect	81	26	82	27
rect	81	34	82	35
rect	81	35	82	36
rect	81	39	82	40
rect	81	45	82	46
rect	81	49	82	50
rect	81	53	82	54
rect	81	54	82	55
rect	81	55	82	56
rect	81	58	82	59
rect	81	59	82	60
rect	81	72	82	73
rect	81	73	82	74
rect	81	74	82	75
rect	81	75	82	76
rect	81	77	82	78
rect	81	80	82	81
rect	81	81	82	82
rect	81	83	82	84
rect	81	84	82	85
rect	81	93	82	94
rect	81	97	82	98
rect	81	103	82	104
rect	81	106	82	107
rect	81	109	82	110
rect	81	112	82	113
rect	81	115	82	116
rect	81	121	82	122
rect	81	125	82	126
rect	81	134	82	135
rect	81	137	82	138
rect	81	140	82	141
rect	81	147	82	148
rect	81	150	82	151
rect	81	153	82	154
rect	81	156	82	157
rect	81	160	82	161
rect	81	163	82	164
rect	81	166	82	167
rect	81	169	82	170
rect	81	178	82	179
rect	81	208	82	209
rect	82	1	83	2
rect	82	7	83	8
rect	82	10	83	11
rect	82	13	83	14
rect	82	16	83	17
rect	82	17	83	18
rect	82	19	83	20
rect	82	20	83	21
rect	82	22	83	23
rect	82	23	83	24
rect	82	25	83	26
rect	82	26	83	27
rect	82	34	83	35
rect	82	35	83	36
rect	82	39	83	40
rect	82	45	83	46
rect	82	49	83	50
rect	82	52	83	53
rect	82	53	83	54
rect	82	54	83	55
rect	82	55	83	56
rect	82	58	83	59
rect	82	59	83	60
rect	82	68	83	69
rect	82	71	83	72
rect	82	72	83	73
rect	82	73	83	74
rect	82	74	83	75
rect	82	75	83	76
rect	82	77	83	78
rect	82	80	83	81
rect	82	81	83	82
rect	82	83	83	84
rect	82	84	83	85
rect	82	93	83	94
rect	82	97	83	98
rect	82	103	83	104
rect	82	106	83	107
rect	82	109	83	110
rect	82	112	83	113
rect	82	115	83	116
rect	82	121	83	122
rect	82	125	83	126
rect	82	134	83	135
rect	82	137	83	138
rect	82	140	83	141
rect	82	147	83	148
rect	82	150	83	151
rect	82	153	83	154
rect	82	156	83	157
rect	82	160	83	161
rect	82	163	83	164
rect	82	166	83	167
rect	82	169	83	170
rect	82	178	83	179
rect	82	208	83	209
rect	83	1	84	2
rect	83	7	84	8
rect	83	10	84	11
rect	83	13	84	14
rect	83	16	84	17
rect	83	17	84	18
rect	83	19	84	20
rect	83	20	84	21
rect	83	22	84	23
rect	83	23	84	24
rect	83	25	84	26
rect	83	26	84	27
rect	83	34	84	35
rect	83	35	84	36
rect	83	45	84	46
rect	83	52	84	53
rect	83	53	84	54
rect	83	54	84	55
rect	83	55	84	56
rect	83	59	84	60
rect	83	68	84	69
rect	83	71	84	72
rect	83	72	84	73
rect	83	73	84	74
rect	83	74	84	75
rect	83	75	84	76
rect	83	77	84	78
rect	83	80	84	81
rect	83	81	84	82
rect	83	83	84	84
rect	83	84	84	85
rect	83	93	84	94
rect	83	97	84	98
rect	83	103	84	104
rect	83	106	84	107
rect	83	109	84	110
rect	83	112	84	113
rect	83	115	84	116
rect	83	125	84	126
rect	83	134	84	135
rect	83	137	84	138
rect	83	140	84	141
rect	83	147	84	148
rect	83	150	84	151
rect	83	153	84	154
rect	83	156	84	157
rect	83	160	84	161
rect	83	166	84	167
rect	83	169	84	170
rect	83	178	84	179
rect	83	208	84	209
rect	84	1	85	2
rect	84	7	85	8
rect	84	10	85	11
rect	84	13	85	14
rect	84	16	85	17
rect	84	17	85	18
rect	84	19	85	20
rect	84	20	85	21
rect	84	22	85	23
rect	84	23	85	24
rect	84	25	85	26
rect	84	26	85	27
rect	84	29	85	30
rect	84	34	85	35
rect	84	35	85	36
rect	84	45	85	46
rect	84	52	85	53
rect	84	53	85	54
rect	84	54	85	55
rect	84	55	85	56
rect	84	58	85	59
rect	84	59	85	60
rect	84	68	85	69
rect	84	71	85	72
rect	84	72	85	73
rect	84	73	85	74
rect	84	74	85	75
rect	84	75	85	76
rect	84	77	85	78
rect	84	80	85	81
rect	84	81	85	82
rect	84	83	85	84
rect	84	84	85	85
rect	84	93	85	94
rect	84	97	85	98
rect	84	100	85	101
rect	84	103	85	104
rect	84	106	85	107
rect	84	109	85	110
rect	84	112	85	113
rect	84	115	85	116
rect	84	125	85	126
rect	84	128	85	129
rect	84	134	85	135
rect	84	137	85	138
rect	84	140	85	141
rect	84	147	85	148
rect	84	150	85	151
rect	84	153	85	154
rect	84	156	85	157
rect	84	160	85	161
rect	84	166	85	167
rect	84	169	85	170
rect	84	172	85	173
rect	84	178	85	179
rect	84	208	85	209
rect	85	7	86	8
rect	85	16	86	17
rect	85	17	86	18
rect	85	19	86	20
rect	85	20	86	21
rect	85	22	86	23
rect	85	23	86	24
rect	85	25	86	26
rect	85	29	86	30
rect	85	34	86	35
rect	85	35	86	36
rect	85	52	86	53
rect	85	53	86	54
rect	85	54	86	55
rect	85	58	86	59
rect	85	59	86	60
rect	85	68	86	69
rect	85	71	86	72
rect	85	72	86	73
rect	85	73	86	74
rect	85	74	86	75
rect	85	75	86	76
rect	85	77	86	78
rect	85	80	86	81
rect	85	81	86	82
rect	85	83	86	84
rect	85	84	86	85
rect	85	93	86	94
rect	85	97	86	98
rect	85	100	86	101
rect	85	103	86	104
rect	85	106	86	107
rect	85	109	86	110
rect	85	112	86	113
rect	85	115	86	116
rect	85	125	86	126
rect	85	128	86	129
rect	85	134	86	135
rect	85	137	86	138
rect	85	140	86	141
rect	85	147	86	148
rect	85	150	86	151
rect	85	153	86	154
rect	85	156	86	157
rect	85	160	86	161
rect	85	166	86	167
rect	85	169	86	170
rect	85	172	86	173
rect	85	178	86	179
rect	85	208	86	209
rect	86	7	87	8
rect	86	16	87	17
rect	86	17	87	18
rect	86	19	87	20
rect	86	20	87	21
rect	86	22	87	23
rect	86	23	87	24
rect	86	25	87	26
rect	86	26	87	27
rect	86	29	87	30
rect	86	34	87	35
rect	86	35	87	36
rect	86	36	87	37
rect	86	39	87	40
rect	86	42	87	43
rect	86	52	87	53
rect	86	53	87	54
rect	86	54	87	55
rect	86	58	87	59
rect	86	59	87	60
rect	86	62	87	63
rect	86	65	87	66
rect	86	68	87	69
rect	86	71	87	72
rect	86	72	87	73
rect	86	73	87	74
rect	86	74	87	75
rect	86	75	87	76
rect	86	77	87	78
rect	86	80	87	81
rect	86	81	87	82
rect	86	83	87	84
rect	86	84	87	85
rect	86	93	87	94
rect	86	97	87	98
rect	86	100	87	101
rect	86	103	87	104
rect	86	106	87	107
rect	86	109	87	110
rect	86	112	87	113
rect	86	115	87	116
rect	86	125	87	126
rect	86	128	87	129
rect	86	134	87	135
rect	86	137	87	138
rect	86	140	87	141
rect	86	147	87	148
rect	86	150	87	151
rect	86	153	87	154
rect	86	156	87	157
rect	86	160	87	161
rect	86	163	87	164
rect	86	166	87	167
rect	86	169	87	170
rect	86	172	87	173
rect	86	178	87	179
rect	86	208	87	209
rect	87	16	88	17
rect	87	17	88	18
rect	87	19	88	20
rect	87	20	88	21
rect	87	22	88	23
rect	87	23	88	24
rect	87	25	88	26
rect	87	26	88	27
rect	87	29	88	30
rect	87	34	88	35
rect	87	35	88	36
rect	87	36	88	37
rect	87	39	88	40
rect	87	42	88	43
rect	87	52	88	53
rect	87	53	88	54
rect	87	54	88	55
rect	87	58	88	59
rect	87	59	88	60
rect	87	62	88	63
rect	87	65	88	66
rect	87	68	88	69
rect	87	71	88	72
rect	87	72	88	73
rect	87	73	88	74
rect	87	74	88	75
rect	87	75	88	76
rect	87	77	88	78
rect	87	80	88	81
rect	87	81	88	82
rect	87	83	88	84
rect	87	84	88	85
rect	87	93	88	94
rect	87	97	88	98
rect	87	100	88	101
rect	87	103	88	104
rect	87	106	88	107
rect	87	109	88	110
rect	87	112	88	113
rect	87	115	88	116
rect	87	125	88	126
rect	87	128	88	129
rect	87	134	88	135
rect	87	137	88	138
rect	87	140	88	141
rect	87	147	88	148
rect	87	150	88	151
rect	87	153	88	154
rect	87	156	88	157
rect	87	163	88	164
rect	87	166	88	167
rect	87	169	88	170
rect	87	172	88	173
rect	87	178	88	179
rect	87	208	88	209
rect	88	4	89	5
rect	88	11	89	12
rect	88	14	89	15
rect	88	16	89	17
rect	88	17	89	18
rect	88	19	89	20
rect	88	20	89	21
rect	88	22	89	23
rect	88	23	89	24
rect	88	25	89	26
rect	88	26	89	27
rect	88	29	89	30
rect	88	33	89	34
rect	88	34	89	35
rect	88	35	89	36
rect	88	36	89	37
rect	88	39	89	40
rect	88	42	89	43
rect	88	52	89	53
rect	88	53	89	54
rect	88	54	89	55
rect	88	58	89	59
rect	88	59	89	60
rect	88	62	89	63
rect	88	65	89	66
rect	88	68	89	69
rect	88	71	89	72
rect	88	72	89	73
rect	88	73	89	74
rect	88	74	89	75
rect	88	75	89	76
rect	88	77	89	78
rect	88	80	89	81
rect	88	81	89	82
rect	88	83	89	84
rect	88	84	89	85
rect	88	93	89	94
rect	88	97	89	98
rect	88	100	89	101
rect	88	103	89	104
rect	88	106	89	107
rect	88	109	89	110
rect	88	112	89	113
rect	88	115	89	116
rect	88	125	89	126
rect	88	128	89	129
rect	88	131	89	132
rect	88	134	89	135
rect	88	137	89	138
rect	88	140	89	141
rect	88	147	89	148
rect	88	150	89	151
rect	88	153	89	154
rect	88	156	89	157
rect	88	163	89	164
rect	88	166	89	167
rect	88	169	89	170
rect	88	172	89	173
rect	88	175	89	176
rect	88	178	89	179
rect	88	208	89	209
rect	89	16	90	17
rect	89	17	90	18
rect	89	19	90	20
rect	89	20	90	21
rect	89	22	90	23
rect	89	23	90	24
rect	89	25	90	26
rect	89	26	90	27
rect	89	34	90	35
rect	89	35	90	36
rect	89	53	90	54
rect	89	54	90	55
rect	89	58	90	59
rect	89	59	90	60
rect	89	72	90	73
rect	89	73	90	74
rect	89	74	90	75
rect	89	75	90	76
rect	89	80	90	81
rect	89	81	90	82
rect	89	83	90	84
rect	89	84	90	85
rect	90	16	91	17
rect	90	17	91	18
rect	90	19	91	20
rect	90	20	91	21
rect	90	22	91	23
rect	90	23	91	24
rect	90	25	91	26
rect	90	26	91	27
rect	90	34	91	35
rect	90	35	91	36
rect	90	53	91	54
rect	90	54	91	55
rect	90	58	91	59
rect	90	59	91	60
rect	90	72	91	73
rect	90	73	91	74
rect	90	74	91	75
rect	90	75	91	76
rect	90	80	91	81
rect	90	81	91	82
rect	90	83	91	84
rect	90	84	91	85
rect	91	16	92	17
rect	91	17	92	18
rect	91	19	92	20
rect	91	20	92	21
rect	91	22	92	23
rect	91	23	92	24
rect	91	25	92	26
rect	91	26	92	27
rect	91	34	92	35
rect	91	35	92	36
rect	91	53	92	54
rect	91	54	92	55
rect	91	58	92	59
rect	91	59	92	60
rect	91	72	92	73
rect	91	73	92	74
rect	91	74	92	75
rect	91	75	92	76
rect	91	80	92	81
rect	91	81	92	82
rect	91	83	92	84
rect	91	84	92	85
rect	92	16	93	17
rect	92	17	93	18
rect	92	19	93	20
rect	92	20	93	21
rect	92	22	93	23
rect	92	23	93	24
rect	92	25	93	26
rect	92	26	93	27
rect	92	34	93	35
rect	92	35	93	36
rect	92	53	93	54
rect	92	54	93	55
rect	92	58	93	59
rect	92	59	93	60
rect	92	72	93	73
rect	92	73	93	74
rect	92	74	93	75
rect	92	75	93	76
rect	92	80	93	81
rect	92	81	93	82
rect	92	83	93	84
rect	92	84	93	85
rect	93	16	94	17
rect	93	17	94	18
rect	93	19	94	20
rect	93	20	94	21
rect	93	22	94	23
rect	93	23	94	24
rect	93	25	94	26
rect	93	26	94	27
rect	93	34	94	35
rect	93	35	94	36
rect	93	53	94	54
rect	93	54	94	55
rect	93	58	94	59
rect	93	59	94	60
rect	93	72	94	73
rect	93	73	94	74
rect	93	74	94	75
rect	93	75	94	76
rect	93	80	94	81
rect	93	81	94	82
rect	93	83	94	84
rect	93	84	94	85
rect	94	16	95	17
rect	94	17	95	18
rect	94	19	95	20
rect	94	20	95	21
rect	94	22	95	23
rect	94	23	95	24
rect	94	25	95	26
rect	94	26	95	27
rect	94	34	95	35
rect	94	35	95	36
rect	94	53	95	54
rect	94	54	95	55
rect	94	58	95	59
rect	94	59	95	60
rect	94	72	95	73
rect	94	73	95	74
rect	94	75	95	76
rect	94	81	95	82
rect	94	83	95	84
rect	94	84	95	85
rect	95	1	96	2
rect	95	11	96	12
rect	95	14	96	15
rect	95	16	96	17
rect	95	17	96	18
rect	95	19	96	20
rect	95	20	96	21
rect	95	22	96	23
rect	95	23	96	24
rect	95	25	96	26
rect	95	26	96	27
rect	95	29	96	30
rect	95	33	96	34
rect	95	34	96	35
rect	95	35	96	36
rect	95	39	96	40
rect	95	42	96	43
rect	95	52	96	53
rect	95	53	96	54
rect	95	54	96	55
rect	95	58	96	59
rect	95	59	96	60
rect	95	62	96	63
rect	95	65	96	66
rect	95	68	96	69
rect	95	71	96	72
rect	95	72	96	73
rect	95	73	96	74
rect	95	75	96	76
rect	95	77	96	78
rect	95	81	96	82
rect	95	83	96	84
rect	95	84	96	85
rect	95	87	96	88
rect	95	90	96	91
rect	95	93	96	94
rect	95	97	96	98
rect	95	100	96	101
rect	95	103	96	104
rect	95	106	96	107
rect	95	109	96	110
rect	95	112	96	113
rect	95	115	96	116
rect	95	119	96	120
rect	95	122	96	123
rect	95	125	96	126
rect	95	128	96	129
rect	95	131	96	132
rect	95	134	96	135
rect	95	137	96	138
rect	95	140	96	141
rect	95	144	96	145
rect	95	147	96	148
rect	95	150	96	151
rect	95	153	96	154
rect	95	156	96	157
rect	95	160	96	161
rect	95	166	96	167
rect	95	169	96	170
rect	95	172	96	173
rect	95	175	96	176
rect	95	178	96	179
rect	95	208	96	209
rect	96	1	97	2
rect	96	11	97	12
rect	96	14	97	15
rect	96	16	97	17
rect	96	17	97	18
rect	96	19	97	20
rect	96	20	97	21
rect	96	22	97	23
rect	96	23	97	24
rect	96	25	97	26
rect	96	26	97	27
rect	96	29	97	30
rect	96	33	97	34
rect	96	34	97	35
rect	96	35	97	36
rect	96	39	97	40
rect	96	42	97	43
rect	96	52	97	53
rect	96	53	97	54
rect	96	54	97	55
rect	96	58	97	59
rect	96	59	97	60
rect	96	62	97	63
rect	96	65	97	66
rect	96	68	97	69
rect	96	71	97	72
rect	96	72	97	73
rect	96	73	97	74
rect	96	75	97	76
rect	96	77	97	78
rect	96	81	97	82
rect	96	83	97	84
rect	96	84	97	85
rect	96	87	97	88
rect	96	90	97	91
rect	96	93	97	94
rect	96	97	97	98
rect	96	100	97	101
rect	96	103	97	104
rect	96	106	97	107
rect	96	109	97	110
rect	96	112	97	113
rect	96	115	97	116
rect	96	119	97	120
rect	96	122	97	123
rect	96	125	97	126
rect	96	128	97	129
rect	96	131	97	132
rect	96	134	97	135
rect	96	137	97	138
rect	96	140	97	141
rect	96	144	97	145
rect	96	147	97	148
rect	96	150	97	151
rect	96	153	97	154
rect	96	156	97	157
rect	96	160	97	161
rect	96	166	97	167
rect	96	169	97	170
rect	96	172	97	173
rect	96	175	97	176
rect	96	178	97	179
rect	96	208	97	209
rect	97	1	98	2
rect	97	11	98	12
rect	97	14	98	15
rect	97	16	98	17
rect	97	17	98	18
rect	97	19	98	20
rect	97	20	98	21
rect	97	22	98	23
rect	97	23	98	24
rect	97	25	98	26
rect	97	26	98	27
rect	97	29	98	30
rect	97	33	98	34
rect	97	34	98	35
rect	97	35	98	36
rect	97	39	98	40
rect	97	42	98	43
rect	97	52	98	53
rect	97	53	98	54
rect	97	54	98	55
rect	97	58	98	59
rect	97	59	98	60
rect	97	62	98	63
rect	97	65	98	66
rect	97	68	98	69
rect	97	71	98	72
rect	97	72	98	73
rect	97	73	98	74
rect	97	75	98	76
rect	97	77	98	78
rect	97	81	98	82
rect	97	83	98	84
rect	97	84	98	85
rect	97	87	98	88
rect	97	90	98	91
rect	97	93	98	94
rect	97	97	98	98
rect	97	100	98	101
rect	97	103	98	104
rect	97	106	98	107
rect	97	109	98	110
rect	97	112	98	113
rect	97	115	98	116
rect	97	119	98	120
rect	97	122	98	123
rect	97	125	98	126
rect	97	128	98	129
rect	97	131	98	132
rect	97	134	98	135
rect	97	137	98	138
rect	97	140	98	141
rect	97	144	98	145
rect	97	147	98	148
rect	97	150	98	151
rect	97	153	98	154
rect	97	156	98	157
rect	97	160	98	161
rect	97	166	98	167
rect	97	169	98	170
rect	97	172	98	173
rect	97	175	98	176
rect	97	178	98	179
rect	97	208	98	209
rect	98	1	99	2
rect	98	11	99	12
rect	98	14	99	15
rect	98	16	99	17
rect	98	17	99	18
rect	98	19	99	20
rect	98	20	99	21
rect	98	22	99	23
rect	98	23	99	24
rect	98	25	99	26
rect	98	26	99	27
rect	98	29	99	30
rect	98	33	99	34
rect	98	34	99	35
rect	98	35	99	36
rect	98	39	99	40
rect	98	42	99	43
rect	98	52	99	53
rect	98	53	99	54
rect	98	54	99	55
rect	98	58	99	59
rect	98	59	99	60
rect	98	62	99	63
rect	98	65	99	66
rect	98	68	99	69
rect	98	71	99	72
rect	98	72	99	73
rect	98	73	99	74
rect	98	75	99	76
rect	98	77	99	78
rect	98	81	99	82
rect	98	83	99	84
rect	98	84	99	85
rect	98	87	99	88
rect	98	90	99	91
rect	98	93	99	94
rect	98	97	99	98
rect	98	100	99	101
rect	98	103	99	104
rect	98	106	99	107
rect	98	109	99	110
rect	98	112	99	113
rect	98	115	99	116
rect	98	119	99	120
rect	98	122	99	123
rect	98	125	99	126
rect	98	128	99	129
rect	98	131	99	132
rect	98	134	99	135
rect	98	137	99	138
rect	98	140	99	141
rect	98	144	99	145
rect	98	147	99	148
rect	98	150	99	151
rect	98	153	99	154
rect	98	156	99	157
rect	98	160	99	161
rect	98	166	99	167
rect	98	169	99	170
rect	98	172	99	173
rect	98	175	99	176
rect	98	178	99	179
rect	98	208	99	209
rect	99	1	100	2
rect	99	11	100	12
rect	99	14	100	15
rect	99	16	100	17
rect	99	17	100	18
rect	99	19	100	20
rect	99	20	100	21
rect	99	22	100	23
rect	99	23	100	24
rect	99	25	100	26
rect	99	26	100	27
rect	99	29	100	30
rect	99	33	100	34
rect	99	34	100	35
rect	99	35	100	36
rect	99	39	100	40
rect	99	42	100	43
rect	99	52	100	53
rect	99	53	100	54
rect	99	54	100	55
rect	99	58	100	59
rect	99	59	100	60
rect	99	62	100	63
rect	99	65	100	66
rect	99	68	100	69
rect	99	71	100	72
rect	99	72	100	73
rect	99	73	100	74
rect	99	75	100	76
rect	99	77	100	78
rect	99	81	100	82
rect	99	83	100	84
rect	99	84	100	85
rect	99	87	100	88
rect	99	90	100	91
rect	99	93	100	94
rect	99	97	100	98
rect	99	100	100	101
rect	99	103	100	104
rect	99	106	100	107
rect	99	109	100	110
rect	99	112	100	113
rect	99	115	100	116
rect	99	119	100	120
rect	99	122	100	123
rect	99	125	100	126
rect	99	128	100	129
rect	99	131	100	132
rect	99	134	100	135
rect	99	137	100	138
rect	99	140	100	141
rect	99	144	100	145
rect	99	147	100	148
rect	99	150	100	151
rect	99	153	100	154
rect	99	156	100	157
rect	99	160	100	161
rect	99	166	100	167
rect	99	169	100	170
rect	99	172	100	173
rect	99	175	100	176
rect	99	178	100	179
rect	99	208	100	209
rect	100	1	101	2
rect	100	11	101	12
rect	100	14	101	15
rect	100	16	101	17
rect	100	17	101	18
rect	100	19	101	20
rect	100	20	101	21
rect	100	22	101	23
rect	100	23	101	24
rect	100	25	101	26
rect	100	26	101	27
rect	100	29	101	30
rect	100	33	101	34
rect	100	34	101	35
rect	100	35	101	36
rect	100	39	101	40
rect	100	42	101	43
rect	100	52	101	53
rect	100	53	101	54
rect	100	54	101	55
rect	100	58	101	59
rect	100	59	101	60
rect	100	62	101	63
rect	100	65	101	66
rect	100	68	101	69
rect	100	71	101	72
rect	100	72	101	73
rect	100	73	101	74
rect	100	75	101	76
rect	100	77	101	78
rect	100	81	101	82
rect	100	83	101	84
rect	100	84	101	85
rect	100	87	101	88
rect	100	90	101	91
rect	100	93	101	94
rect	100	97	101	98
rect	100	100	101	101
rect	100	103	101	104
rect	100	106	101	107
rect	100	109	101	110
rect	100	112	101	113
rect	100	115	101	116
rect	100	119	101	120
rect	100	122	101	123
rect	100	125	101	126
rect	100	128	101	129
rect	100	131	101	132
rect	100	134	101	135
rect	100	137	101	138
rect	100	140	101	141
rect	100	144	101	145
rect	100	147	101	148
rect	100	150	101	151
rect	100	153	101	154
rect	100	156	101	157
rect	100	160	101	161
rect	100	166	101	167
rect	100	169	101	170
rect	100	172	101	173
rect	100	175	101	176
rect	100	178	101	179
rect	100	208	101	209
rect	101	1	102	2
rect	101	11	102	12
rect	101	14	102	15
rect	101	16	102	17
rect	101	17	102	18
rect	101	19	102	20
rect	101	20	102	21
rect	101	22	102	23
rect	101	23	102	24
rect	101	25	102	26
rect	101	26	102	27
rect	101	29	102	30
rect	101	33	102	34
rect	101	34	102	35
rect	101	35	102	36
rect	101	39	102	40
rect	101	42	102	43
rect	101	52	102	53
rect	101	53	102	54
rect	101	54	102	55
rect	101	58	102	59
rect	101	59	102	60
rect	101	62	102	63
rect	101	65	102	66
rect	101	68	102	69
rect	101	71	102	72
rect	101	72	102	73
rect	101	73	102	74
rect	101	75	102	76
rect	101	77	102	78
rect	101	81	102	82
rect	101	83	102	84
rect	101	84	102	85
rect	101	87	102	88
rect	101	90	102	91
rect	101	93	102	94
rect	101	97	102	98
rect	101	100	102	101
rect	101	103	102	104
rect	101	106	102	107
rect	101	109	102	110
rect	101	112	102	113
rect	101	115	102	116
rect	101	119	102	120
rect	101	122	102	123
rect	101	125	102	126
rect	101	128	102	129
rect	101	131	102	132
rect	101	134	102	135
rect	101	137	102	138
rect	101	140	102	141
rect	101	144	102	145
rect	101	147	102	148
rect	101	150	102	151
rect	101	153	102	154
rect	101	156	102	157
rect	101	160	102	161
rect	101	166	102	167
rect	101	169	102	170
rect	101	172	102	173
rect	101	175	102	176
rect	101	178	102	179
rect	101	208	102	209
rect	102	1	103	2
rect	102	11	103	12
rect	102	14	103	15
rect	102	16	103	17
rect	102	17	103	18
rect	102	19	103	20
rect	102	20	103	21
rect	102	22	103	23
rect	102	23	103	24
rect	102	25	103	26
rect	102	26	103	27
rect	102	29	103	30
rect	102	33	103	34
rect	102	34	103	35
rect	102	35	103	36
rect	102	42	103	43
rect	102	52	103	53
rect	102	53	103	54
rect	102	54	103	55
rect	102	58	103	59
rect	102	59	103	60
rect	102	62	103	63
rect	102	65	103	66
rect	102	68	103	69
rect	102	71	103	72
rect	102	72	103	73
rect	102	73	103	74
rect	102	75	103	76
rect	102	77	103	78
rect	102	81	103	82
rect	102	83	103	84
rect	102	84	103	85
rect	102	87	103	88
rect	102	90	103	91
rect	102	93	103	94
rect	102	97	103	98
rect	102	103	103	104
rect	102	106	103	107
rect	102	109	103	110
rect	102	112	103	113
rect	102	115	103	116
rect	102	119	103	120
rect	102	125	103	126
rect	102	131	103	132
rect	102	134	103	135
rect	102	137	103	138
rect	102	140	103	141
rect	102	144	103	145
rect	102	147	103	148
rect	102	150	103	151
rect	102	153	103	154
rect	102	156	103	157
rect	102	160	103	161
rect	102	166	103	167
rect	102	169	103	170
rect	102	172	103	173
rect	102	175	103	176
rect	102	178	103	179
rect	102	208	103	209
rect	103	1	104	2
rect	103	11	104	12
rect	103	14	104	15
rect	103	16	104	17
rect	103	17	104	18
rect	103	19	104	20
rect	103	20	104	21
rect	103	22	104	23
rect	103	23	104	24
rect	103	25	104	26
rect	103	26	104	27
rect	103	29	104	30
rect	103	33	104	34
rect	103	34	104	35
rect	103	35	104	36
rect	103	42	104	43
rect	103	52	104	53
rect	103	53	104	54
rect	103	54	104	55
rect	103	58	104	59
rect	103	59	104	60
rect	103	62	104	63
rect	103	65	104	66
rect	103	68	104	69
rect	103	71	104	72
rect	103	72	104	73
rect	103	73	104	74
rect	103	75	104	76
rect	103	77	104	78
rect	103	81	104	82
rect	103	83	104	84
rect	103	84	104	85
rect	103	87	104	88
rect	103	90	104	91
rect	103	93	104	94
rect	103	97	104	98
rect	103	103	104	104
rect	103	106	104	107
rect	103	109	104	110
rect	103	112	104	113
rect	103	115	104	116
rect	103	119	104	120
rect	103	125	104	126
rect	103	131	104	132
rect	103	134	104	135
rect	103	137	104	138
rect	103	140	104	141
rect	103	144	104	145
rect	103	147	104	148
rect	103	150	104	151
rect	103	153	104	154
rect	103	156	104	157
rect	103	160	104	161
rect	103	166	104	167
rect	103	169	104	170
rect	103	172	104	173
rect	103	175	104	176
rect	103	178	104	179
rect	103	208	104	209
rect	104	1	105	2
rect	104	11	105	12
rect	104	14	105	15
rect	104	16	105	17
rect	104	17	105	18
rect	104	19	105	20
rect	104	20	105	21
rect	104	22	105	23
rect	104	23	105	24
rect	104	25	105	26
rect	104	26	105	27
rect	104	29	105	30
rect	104	33	105	34
rect	104	34	105	35
rect	104	35	105	36
rect	104	42	105	43
rect	104	52	105	53
rect	104	53	105	54
rect	104	54	105	55
rect	104	58	105	59
rect	104	59	105	60
rect	104	62	105	63
rect	104	65	105	66
rect	104	68	105	69
rect	104	71	105	72
rect	104	72	105	73
rect	104	73	105	74
rect	104	75	105	76
rect	104	77	105	78
rect	104	81	105	82
rect	104	83	105	84
rect	104	84	105	85
rect	104	93	105	94
rect	104	97	105	98
rect	104	103	105	104
rect	104	106	105	107
rect	104	112	105	113
rect	104	115	105	116
rect	104	119	105	120
rect	104	125	105	126
rect	104	131	105	132
rect	104	134	105	135
rect	104	137	105	138
rect	104	140	105	141
rect	104	144	105	145
rect	104	147	105	148
rect	104	150	105	151
rect	104	153	105	154
rect	104	156	105	157
rect	104	160	105	161
rect	104	166	105	167
rect	104	169	105	170
rect	104	172	105	173
rect	104	175	105	176
rect	104	178	105	179
rect	104	208	105	209
rect	105	1	106	2
rect	105	11	106	12
rect	105	14	106	15
rect	105	16	106	17
rect	105	17	106	18
rect	105	19	106	20
rect	105	20	106	21
rect	105	22	106	23
rect	105	23	106	24
rect	105	25	106	26
rect	105	26	106	27
rect	105	29	106	30
rect	105	33	106	34
rect	105	34	106	35
rect	105	35	106	36
rect	105	38	106	39
rect	105	42	106	43
rect	105	52	106	53
rect	105	53	106	54
rect	105	54	106	55
rect	105	58	106	59
rect	105	59	106	60
rect	105	62	106	63
rect	105	65	106	66
rect	105	68	106	69
rect	105	71	106	72
rect	105	72	106	73
rect	105	73	106	74
rect	105	75	106	76
rect	105	77	106	78
rect	105	81	106	82
rect	105	83	106	84
rect	105	84	106	85
rect	105	93	106	94
rect	105	97	106	98
rect	105	100	106	101
rect	105	103	106	104
rect	105	106	106	107
rect	105	112	106	113
rect	105	115	106	116
rect	105	119	106	120
rect	105	125	106	126
rect	105	129	106	130
rect	105	131	106	132
rect	105	134	106	135
rect	105	137	106	138
rect	105	140	106	141
rect	105	144	106	145
rect	105	147	106	148
rect	105	150	106	151
rect	105	153	106	154
rect	105	156	106	157
rect	105	160	106	161
rect	105	166	106	167
rect	105	169	106	170
rect	105	172	106	173
rect	105	175	106	176
rect	105	178	106	179
rect	105	208	106	209
rect	106	1	107	2
rect	106	11	107	12
rect	106	14	107	15
rect	106	16	107	17
rect	106	17	107	18
rect	106	19	107	20
rect	106	20	107	21
rect	106	22	107	23
rect	106	23	107	24
rect	106	25	107	26
rect	106	26	107	27
rect	106	29	107	30
rect	106	33	107	34
rect	106	34	107	35
rect	106	35	107	36
rect	106	38	107	39
rect	106	42	107	43
rect	106	52	107	53
rect	106	53	107	54
rect	106	54	107	55
rect	106	58	107	59
rect	106	59	107	60
rect	106	62	107	63
rect	106	71	107	72
rect	106	72	107	73
rect	106	73	107	74
rect	106	75	107	76
rect	106	77	107	78
rect	106	81	107	82
rect	106	83	107	84
rect	106	84	107	85
rect	106	93	107	94
rect	106	97	107	98
rect	106	100	107	101
rect	106	103	107	104
rect	106	106	107	107
rect	106	112	107	113
rect	106	115	107	116
rect	106	119	107	120
rect	106	129	107	130
rect	106	131	107	132
rect	106	134	107	135
rect	106	137	107	138
rect	106	140	107	141
rect	106	144	107	145
rect	106	147	107	148
rect	106	150	107	151
rect	106	153	107	154
rect	106	156	107	157
rect	106	160	107	161
rect	106	166	107	167
rect	106	169	107	170
rect	106	172	107	173
rect	106	175	107	176
rect	106	178	107	179
rect	106	208	107	209
rect	107	1	108	2
rect	107	11	108	12
rect	107	14	108	15
rect	107	16	108	17
rect	107	17	108	18
rect	107	19	108	20
rect	107	20	108	21
rect	107	22	108	23
rect	107	23	108	24
rect	107	25	108	26
rect	107	26	108	27
rect	107	29	108	30
rect	107	33	108	34
rect	107	34	108	35
rect	107	35	108	36
rect	107	38	108	39
rect	107	42	108	43
rect	107	47	108	48
rect	107	52	108	53
rect	107	53	108	54
rect	107	54	108	55
rect	107	58	108	59
rect	107	59	108	60
rect	107	62	108	63
rect	107	71	108	72
rect	107	72	108	73
rect	107	73	108	74
rect	107	75	108	76
rect	107	77	108	78
rect	107	81	108	82
rect	107	83	108	84
rect	107	84	108	85
rect	107	88	108	89
rect	107	93	108	94
rect	107	97	108	98
rect	107	100	108	101
rect	107	103	108	104
rect	107	106	108	107
rect	107	110	108	111
rect	107	112	108	113
rect	107	115	108	116
rect	107	119	108	120
rect	107	129	108	130
rect	107	131	108	132
rect	107	134	108	135
rect	107	137	108	138
rect	107	140	108	141
rect	107	144	108	145
rect	107	147	108	148
rect	107	150	108	151
rect	107	153	108	154
rect	107	156	108	157
rect	107	160	108	161
rect	107	166	108	167
rect	107	169	108	170
rect	107	172	108	173
rect	107	175	108	176
rect	107	178	108	179
rect	107	208	108	209
rect	108	1	109	2
rect	108	11	109	12
rect	108	14	109	15
rect	108	16	109	17
rect	108	17	109	18
rect	108	19	109	20
rect	108	20	109	21
rect	108	22	109	23
rect	108	23	109	24
rect	108	25	109	26
rect	108	26	109	27
rect	108	29	109	30
rect	108	33	109	34
rect	108	34	109	35
rect	108	35	109	36
rect	108	38	109	39
rect	108	42	109	43
rect	108	47	109	48
rect	108	52	109	53
rect	108	53	109	54
rect	108	54	109	55
rect	108	58	109	59
rect	108	59	109	60
rect	108	62	109	63
rect	108	71	109	72
rect	108	72	109	73
rect	108	73	109	74
rect	108	75	109	76
rect	108	77	109	78
rect	108	81	109	82
rect	108	83	109	84
rect	108	84	109	85
rect	108	88	109	89
rect	108	97	109	98
rect	108	100	109	101
rect	108	103	109	104
rect	108	106	109	107
rect	108	110	109	111
rect	108	112	109	113
rect	108	115	109	116
rect	108	119	109	120
rect	108	129	109	130
rect	108	134	109	135
rect	108	137	109	138
rect	108	140	109	141
rect	108	144	109	145
rect	108	153	109	154
rect	108	156	109	157
rect	108	160	109	161
rect	108	166	109	167
rect	108	169	109	170
rect	108	172	109	173
rect	108	175	109	176
rect	108	178	109	179
rect	108	208	109	209
rect	109	1	110	2
rect	109	11	110	12
rect	109	14	110	15
rect	109	16	110	17
rect	109	17	110	18
rect	109	19	110	20
rect	109	20	110	21
rect	109	22	110	23
rect	109	23	110	24
rect	109	25	110	26
rect	109	26	110	27
rect	109	29	110	30
rect	109	33	110	34
rect	109	34	110	35
rect	109	35	110	36
rect	109	38	110	39
rect	109	42	110	43
rect	109	47	110	48
rect	109	52	110	53
rect	109	53	110	54
rect	109	54	110	55
rect	109	58	110	59
rect	109	59	110	60
rect	109	62	110	63
rect	109	66	110	67
rect	109	71	110	72
rect	109	72	110	73
rect	109	73	110	74
rect	109	75	110	76
rect	109	77	110	78
rect	109	81	110	82
rect	109	83	110	84
rect	109	84	110	85
rect	109	88	110	89
rect	109	97	110	98
rect	109	100	110	101
rect	109	103	110	104
rect	109	106	110	107
rect	109	110	110	111
rect	109	112	110	113
rect	109	115	110	116
rect	109	119	110	120
rect	109	126	110	127
rect	109	129	110	130
rect	109	134	110	135
rect	109	137	110	138
rect	109	140	110	141
rect	109	144	110	145
rect	109	153	110	154
rect	109	156	110	157
rect	109	160	110	161
rect	109	166	110	167
rect	109	169	110	170
rect	109	172	110	173
rect	109	175	110	176
rect	109	178	110	179
rect	109	208	110	209
rect	110	1	111	2
rect	110	11	111	12
rect	110	14	111	15
rect	110	16	111	17
rect	110	17	111	18
rect	110	19	111	20
rect	110	20	111	21
rect	110	22	111	23
rect	110	23	111	24
rect	110	25	111	26
rect	110	26	111	27
rect	110	29	111	30
rect	110	33	111	34
rect	110	34	111	35
rect	110	35	111	36
rect	110	38	111	39
rect	110	42	111	43
rect	110	47	111	48
rect	110	52	111	53
rect	110	53	111	54
rect	110	54	111	55
rect	110	58	111	59
rect	110	59	111	60
rect	110	66	111	67
rect	110	71	111	72
rect	110	72	111	73
rect	110	73	111	74
rect	110	75	111	76
rect	110	77	111	78
rect	110	81	111	82
rect	110	83	111	84
rect	110	84	111	85
rect	110	88	111	89
rect	110	97	111	98
rect	110	100	111	101
rect	110	103	111	104
rect	110	106	111	107
rect	110	110	111	111
rect	110	112	111	113
rect	110	115	111	116
rect	110	119	111	120
rect	110	126	111	127
rect	110	129	111	130
rect	110	134	111	135
rect	110	137	111	138
rect	110	140	111	141
rect	110	144	111	145
rect	110	153	111	154
rect	110	156	111	157
rect	110	160	111	161
rect	110	166	111	167
rect	110	169	111	170
rect	110	172	111	173
rect	110	175	111	176
rect	110	178	111	179
rect	110	208	111	209
rect	111	1	112	2
rect	111	11	112	12
rect	111	14	112	15
rect	111	16	112	17
rect	111	17	112	18
rect	111	19	112	20
rect	111	20	112	21
rect	111	22	112	23
rect	111	23	112	24
rect	111	25	112	26
rect	111	26	112	27
rect	111	29	112	30
rect	111	33	112	34
rect	111	34	112	35
rect	111	35	112	36
rect	111	38	112	39
rect	111	42	112	43
rect	111	47	112	48
rect	111	52	112	53
rect	111	53	112	54
rect	111	54	112	55
rect	111	58	112	59
rect	111	59	112	60
rect	111	66	112	67
rect	111	71	112	72
rect	111	72	112	73
rect	111	73	112	74
rect	111	75	112	76
rect	111	77	112	78
rect	111	81	112	82
rect	111	83	112	84
rect	111	84	112	85
rect	111	88	112	89
rect	111	97	112	98
rect	111	100	112	101
rect	111	103	112	104
rect	111	106	112	107
rect	111	110	112	111
rect	111	112	112	113
rect	111	115	112	116
rect	111	119	112	120
rect	111	126	112	127
rect	111	129	112	130
rect	111	134	112	135
rect	111	137	112	138
rect	111	140	112	141
rect	111	144	112	145
rect	111	153	112	154
rect	111	156	112	157
rect	111	160	112	161
rect	111	166	112	167
rect	111	169	112	170
rect	111	172	112	173
rect	111	175	112	176
rect	111	178	112	179
rect	111	196	112	197
rect	111	208	112	209
rect	112	1	113	2
rect	112	11	113	12
rect	112	14	113	15
rect	112	16	113	17
rect	112	17	113	18
rect	112	19	113	20
rect	112	20	113	21
rect	112	22	113	23
rect	112	23	113	24
rect	112	25	113	26
rect	112	26	113	27
rect	112	29	113	30
rect	112	33	113	34
rect	112	34	113	35
rect	112	35	113	36
rect	112	38	113	39
rect	112	42	113	43
rect	112	47	113	48
rect	112	52	113	53
rect	112	53	113	54
rect	112	54	113	55
rect	112	58	113	59
rect	112	59	113	60
rect	112	66	113	67
rect	112	72	113	73
rect	112	73	113	74
rect	112	75	113	76
rect	112	81	113	82
rect	112	83	113	84
rect	112	84	113	85
rect	112	88	113	89
rect	112	100	113	101
rect	112	106	113	107
rect	112	110	113	111
rect	112	112	113	113
rect	112	115	113	116
rect	112	126	113	127
rect	112	129	113	130
rect	112	134	113	135
rect	112	137	113	138
rect	112	140	113	141
rect	112	144	113	145
rect	112	153	113	154
rect	112	160	113	161
rect	112	166	113	167
rect	112	169	113	170
rect	112	172	113	173
rect	112	175	113	176
rect	112	178	113	179
rect	112	196	113	197
rect	112	208	113	209
rect	113	1	114	2
rect	113	11	114	12
rect	113	14	114	15
rect	113	16	114	17
rect	113	17	114	18
rect	113	19	114	20
rect	113	20	114	21
rect	113	22	114	23
rect	113	23	114	24
rect	113	25	114	26
rect	113	26	114	27
rect	113	29	114	30
rect	113	31	114	32
rect	113	33	114	34
rect	113	34	114	35
rect	113	35	114	36
rect	113	38	114	39
rect	113	42	114	43
rect	113	47	114	48
rect	113	52	114	53
rect	113	53	114	54
rect	113	54	114	55
rect	113	58	114	59
rect	113	59	114	60
rect	113	60	114	61
rect	113	63	114	64
rect	113	66	114	67
rect	113	72	114	73
rect	113	73	114	74
rect	113	75	114	76
rect	113	81	114	82
rect	113	83	114	84
rect	113	84	114	85
rect	113	88	114	89
rect	113	100	114	101
rect	113	106	114	107
rect	113	110	114	111
rect	113	112	114	113
rect	113	115	114	116
rect	113	126	114	127
rect	113	129	114	130
rect	113	132	114	133
rect	113	134	114	135
rect	113	137	114	138
rect	113	140	114	141
rect	113	144	114	145
rect	113	153	114	154
rect	113	160	114	161
rect	113	166	114	167
rect	113	169	114	170
rect	113	172	114	173
rect	113	175	114	176
rect	113	178	114	179
rect	113	196	114	197
rect	113	208	114	209
rect	114	1	115	2
rect	114	11	115	12
rect	114	14	115	15
rect	114	16	115	17
rect	114	17	115	18
rect	114	19	115	20
rect	114	22	115	23
rect	114	23	115	24
rect	114	25	115	26
rect	114	26	115	27
rect	114	29	115	30
rect	114	31	115	32
rect	114	34	115	35
rect	114	35	115	36
rect	114	38	115	39
rect	114	47	115	48
rect	114	52	115	53
rect	114	53	115	54
rect	114	54	115	55
rect	114	58	115	59
rect	114	59	115	60
rect	114	60	115	61
rect	114	63	115	64
rect	114	66	115	67
rect	114	72	115	73
rect	114	73	115	74
rect	114	75	115	76
rect	114	81	115	82
rect	114	83	115	84
rect	114	84	115	85
rect	114	88	115	89
rect	114	100	115	101
rect	114	110	115	111
rect	114	112	115	113
rect	114	126	115	127
rect	114	129	115	130
rect	114	132	115	133
rect	114	137	115	138
rect	114	140	115	141
rect	114	160	115	161
rect	114	166	115	167
rect	114	169	115	170
rect	114	172	115	173
rect	114	178	115	179
rect	114	196	115	197
rect	114	208	115	209
rect	115	1	116	2
rect	115	11	116	12
rect	115	14	116	15
rect	115	16	116	17
rect	115	17	116	18
rect	115	19	116	20
rect	115	20	116	21
rect	115	22	116	23
rect	115	23	116	24
rect	115	25	116	26
rect	115	26	116	27
rect	115	29	116	30
rect	115	31	116	32
rect	115	34	116	35
rect	115	35	116	36
rect	115	38	116	39
rect	115	47	116	48
rect	115	52	116	53
rect	115	53	116	54
rect	115	54	116	55
rect	115	57	116	58
rect	115	58	116	59
rect	115	59	116	60
rect	115	60	116	61
rect	115	63	116	64
rect	115	66	116	67
rect	115	72	116	73
rect	115	73	116	74
rect	115	75	116	76
rect	115	81	116	82
rect	115	83	116	84
rect	115	84	116	85
rect	115	88	116	89
rect	115	91	116	92
rect	115	97	116	98
rect	115	100	116	101
rect	115	110	116	111
rect	115	112	116	113
rect	115	116	116	117
rect	115	126	116	127
rect	115	129	116	130
rect	115	132	116	133
rect	115	137	116	138
rect	115	140	116	141
rect	115	148	116	149
rect	115	157	116	158
rect	115	160	116	161
rect	115	166	116	167
rect	115	169	116	170
rect	115	172	116	173
rect	115	178	116	179
rect	115	196	116	197
rect	115	208	116	209
rect	116	1	117	2
rect	116	11	117	12
rect	116	14	117	15
rect	116	16	117	17
rect	116	17	117	18
rect	116	19	117	20
rect	116	20	117	21
rect	116	22	117	23
rect	116	23	117	24
rect	116	25	117	26
rect	116	26	117	27
rect	116	31	117	32
rect	116	34	117	35
rect	116	35	117	36
rect	116	38	117	39
rect	116	47	117	48
rect	116	52	117	53
rect	116	53	117	54
rect	116	54	117	55
rect	116	57	117	58
rect	116	58	117	59
rect	116	59	117	60
rect	116	60	117	61
rect	116	63	117	64
rect	116	66	117	67
rect	116	73	117	74
rect	116	75	117	76
rect	116	81	117	82
rect	116	88	117	89
rect	116	91	117	92
rect	116	97	117	98
rect	116	100	117	101
rect	116	110	117	111
rect	116	116	117	117
rect	116	126	117	127
rect	116	129	117	130
rect	116	132	117	133
rect	116	140	117	141
rect	116	148	117	149
rect	116	157	117	158
rect	116	160	117	161
rect	116	166	117	167
rect	116	169	117	170
rect	116	178	117	179
rect	116	196	117	197
rect	116	208	117	209
rect	117	1	118	2
rect	117	11	118	12
rect	117	14	118	15
rect	117	16	118	17
rect	117	17	118	18
rect	117	19	118	20
rect	117	20	118	21
rect	117	22	118	23
rect	117	23	118	24
rect	117	25	118	26
rect	117	26	118	27
rect	117	31	118	32
rect	117	34	118	35
rect	117	35	118	36
rect	117	38	118	39
rect	117	47	118	48
rect	117	52	118	53
rect	117	53	118	54
rect	117	54	118	55
rect	117	57	118	58
rect	117	58	118	59
rect	117	59	118	60
rect	117	60	118	61
rect	117	63	118	64
rect	117	66	118	67
rect	117	72	118	73
rect	117	73	118	74
rect	117	75	118	76
rect	117	81	118	82
rect	117	83	118	84
rect	117	84	118	85
rect	117	88	118	89
rect	117	91	118	92
rect	117	94	118	95
rect	117	97	118	98
rect	117	100	118	101
rect	117	104	118	105
rect	117	110	118	111
rect	117	113	118	114
rect	117	116	118	117
rect	117	126	118	127
rect	117	129	118	130
rect	117	132	118	133
rect	117	135	118	136
rect	117	140	118	141
rect	117	142	118	143
rect	117	148	118	149
rect	117	151	118	152
rect	117	157	118	158
rect	117	160	118	161
rect	117	166	118	167
rect	117	169	118	170
rect	117	176	118	177
rect	117	178	118	179
rect	117	196	118	197
rect	117	208	118	209
rect	118	1	119	2
rect	118	11	119	12
rect	118	16	119	17
rect	118	17	119	18
rect	118	19	119	20
rect	118	20	119	21
rect	118	22	119	23
rect	118	23	119	24
rect	118	25	119	26
rect	118	26	119	27
rect	118	31	119	32
rect	118	34	119	35
rect	118	35	119	36
rect	118	38	119	39
rect	118	47	119	48
rect	118	53	119	54
rect	118	54	119	55
rect	118	57	119	58
rect	118	58	119	59
rect	118	59	119	60
rect	118	60	119	61
rect	118	63	119	64
rect	118	66	119	67
rect	118	72	119	73
rect	118	73	119	74
rect	118	75	119	76
rect	118	81	119	82
rect	118	83	119	84
rect	118	84	119	85
rect	118	88	119	89
rect	118	91	119	92
rect	118	94	119	95
rect	118	97	119	98
rect	118	100	119	101
rect	118	104	119	105
rect	118	110	119	111
rect	118	113	119	114
rect	118	116	119	117
rect	118	126	119	127
rect	118	129	119	130
rect	118	132	119	133
rect	118	135	119	136
rect	118	142	119	143
rect	118	148	119	149
rect	118	151	119	152
rect	118	157	119	158
rect	118	160	119	161
rect	118	176	119	177
rect	118	178	119	179
rect	118	196	119	197
rect	118	208	119	209
rect	119	1	120	2
rect	119	11	120	12
rect	119	16	120	17
rect	119	17	120	18
rect	119	19	120	20
rect	119	20	120	21
rect	119	22	120	23
rect	119	23	120	24
rect	119	25	120	26
rect	119	26	120	27
rect	119	28	120	29
rect	119	31	120	32
rect	119	34	120	35
rect	119	35	120	36
rect	119	38	120	39
rect	119	47	120	48
rect	119	53	120	54
rect	119	54	120	55
rect	119	57	120	58
rect	119	58	120	59
rect	119	59	120	60
rect	119	60	120	61
rect	119	63	120	64
rect	119	66	120	67
rect	119	72	120	73
rect	119	73	120	74
rect	119	75	120	76
rect	119	81	120	82
rect	119	83	120	84
rect	119	84	120	85
rect	119	88	120	89
rect	119	91	120	92
rect	119	94	120	95
rect	119	97	120	98
rect	119	100	120	101
rect	119	104	120	105
rect	119	110	120	111
rect	119	113	120	114
rect	119	116	120	117
rect	119	120	120	121
rect	119	126	120	127
rect	119	129	120	130
rect	119	132	120	133
rect	119	135	120	136
rect	119	138	120	139
rect	119	142	120	143
rect	119	148	120	149
rect	119	151	120	152
rect	119	154	120	155
rect	119	157	120	158
rect	119	160	120	161
rect	119	173	120	174
rect	119	176	120	177
rect	119	178	120	179
rect	119	196	120	197
rect	119	208	120	209
rect	120	1	121	2
rect	120	11	121	12
rect	120	16	121	17
rect	120	17	121	18
rect	120	19	121	20
rect	120	20	121	21
rect	120	22	121	23
rect	120	23	121	24
rect	120	25	121	26
rect	120	26	121	27
rect	120	28	121	29
rect	120	31	121	32
rect	120	34	121	35
rect	120	35	121	36
rect	120	38	121	39
rect	120	47	121	48
rect	120	53	121	54
rect	120	54	121	55
rect	120	57	121	58
rect	120	58	121	59
rect	120	59	121	60
rect	120	60	121	61
rect	120	63	121	64
rect	120	66	121	67
rect	120	72	121	73
rect	120	73	121	74
rect	120	75	121	76
rect	120	81	121	82
rect	120	83	121	84
rect	120	84	121	85
rect	120	88	121	89
rect	120	91	121	92
rect	120	94	121	95
rect	120	97	121	98
rect	120	100	121	101
rect	120	104	121	105
rect	120	110	121	111
rect	120	113	121	114
rect	120	116	121	117
rect	120	120	121	121
rect	120	126	121	127
rect	120	129	121	130
rect	120	132	121	133
rect	120	135	121	136
rect	120	138	121	139
rect	120	142	121	143
rect	120	148	121	149
rect	120	151	121	152
rect	120	154	121	155
rect	120	157	121	158
rect	120	173	121	174
rect	120	176	121	177
rect	120	196	121	197
rect	120	208	121	209
rect	121	1	122	2
rect	121	4	122	5
rect	121	11	122	12
rect	121	16	122	17
rect	121	17	122	18
rect	121	19	122	20
rect	121	20	122	21
rect	121	22	122	23
rect	121	23	122	24
rect	121	25	122	26
rect	121	26	122	27
rect	121	28	122	29
rect	121	31	122	32
rect	121	34	122	35
rect	121	35	122	36
rect	121	38	122	39
rect	121	41	122	42
rect	121	44	122	45
rect	121	47	122	48
rect	121	51	122	52
rect	121	53	122	54
rect	121	54	122	55
rect	121	57	122	58
rect	121	58	122	59
rect	121	59	122	60
rect	121	60	122	61
rect	121	63	122	64
rect	121	66	122	67
rect	121	69	122	70
rect	121	72	122	73
rect	121	73	122	74
rect	121	75	122	76
rect	121	78	122	79
rect	121	81	122	82
rect	121	83	122	84
rect	121	84	122	85
rect	121	88	122	89
rect	121	91	122	92
rect	121	94	122	95
rect	121	97	122	98
rect	121	100	122	101
rect	121	104	122	105
rect	121	110	122	111
rect	121	113	122	114
rect	121	116	122	117
rect	121	120	122	121
rect	121	126	122	127
rect	121	129	122	130
rect	121	132	122	133
rect	121	135	122	136
rect	121	138	122	139
rect	121	142	122	143
rect	121	148	122	149
rect	121	151	122	152
rect	121	154	122	155
rect	121	157	122	158
rect	121	164	122	165
rect	121	170	122	171
rect	121	173	122	174
rect	121	176	122	177
rect	121	182	122	183
rect	121	196	122	197
rect	121	208	122	209
rect	122	4	123	5
rect	122	16	123	17
rect	122	17	123	18
rect	122	19	123	20
rect	122	20	123	21
rect	122	22	123	23
rect	122	25	123	26
rect	122	26	123	27
rect	122	28	123	29
rect	122	31	123	32
rect	122	34	123	35
rect	122	35	123	36
rect	122	38	123	39
rect	122	41	123	42
rect	122	44	123	45
rect	122	47	123	48
rect	122	51	123	52
rect	122	53	123	54
rect	122	54	123	55
rect	122	57	123	58
rect	122	58	123	59
rect	122	59	123	60
rect	122	60	123	61
rect	122	63	123	64
rect	122	66	123	67
rect	122	69	123	70
rect	122	72	123	73
rect	122	73	123	74
rect	122	75	123	76
rect	122	78	123	79
rect	122	81	123	82
rect	122	83	123	84
rect	122	84	123	85
rect	122	88	123	89
rect	122	91	123	92
rect	122	94	123	95
rect	122	97	123	98
rect	122	100	123	101
rect	122	104	123	105
rect	122	110	123	111
rect	122	113	123	114
rect	122	116	123	117
rect	122	120	123	121
rect	122	126	123	127
rect	122	129	123	130
rect	122	132	123	133
rect	122	135	123	136
rect	122	138	123	139
rect	122	142	123	143
rect	122	148	123	149
rect	122	151	123	152
rect	122	154	123	155
rect	122	157	123	158
rect	122	164	123	165
rect	122	170	123	171
rect	122	173	123	174
rect	122	176	123	177
rect	122	182	123	183
rect	122	196	123	197
rect	122	208	123	209
rect	123	4	124	5
rect	123	7	124	8
rect	123	13	124	14
rect	123	16	124	17
rect	123	17	124	18
rect	123	19	124	20
rect	123	20	124	21
rect	123	22	124	23
rect	123	23	124	24
rect	123	25	124	26
rect	123	26	124	27
rect	123	28	124	29
rect	123	31	124	32
rect	123	34	124	35
rect	123	35	124	36
rect	123	38	124	39
rect	123	41	124	42
rect	123	44	124	45
rect	123	47	124	48
rect	123	51	124	52
rect	123	53	124	54
rect	123	54	124	55
rect	123	57	124	58
rect	123	58	124	59
rect	123	59	124	60
rect	123	60	124	61
rect	123	63	124	64
rect	123	66	124	67
rect	123	69	124	70
rect	123	72	124	73
rect	123	73	124	74
rect	123	75	124	76
rect	123	78	124	79
rect	123	81	124	82
rect	123	83	124	84
rect	123	84	124	85
rect	123	88	124	89
rect	123	91	124	92
rect	123	94	124	95
rect	123	97	124	98
rect	123	100	124	101
rect	123	104	124	105
rect	123	110	124	111
rect	123	113	124	114
rect	123	116	124	117
rect	123	120	124	121
rect	123	126	124	127
rect	123	129	124	130
rect	123	132	124	133
rect	123	135	124	136
rect	123	138	124	139
rect	123	142	124	143
rect	123	148	124	149
rect	123	151	124	152
rect	123	154	124	155
rect	123	157	124	158
rect	123	164	124	165
rect	123	170	124	171
rect	123	173	124	174
rect	123	176	124	177
rect	123	182	124	183
rect	123	193	124	194
rect	123	196	124	197
rect	123	208	124	209
rect	124	4	125	5
rect	124	7	125	8
rect	124	13	125	14
rect	124	16	125	17
rect	124	17	125	18
rect	124	19	125	20
rect	124	20	125	21
rect	124	22	125	23
rect	124	23	125	24
rect	124	25	125	26
rect	124	26	125	27
rect	124	28	125	29
rect	124	31	125	32
rect	124	34	125	35
rect	124	35	125	36
rect	124	38	125	39
rect	124	41	125	42
rect	124	44	125	45
rect	124	47	125	48
rect	124	51	125	52
rect	124	53	125	54
rect	124	54	125	55
rect	124	57	125	58
rect	124	58	125	59
rect	124	59	125	60
rect	124	60	125	61
rect	124	63	125	64
rect	124	66	125	67
rect	124	69	125	70
rect	124	72	125	73
rect	124	73	125	74
rect	124	75	125	76
rect	124	78	125	79
rect	124	81	125	82
rect	124	83	125	84
rect	124	84	125	85
rect	124	88	125	89
rect	124	91	125	92
rect	124	94	125	95
rect	124	97	125	98
rect	124	100	125	101
rect	124	104	125	105
rect	124	110	125	111
rect	124	113	125	114
rect	124	116	125	117
rect	124	120	125	121
rect	124	126	125	127
rect	124	129	125	130
rect	124	132	125	133
rect	124	135	125	136
rect	124	138	125	139
rect	124	142	125	143
rect	124	148	125	149
rect	124	151	125	152
rect	124	154	125	155
rect	124	157	125	158
rect	124	164	125	165
rect	124	170	125	171
rect	124	173	125	174
rect	124	176	125	177
rect	124	182	125	183
rect	124	193	125	194
rect	124	196	125	197
rect	125	1	126	2
rect	125	4	126	5
rect	125	7	126	8
rect	125	10	126	11
rect	125	13	126	14
rect	125	16	126	17
rect	125	17	126	18
rect	125	19	126	20
rect	125	20	126	21
rect	125	22	126	23
rect	125	23	126	24
rect	125	25	126	26
rect	125	26	126	27
rect	125	28	126	29
rect	125	31	126	32
rect	125	34	126	35
rect	125	35	126	36
rect	125	38	126	39
rect	125	41	126	42
rect	125	44	126	45
rect	125	47	126	48
rect	125	51	126	52
rect	125	53	126	54
rect	125	54	126	55
rect	125	57	126	58
rect	125	58	126	59
rect	125	59	126	60
rect	125	60	126	61
rect	125	63	126	64
rect	125	66	126	67
rect	125	69	126	70
rect	125	72	126	73
rect	125	73	126	74
rect	125	75	126	76
rect	125	78	126	79
rect	125	81	126	82
rect	125	83	126	84
rect	125	84	126	85
rect	125	88	126	89
rect	125	91	126	92
rect	125	94	126	95
rect	125	97	126	98
rect	125	100	126	101
rect	125	104	126	105
rect	125	110	126	111
rect	125	113	126	114
rect	125	116	126	117
rect	125	120	126	121
rect	125	126	126	127
rect	125	129	126	130
rect	125	132	126	133
rect	125	135	126	136
rect	125	138	126	139
rect	125	142	126	143
rect	125	145	126	146
rect	125	148	126	149
rect	125	151	126	152
rect	125	154	126	155
rect	125	157	126	158
rect	125	161	126	162
rect	125	164	126	165
rect	125	167	126	168
rect	125	170	126	171
rect	125	173	126	174
rect	125	176	126	177
rect	125	179	126	180
rect	125	182	126	183
rect	125	193	126	194
rect	125	196	126	197
rect	126	16	127	17
rect	126	17	127	18
rect	126	19	127	20
rect	126	20	127	21
rect	126	22	127	23
rect	126	23	127	24
rect	126	25	127	26
rect	126	26	127	27
rect	126	34	127	35
rect	126	35	127	36
rect	126	53	127	54
rect	126	54	127	55
rect	126	58	127	59
rect	126	59	127	60
rect	126	72	127	73
rect	126	73	127	74
rect	126	83	127	84
rect	126	84	127	85
rect	127	16	128	17
rect	127	17	128	18
rect	127	19	128	20
rect	127	20	128	21
rect	127	22	128	23
rect	127	23	128	24
rect	127	25	128	26
rect	127	26	128	27
rect	127	34	128	35
rect	127	35	128	36
rect	127	53	128	54
rect	127	54	128	55
rect	127	58	128	59
rect	127	59	128	60
rect	127	72	128	73
rect	127	73	128	74
rect	127	83	128	84
rect	127	84	128	85
rect	128	16	129	17
rect	128	17	129	18
rect	128	19	129	20
rect	128	20	129	21
rect	128	22	129	23
rect	128	23	129	24
rect	128	25	129	26
rect	128	26	129	27
rect	128	34	129	35
rect	128	35	129	36
rect	128	53	129	54
rect	128	54	129	55
rect	128	58	129	59
rect	128	59	129	60
rect	128	72	129	73
rect	128	73	129	74
rect	128	83	129	84
rect	128	84	129	85
rect	129	16	130	17
rect	129	17	130	18
rect	129	19	130	20
rect	129	20	130	21
rect	129	22	130	23
rect	129	23	130	24
rect	129	25	130	26
rect	129	26	130	27
rect	129	34	130	35
rect	129	35	130	36
rect	129	53	130	54
rect	129	54	130	55
rect	129	58	130	59
rect	129	59	130	60
rect	129	72	130	73
rect	129	73	130	74
rect	129	83	130	84
rect	129	84	130	85
rect	130	16	131	17
rect	130	17	131	18
rect	130	19	131	20
rect	130	20	131	21
rect	130	22	131	23
rect	130	23	131	24
rect	130	25	131	26
rect	130	26	131	27
rect	130	34	131	35
rect	130	35	131	36
rect	130	53	131	54
rect	130	54	131	55
rect	130	58	131	59
rect	130	59	131	60
rect	130	72	131	73
rect	130	73	131	74
rect	130	83	131	84
rect	130	84	131	85
rect	131	16	132	17
rect	131	17	132	18
rect	131	19	132	20
rect	131	20	132	21
rect	131	22	132	23
rect	131	23	132	24
rect	131	25	132	26
rect	131	26	132	27
rect	131	35	132	36
rect	131	53	132	54
rect	131	54	132	55
rect	131	58	132	59
rect	131	59	132	60
rect	131	72	132	73
rect	131	73	132	74
rect	131	83	132	84
rect	131	84	132	85
rect	132	1	133	2
rect	132	4	133	5
rect	132	7	133	8
rect	132	10	133	11
rect	132	13	133	14
rect	132	16	133	17
rect	132	17	133	18
rect	132	19	133	20
rect	132	20	133	21
rect	132	22	133	23
rect	132	23	133	24
rect	132	25	133	26
rect	132	26	133	27
rect	132	28	133	29
rect	132	31	133	32
rect	132	35	133	36
rect	132	41	133	42
rect	132	44	133	45
rect	132	47	133	48
rect	132	53	133	54
rect	132	54	133	55
rect	132	57	133	58
rect	132	58	133	59
rect	132	59	133	60
rect	132	60	133	61
rect	132	63	133	64
rect	132	66	133	67
rect	132	69	133	70
rect	132	72	133	73
rect	132	73	133	74
rect	132	75	133	76
rect	132	78	133	79
rect	132	81	133	82
rect	132	83	133	84
rect	132	84	133	85
rect	132	88	133	89
rect	132	94	133	95
rect	132	97	133	98
rect	132	100	133	101
rect	132	104	133	105
rect	132	110	133	111
rect	132	113	133	114
rect	132	116	133	117
rect	132	126	133	127
rect	132	129	133	130
rect	132	132	133	133
rect	132	135	133	136
rect	132	138	133	139
rect	132	145	133	146
rect	132	148	133	149
rect	132	151	133	152
rect	132	154	133	155
rect	132	157	133	158
rect	132	161	133	162
rect	132	164	133	165
rect	132	167	133	168
rect	132	170	133	171
rect	132	173	133	174
rect	132	176	133	177
rect	132	179	133	180
rect	132	182	133	183
rect	132	186	133	187
rect	132	193	133	194
rect	132	196	133	197
rect	133	1	134	2
rect	133	4	134	5
rect	133	7	134	8
rect	133	10	134	11
rect	133	13	134	14
rect	133	16	134	17
rect	133	17	134	18
rect	133	19	134	20
rect	133	20	134	21
rect	133	22	134	23
rect	133	23	134	24
rect	133	25	134	26
rect	133	26	134	27
rect	133	28	134	29
rect	133	31	134	32
rect	133	35	134	36
rect	133	41	134	42
rect	133	44	134	45
rect	133	47	134	48
rect	133	53	134	54
rect	133	54	134	55
rect	133	57	134	58
rect	133	58	134	59
rect	133	59	134	60
rect	133	60	134	61
rect	133	63	134	64
rect	133	66	134	67
rect	133	69	134	70
rect	133	72	134	73
rect	133	73	134	74
rect	133	75	134	76
rect	133	78	134	79
rect	133	81	134	82
rect	133	83	134	84
rect	133	84	134	85
rect	133	88	134	89
rect	133	94	134	95
rect	133	97	134	98
rect	133	100	134	101
rect	133	104	134	105
rect	133	110	134	111
rect	133	113	134	114
rect	133	116	134	117
rect	133	126	134	127
rect	133	129	134	130
rect	133	132	134	133
rect	133	135	134	136
rect	133	138	134	139
rect	133	145	134	146
rect	133	148	134	149
rect	133	151	134	152
rect	133	154	134	155
rect	133	157	134	158
rect	133	161	134	162
rect	133	164	134	165
rect	133	167	134	168
rect	133	170	134	171
rect	133	173	134	174
rect	133	176	134	177
rect	133	179	134	180
rect	133	182	134	183
rect	133	186	134	187
rect	133	193	134	194
rect	133	196	134	197
rect	134	1	135	2
rect	134	4	135	5
rect	134	7	135	8
rect	134	10	135	11
rect	134	13	135	14
rect	134	16	135	17
rect	134	17	135	18
rect	134	19	135	20
rect	134	20	135	21
rect	134	22	135	23
rect	134	23	135	24
rect	134	25	135	26
rect	134	26	135	27
rect	134	28	135	29
rect	134	31	135	32
rect	134	35	135	36
rect	134	41	135	42
rect	134	44	135	45
rect	134	47	135	48
rect	134	53	135	54
rect	134	54	135	55
rect	134	57	135	58
rect	134	58	135	59
rect	134	59	135	60
rect	134	60	135	61
rect	134	63	135	64
rect	134	66	135	67
rect	134	69	135	70
rect	134	72	135	73
rect	134	73	135	74
rect	134	75	135	76
rect	134	78	135	79
rect	134	81	135	82
rect	134	83	135	84
rect	134	84	135	85
rect	134	88	135	89
rect	134	94	135	95
rect	134	97	135	98
rect	134	100	135	101
rect	134	104	135	105
rect	134	110	135	111
rect	134	113	135	114
rect	134	116	135	117
rect	134	126	135	127
rect	134	129	135	130
rect	134	132	135	133
rect	134	135	135	136
rect	134	138	135	139
rect	134	145	135	146
rect	134	148	135	149
rect	134	151	135	152
rect	134	154	135	155
rect	134	157	135	158
rect	134	161	135	162
rect	134	164	135	165
rect	134	167	135	168
rect	134	170	135	171
rect	134	173	135	174
rect	134	176	135	177
rect	134	179	135	180
rect	134	182	135	183
rect	134	186	135	187
rect	134	193	135	194
rect	134	196	135	197
rect	135	1	136	2
rect	135	4	136	5
rect	135	7	136	8
rect	135	10	136	11
rect	135	13	136	14
rect	135	16	136	17
rect	135	17	136	18
rect	135	19	136	20
rect	135	20	136	21
rect	135	22	136	23
rect	135	23	136	24
rect	135	25	136	26
rect	135	26	136	27
rect	135	28	136	29
rect	135	31	136	32
rect	135	35	136	36
rect	135	41	136	42
rect	135	44	136	45
rect	135	47	136	48
rect	135	53	136	54
rect	135	54	136	55
rect	135	57	136	58
rect	135	58	136	59
rect	135	59	136	60
rect	135	60	136	61
rect	135	63	136	64
rect	135	66	136	67
rect	135	69	136	70
rect	135	72	136	73
rect	135	73	136	74
rect	135	75	136	76
rect	135	78	136	79
rect	135	81	136	82
rect	135	83	136	84
rect	135	84	136	85
rect	135	88	136	89
rect	135	94	136	95
rect	135	97	136	98
rect	135	100	136	101
rect	135	104	136	105
rect	135	110	136	111
rect	135	113	136	114
rect	135	116	136	117
rect	135	126	136	127
rect	135	129	136	130
rect	135	132	136	133
rect	135	135	136	136
rect	135	138	136	139
rect	135	145	136	146
rect	135	148	136	149
rect	135	151	136	152
rect	135	154	136	155
rect	135	157	136	158
rect	135	161	136	162
rect	135	164	136	165
rect	135	167	136	168
rect	135	170	136	171
rect	135	173	136	174
rect	135	176	136	177
rect	135	179	136	180
rect	135	182	136	183
rect	135	186	136	187
rect	135	193	136	194
rect	135	196	136	197
rect	136	1	137	2
rect	136	4	137	5
rect	136	7	137	8
rect	136	10	137	11
rect	136	13	137	14
rect	136	16	137	17
rect	136	17	137	18
rect	136	19	137	20
rect	136	20	137	21
rect	136	22	137	23
rect	136	23	137	24
rect	136	25	137	26
rect	136	26	137	27
rect	136	28	137	29
rect	136	31	137	32
rect	136	35	137	36
rect	136	41	137	42
rect	136	44	137	45
rect	136	47	137	48
rect	136	53	137	54
rect	136	54	137	55
rect	136	57	137	58
rect	136	58	137	59
rect	136	59	137	60
rect	136	60	137	61
rect	136	63	137	64
rect	136	66	137	67
rect	136	69	137	70
rect	136	72	137	73
rect	136	73	137	74
rect	136	75	137	76
rect	136	78	137	79
rect	136	81	137	82
rect	136	83	137	84
rect	136	84	137	85
rect	136	88	137	89
rect	136	94	137	95
rect	136	97	137	98
rect	136	100	137	101
rect	136	104	137	105
rect	136	110	137	111
rect	136	113	137	114
rect	136	116	137	117
rect	136	126	137	127
rect	136	129	137	130
rect	136	132	137	133
rect	136	135	137	136
rect	136	138	137	139
rect	136	145	137	146
rect	136	148	137	149
rect	136	151	137	152
rect	136	154	137	155
rect	136	157	137	158
rect	136	161	137	162
rect	136	164	137	165
rect	136	167	137	168
rect	136	170	137	171
rect	136	173	137	174
rect	136	176	137	177
rect	136	179	137	180
rect	136	182	137	183
rect	136	186	137	187
rect	136	193	137	194
rect	136	196	137	197
rect	137	1	138	2
rect	137	4	138	5
rect	137	7	138	8
rect	137	10	138	11
rect	137	13	138	14
rect	137	16	138	17
rect	137	17	138	18
rect	137	19	138	20
rect	137	20	138	21
rect	137	22	138	23
rect	137	23	138	24
rect	137	25	138	26
rect	137	26	138	27
rect	137	28	138	29
rect	137	31	138	32
rect	137	35	138	36
rect	137	41	138	42
rect	137	44	138	45
rect	137	47	138	48
rect	137	53	138	54
rect	137	54	138	55
rect	137	57	138	58
rect	137	58	138	59
rect	137	59	138	60
rect	137	60	138	61
rect	137	63	138	64
rect	137	66	138	67
rect	137	69	138	70
rect	137	72	138	73
rect	137	73	138	74
rect	137	75	138	76
rect	137	78	138	79
rect	137	81	138	82
rect	137	83	138	84
rect	137	84	138	85
rect	137	88	138	89
rect	137	94	138	95
rect	137	97	138	98
rect	137	100	138	101
rect	137	104	138	105
rect	137	110	138	111
rect	137	113	138	114
rect	137	116	138	117
rect	137	126	138	127
rect	137	129	138	130
rect	137	132	138	133
rect	137	135	138	136
rect	137	138	138	139
rect	137	145	138	146
rect	137	148	138	149
rect	137	151	138	152
rect	137	154	138	155
rect	137	157	138	158
rect	137	161	138	162
rect	137	164	138	165
rect	137	167	138	168
rect	137	170	138	171
rect	137	173	138	174
rect	137	176	138	177
rect	137	179	138	180
rect	137	182	138	183
rect	137	186	138	187
rect	137	193	138	194
rect	137	196	138	197
rect	138	1	139	2
rect	138	4	139	5
rect	138	7	139	8
rect	138	10	139	11
rect	138	13	139	14
rect	138	16	139	17
rect	138	17	139	18
rect	138	19	139	20
rect	138	20	139	21
rect	138	22	139	23
rect	138	23	139	24
rect	138	25	139	26
rect	138	26	139	27
rect	138	28	139	29
rect	138	31	139	32
rect	138	35	139	36
rect	138	41	139	42
rect	138	44	139	45
rect	138	47	139	48
rect	138	53	139	54
rect	138	54	139	55
rect	138	57	139	58
rect	138	58	139	59
rect	138	59	139	60
rect	138	60	139	61
rect	138	63	139	64
rect	138	66	139	67
rect	138	69	139	70
rect	138	72	139	73
rect	138	73	139	74
rect	138	75	139	76
rect	138	78	139	79
rect	138	81	139	82
rect	138	83	139	84
rect	138	84	139	85
rect	138	88	139	89
rect	138	94	139	95
rect	138	97	139	98
rect	138	100	139	101
rect	138	104	139	105
rect	138	110	139	111
rect	138	113	139	114
rect	138	116	139	117
rect	138	126	139	127
rect	138	129	139	130
rect	138	132	139	133
rect	138	135	139	136
rect	138	138	139	139
rect	138	145	139	146
rect	138	148	139	149
rect	138	151	139	152
rect	138	154	139	155
rect	138	157	139	158
rect	138	161	139	162
rect	138	164	139	165
rect	138	167	139	168
rect	138	170	139	171
rect	138	173	139	174
rect	138	176	139	177
rect	138	179	139	180
rect	138	182	139	183
rect	138	186	139	187
rect	138	193	139	194
rect	138	196	139	197
rect	139	1	140	2
rect	139	4	140	5
rect	139	7	140	8
rect	139	10	140	11
rect	139	13	140	14
rect	139	16	140	17
rect	139	17	140	18
rect	139	19	140	20
rect	139	20	140	21
rect	139	22	140	23
rect	139	23	140	24
rect	139	25	140	26
rect	139	26	140	27
rect	139	28	140	29
rect	139	31	140	32
rect	139	35	140	36
rect	139	41	140	42
rect	139	44	140	45
rect	139	47	140	48
rect	139	53	140	54
rect	139	54	140	55
rect	139	57	140	58
rect	139	58	140	59
rect	139	59	140	60
rect	139	60	140	61
rect	139	63	140	64
rect	139	66	140	67
rect	139	69	140	70
rect	139	72	140	73
rect	139	73	140	74
rect	139	75	140	76
rect	139	78	140	79
rect	139	81	140	82
rect	139	83	140	84
rect	139	84	140	85
rect	139	88	140	89
rect	139	94	140	95
rect	139	100	140	101
rect	139	110	140	111
rect	139	113	140	114
rect	139	116	140	117
rect	139	126	140	127
rect	139	129	140	130
rect	139	132	140	133
rect	139	135	140	136
rect	139	138	140	139
rect	139	145	140	146
rect	139	148	140	149
rect	139	151	140	152
rect	139	154	140	155
rect	139	157	140	158
rect	139	161	140	162
rect	139	164	140	165
rect	139	167	140	168
rect	139	170	140	171
rect	139	173	140	174
rect	139	176	140	177
rect	139	179	140	180
rect	139	182	140	183
rect	139	186	140	187
rect	139	193	140	194
rect	139	196	140	197
rect	140	1	141	2
rect	140	4	141	5
rect	140	7	141	8
rect	140	10	141	11
rect	140	13	141	14
rect	140	16	141	17
rect	140	17	141	18
rect	140	19	141	20
rect	140	20	141	21
rect	140	22	141	23
rect	140	23	141	24
rect	140	25	141	26
rect	140	26	141	27
rect	140	28	141	29
rect	140	31	141	32
rect	140	35	141	36
rect	140	41	141	42
rect	140	44	141	45
rect	140	47	141	48
rect	140	53	141	54
rect	140	54	141	55
rect	140	57	141	58
rect	140	58	141	59
rect	140	59	141	60
rect	140	60	141	61
rect	140	63	141	64
rect	140	66	141	67
rect	140	69	141	70
rect	140	72	141	73
rect	140	73	141	74
rect	140	75	141	76
rect	140	78	141	79
rect	140	81	141	82
rect	140	83	141	84
rect	140	84	141	85
rect	140	88	141	89
rect	140	94	141	95
rect	140	100	141	101
rect	140	110	141	111
rect	140	113	141	114
rect	140	116	141	117
rect	140	126	141	127
rect	140	129	141	130
rect	140	132	141	133
rect	140	135	141	136
rect	140	138	141	139
rect	140	145	141	146
rect	140	148	141	149
rect	140	151	141	152
rect	140	154	141	155
rect	140	157	141	158
rect	140	161	141	162
rect	140	164	141	165
rect	140	167	141	168
rect	140	170	141	171
rect	140	173	141	174
rect	140	176	141	177
rect	140	179	141	180
rect	140	182	141	183
rect	140	186	141	187
rect	140	193	141	194
rect	140	196	141	197
rect	141	1	142	2
rect	141	4	142	5
rect	141	7	142	8
rect	141	10	142	11
rect	141	13	142	14
rect	141	16	142	17
rect	141	17	142	18
rect	141	19	142	20
rect	141	20	142	21
rect	141	22	142	23
rect	141	23	142	24
rect	141	25	142	26
rect	141	26	142	27
rect	141	28	142	29
rect	141	31	142	32
rect	141	35	142	36
rect	141	41	142	42
rect	141	44	142	45
rect	141	47	142	48
rect	141	53	142	54
rect	141	54	142	55
rect	141	58	142	59
rect	141	59	142	60
rect	141	60	142	61
rect	141	63	142	64
rect	141	66	142	67
rect	141	69	142	70
rect	141	72	142	73
rect	141	73	142	74
rect	141	75	142	76
rect	141	78	142	79
rect	141	81	142	82
rect	141	83	142	84
rect	141	84	142	85
rect	141	88	142	89
rect	141	94	142	95
rect	141	100	142	101
rect	141	110	142	111
rect	141	113	142	114
rect	141	116	142	117
rect	141	126	142	127
rect	141	129	142	130
rect	141	132	142	133
rect	141	135	142	136
rect	141	138	142	139
rect	141	145	142	146
rect	141	148	142	149
rect	141	151	142	152
rect	141	154	142	155
rect	141	157	142	158
rect	141	161	142	162
rect	141	164	142	165
rect	141	167	142	168
rect	141	170	142	171
rect	141	173	142	174
rect	141	176	142	177
rect	141	179	142	180
rect	141	182	142	183
rect	141	186	142	187
rect	141	193	142	194
rect	141	196	142	197
rect	142	1	143	2
rect	142	4	143	5
rect	142	7	143	8
rect	142	10	143	11
rect	142	13	143	14
rect	142	16	143	17
rect	142	17	143	18
rect	142	19	143	20
rect	142	20	143	21
rect	142	22	143	23
rect	142	23	143	24
rect	142	25	143	26
rect	142	26	143	27
rect	142	28	143	29
rect	142	31	143	32
rect	142	35	143	36
rect	142	41	143	42
rect	142	44	143	45
rect	142	47	143	48
rect	142	53	143	54
rect	142	54	143	55
rect	142	58	143	59
rect	142	59	143	60
rect	142	60	143	61
rect	142	63	143	64
rect	142	66	143	67
rect	142	69	143	70
rect	142	72	143	73
rect	142	73	143	74
rect	142	75	143	76
rect	142	78	143	79
rect	142	81	143	82
rect	142	83	143	84
rect	142	84	143	85
rect	142	88	143	89
rect	142	94	143	95
rect	142	97	143	98
rect	142	100	143	101
rect	142	110	143	111
rect	142	113	143	114
rect	142	116	143	117
rect	142	126	143	127
rect	142	129	143	130
rect	142	132	143	133
rect	142	135	143	136
rect	142	138	143	139
rect	142	145	143	146
rect	142	148	143	149
rect	142	151	143	152
rect	142	154	143	155
rect	142	157	143	158
rect	142	161	143	162
rect	142	164	143	165
rect	142	167	143	168
rect	142	170	143	171
rect	142	173	143	174
rect	142	176	143	177
rect	142	179	143	180
rect	142	182	143	183
rect	142	186	143	187
rect	142	193	143	194
rect	142	196	143	197
rect	143	1	144	2
rect	143	4	144	5
rect	143	7	144	8
rect	143	10	144	11
rect	143	13	144	14
rect	143	16	144	17
rect	143	17	144	18
rect	143	19	144	20
rect	143	20	144	21
rect	143	22	144	23
rect	143	23	144	24
rect	143	25	144	26
rect	143	26	144	27
rect	143	28	144	29
rect	143	31	144	32
rect	143	35	144	36
rect	143	41	144	42
rect	143	44	144	45
rect	143	47	144	48
rect	143	53	144	54
rect	143	54	144	55
rect	143	58	144	59
rect	143	59	144	60
rect	143	60	144	61
rect	143	63	144	64
rect	143	66	144	67
rect	143	69	144	70
rect	143	72	144	73
rect	143	73	144	74
rect	143	75	144	76
rect	143	81	144	82
rect	143	83	144	84
rect	143	84	144	85
rect	143	88	144	89
rect	143	94	144	95
rect	143	97	144	98
rect	143	100	144	101
rect	143	110	144	111
rect	143	113	144	114
rect	143	116	144	117
rect	143	126	144	127
rect	143	129	144	130
rect	143	132	144	133
rect	143	135	144	136
rect	143	138	144	139
rect	143	145	144	146
rect	143	148	144	149
rect	143	151	144	152
rect	143	154	144	155
rect	143	157	144	158
rect	143	161	144	162
rect	143	164	144	165
rect	143	167	144	168
rect	143	170	144	171
rect	143	173	144	174
rect	143	176	144	177
rect	143	179	144	180
rect	143	182	144	183
rect	143	186	144	187
rect	143	193	144	194
rect	143	196	144	197
rect	144	1	145	2
rect	144	4	145	5
rect	144	7	145	8
rect	144	10	145	11
rect	144	13	145	14
rect	144	16	145	17
rect	144	17	145	18
rect	144	19	145	20
rect	144	20	145	21
rect	144	22	145	23
rect	144	23	145	24
rect	144	25	145	26
rect	144	26	145	27
rect	144	28	145	29
rect	144	31	145	32
rect	144	35	145	36
rect	144	41	145	42
rect	144	44	145	45
rect	144	47	145	48
rect	144	53	145	54
rect	144	54	145	55
rect	144	56	145	57
rect	144	58	145	59
rect	144	59	145	60
rect	144	60	145	61
rect	144	63	145	64
rect	144	66	145	67
rect	144	69	145	70
rect	144	72	145	73
rect	144	73	145	74
rect	144	75	145	76
rect	144	81	145	82
rect	144	83	145	84
rect	144	84	145	85
rect	144	88	145	89
rect	144	94	145	95
rect	144	97	145	98
rect	144	100	145	101
rect	144	110	145	111
rect	144	113	145	114
rect	144	116	145	117
rect	144	126	145	127
rect	144	129	145	130
rect	144	132	145	133
rect	144	135	145	136
rect	144	138	145	139
rect	144	145	145	146
rect	144	148	145	149
rect	144	151	145	152
rect	144	154	145	155
rect	144	157	145	158
rect	144	161	145	162
rect	144	164	145	165
rect	144	167	145	168
rect	144	170	145	171
rect	144	173	145	174
rect	144	176	145	177
rect	144	179	145	180
rect	144	182	145	183
rect	144	186	145	187
rect	144	193	145	194
rect	144	196	145	197
rect	145	1	146	2
rect	145	4	146	5
rect	145	7	146	8
rect	145	10	146	11
rect	145	13	146	14
rect	145	16	146	17
rect	145	17	146	18
rect	145	19	146	20
rect	145	20	146	21
rect	145	22	146	23
rect	145	23	146	24
rect	145	25	146	26
rect	145	26	146	27
rect	145	28	146	29
rect	145	31	146	32
rect	145	35	146	36
rect	145	41	146	42
rect	145	44	146	45
rect	145	47	146	48
rect	145	53	146	54
rect	145	54	146	55
rect	145	56	146	57
rect	145	58	146	59
rect	145	59	146	60
rect	145	60	146	61
rect	145	63	146	64
rect	145	66	146	67
rect	145	69	146	70
rect	145	72	146	73
rect	145	73	146	74
rect	145	75	146	76
rect	145	81	146	82
rect	145	83	146	84
rect	145	84	146	85
rect	145	94	146	95
rect	145	97	146	98
rect	145	100	146	101
rect	145	110	146	111
rect	145	113	146	114
rect	145	116	146	117
rect	145	126	146	127
rect	145	129	146	130
rect	145	132	146	133
rect	145	135	146	136
rect	145	138	146	139
rect	145	145	146	146
rect	145	148	146	149
rect	145	151	146	152
rect	145	154	146	155
rect	145	157	146	158
rect	145	161	146	162
rect	145	164	146	165
rect	145	167	146	168
rect	145	170	146	171
rect	145	173	146	174
rect	145	176	146	177
rect	145	179	146	180
rect	145	182	146	183
rect	145	186	146	187
rect	145	193	146	194
rect	145	196	146	197
rect	146	1	147	2
rect	146	4	147	5
rect	146	7	147	8
rect	146	10	147	11
rect	146	13	147	14
rect	146	16	147	17
rect	146	17	147	18
rect	146	19	147	20
rect	146	20	147	21
rect	146	22	147	23
rect	146	23	147	24
rect	146	25	147	26
rect	146	26	147	27
rect	146	28	147	29
rect	146	31	147	32
rect	146	35	147	36
rect	146	41	147	42
rect	146	44	147	45
rect	146	47	147	48
rect	146	53	147	54
rect	146	54	147	55
rect	146	56	147	57
rect	146	58	147	59
rect	146	59	147	60
rect	146	60	147	61
rect	146	63	147	64
rect	146	66	147	67
rect	146	69	147	70
rect	146	72	147	73
rect	146	73	147	74
rect	146	75	147	76
rect	146	78	147	79
rect	146	81	147	82
rect	146	83	147	84
rect	146	84	147	85
rect	146	94	147	95
rect	146	97	147	98
rect	146	100	147	101
rect	146	110	147	111
rect	146	113	147	114
rect	146	116	147	117
rect	146	126	147	127
rect	146	129	147	130
rect	146	132	147	133
rect	146	135	147	136
rect	146	138	147	139
rect	146	145	147	146
rect	146	148	147	149
rect	146	151	147	152
rect	146	154	147	155
rect	146	157	147	158
rect	146	161	147	162
rect	146	164	147	165
rect	146	167	147	168
rect	146	170	147	171
rect	146	173	147	174
rect	146	176	147	177
rect	146	179	147	180
rect	146	182	147	183
rect	146	186	147	187
rect	146	193	147	194
rect	146	196	147	197
rect	147	1	148	2
rect	147	4	148	5
rect	147	7	148	8
rect	147	10	148	11
rect	147	13	148	14
rect	147	16	148	17
rect	147	17	148	18
rect	147	19	148	20
rect	147	20	148	21
rect	147	22	148	23
rect	147	23	148	24
rect	147	25	148	26
rect	147	26	148	27
rect	147	28	148	29
rect	147	31	148	32
rect	147	35	148	36
rect	147	41	148	42
rect	147	44	148	45
rect	147	47	148	48
rect	147	53	148	54
rect	147	54	148	55
rect	147	56	148	57
rect	147	58	148	59
rect	147	59	148	60
rect	147	60	148	61
rect	147	63	148	64
rect	147	66	148	67
rect	147	69	148	70
rect	147	72	148	73
rect	147	73	148	74
rect	147	78	148	79
rect	147	81	148	82
rect	147	83	148	84
rect	147	84	148	85
rect	147	94	148	95
rect	147	97	148	98
rect	147	100	148	101
rect	147	110	148	111
rect	147	113	148	114
rect	147	116	148	117
rect	147	126	148	127
rect	147	129	148	130
rect	147	132	148	133
rect	147	135	148	136
rect	147	138	148	139
rect	147	145	148	146
rect	147	148	148	149
rect	147	151	148	152
rect	147	154	148	155
rect	147	157	148	158
rect	147	161	148	162
rect	147	164	148	165
rect	147	167	148	168
rect	147	170	148	171
rect	147	173	148	174
rect	147	176	148	177
rect	147	179	148	180
rect	147	182	148	183
rect	147	186	148	187
rect	147	193	148	194
rect	147	196	148	197
rect	148	1	149	2
rect	148	4	149	5
rect	148	7	149	8
rect	148	10	149	11
rect	148	13	149	14
rect	148	16	149	17
rect	148	17	149	18
rect	148	19	149	20
rect	148	20	149	21
rect	148	22	149	23
rect	148	23	149	24
rect	148	25	149	26
rect	148	26	149	27
rect	148	28	149	29
rect	148	31	149	32
rect	148	35	149	36
rect	148	41	149	42
rect	148	44	149	45
rect	148	47	149	48
rect	148	53	149	54
rect	148	54	149	55
rect	148	56	149	57
rect	148	58	149	59
rect	148	59	149	60
rect	148	60	149	61
rect	148	63	149	64
rect	148	66	149	67
rect	148	69	149	70
rect	148	72	149	73
rect	148	73	149	74
rect	148	78	149	79
rect	148	81	149	82
rect	148	83	149	84
rect	148	84	149	85
rect	148	90	149	91
rect	148	94	149	95
rect	148	97	149	98
rect	148	100	149	101
rect	148	110	149	111
rect	148	113	149	114
rect	148	116	149	117
rect	148	126	149	127
rect	148	129	149	130
rect	148	132	149	133
rect	148	135	149	136
rect	148	138	149	139
rect	148	145	149	146
rect	148	148	149	149
rect	148	151	149	152
rect	148	154	149	155
rect	148	157	149	158
rect	148	161	149	162
rect	148	164	149	165
rect	148	167	149	168
rect	148	170	149	171
rect	148	173	149	174
rect	148	176	149	177
rect	148	179	149	180
rect	148	182	149	183
rect	148	186	149	187
rect	148	193	149	194
rect	148	196	149	197
rect	149	1	150	2
rect	149	4	150	5
rect	149	7	150	8
rect	149	10	150	11
rect	149	13	150	14
rect	149	16	150	17
rect	149	17	150	18
rect	149	19	150	20
rect	149	20	150	21
rect	149	22	150	23
rect	149	23	150	24
rect	149	25	150	26
rect	149	26	150	27
rect	149	28	150	29
rect	149	31	150	32
rect	149	35	150	36
rect	149	41	150	42
rect	149	44	150	45
rect	149	47	150	48
rect	149	53	150	54
rect	149	54	150	55
rect	149	56	150	57
rect	149	58	150	59
rect	149	59	150	60
rect	149	60	150	61
rect	149	63	150	64
rect	149	66	150	67
rect	149	69	150	70
rect	149	73	150	74
rect	149	78	150	79
rect	149	81	150	82
rect	149	83	150	84
rect	149	84	150	85
rect	149	90	150	91
rect	149	94	150	95
rect	149	97	150	98
rect	149	100	150	101
rect	149	110	150	111
rect	149	126	150	127
rect	149	129	150	130
rect	149	132	150	133
rect	149	135	150	136
rect	149	138	150	139
rect	149	145	150	146
rect	149	148	150	149
rect	149	151	150	152
rect	149	154	150	155
rect	149	157	150	158
rect	149	161	150	162
rect	149	164	150	165
rect	149	167	150	168
rect	149	170	150	171
rect	149	173	150	174
rect	149	176	150	177
rect	149	179	150	180
rect	149	182	150	183
rect	149	186	150	187
rect	149	193	150	194
rect	149	196	150	197
rect	150	1	151	2
rect	150	4	151	5
rect	150	7	151	8
rect	150	10	151	11
rect	150	13	151	14
rect	150	16	151	17
rect	150	17	151	18
rect	150	19	151	20
rect	150	20	151	21
rect	150	22	151	23
rect	150	23	151	24
rect	150	25	151	26
rect	150	26	151	27
rect	150	28	151	29
rect	150	31	151	32
rect	150	35	151	36
rect	150	41	151	42
rect	150	44	151	45
rect	150	47	151	48
rect	150	53	151	54
rect	150	54	151	55
rect	150	56	151	57
rect	150	58	151	59
rect	150	59	151	60
rect	150	60	151	61
rect	150	63	151	64
rect	150	66	151	67
rect	150	69	151	70
rect	150	72	151	73
rect	150	73	151	74
rect	150	78	151	79
rect	150	81	151	82
rect	150	83	151	84
rect	150	84	151	85
rect	150	87	151	88
rect	150	90	151	91
rect	150	94	151	95
rect	150	97	151	98
rect	150	100	151	101
rect	150	106	151	107
rect	150	110	151	111
rect	150	119	151	120
rect	150	126	151	127
rect	150	129	151	130
rect	150	132	151	133
rect	150	135	151	136
rect	150	138	151	139
rect	150	145	151	146
rect	150	148	151	149
rect	150	151	151	152
rect	150	154	151	155
rect	150	157	151	158
rect	150	161	151	162
rect	150	164	151	165
rect	150	167	151	168
rect	150	170	151	171
rect	150	173	151	174
rect	150	176	151	177
rect	150	179	151	180
rect	150	182	151	183
rect	150	186	151	187
rect	150	193	151	194
rect	150	196	151	197
rect	151	1	152	2
rect	151	4	152	5
rect	151	7	152	8
rect	151	10	152	11
rect	151	13	152	14
rect	151	16	152	17
rect	151	17	152	18
rect	151	19	152	20
rect	151	20	152	21
rect	151	22	152	23
rect	151	23	152	24
rect	151	25	152	26
rect	151	26	152	27
rect	151	28	152	29
rect	151	31	152	32
rect	151	35	152	36
rect	151	41	152	42
rect	151	44	152	45
rect	151	47	152	48
rect	151	53	152	54
rect	151	54	152	55
rect	151	56	152	57
rect	151	58	152	59
rect	151	59	152	60
rect	151	60	152	61
rect	151	66	152	67
rect	151	69	152	70
rect	151	72	152	73
rect	151	73	152	74
rect	151	78	152	79
rect	151	81	152	82
rect	151	83	152	84
rect	151	84	152	85
rect	151	87	152	88
rect	151	90	152	91
rect	151	94	152	95
rect	151	97	152	98
rect	151	100	152	101
rect	151	106	152	107
rect	151	110	152	111
rect	151	119	152	120
rect	151	126	152	127
rect	151	129	152	130
rect	151	135	152	136
rect	151	138	152	139
rect	151	145	152	146
rect	151	148	152	149
rect	151	151	152	152
rect	151	154	152	155
rect	151	157	152	158
rect	151	161	152	162
rect	151	164	152	165
rect	151	170	152	171
rect	151	173	152	174
rect	151	176	152	177
rect	151	179	152	180
rect	151	182	152	183
rect	151	186	152	187
rect	151	193	152	194
rect	152	1	153	2
rect	152	4	153	5
rect	152	7	153	8
rect	152	10	153	11
rect	152	13	153	14
rect	152	16	153	17
rect	152	17	153	18
rect	152	19	153	20
rect	152	20	153	21
rect	152	22	153	23
rect	152	23	153	24
rect	152	25	153	26
rect	152	26	153	27
rect	152	28	153	29
rect	152	31	153	32
rect	152	35	153	36
rect	152	41	153	42
rect	152	44	153	45
rect	152	47	153	48
rect	152	53	153	54
rect	152	54	153	55
rect	152	56	153	57
rect	152	58	153	59
rect	152	59	153	60
rect	152	60	153	61
rect	152	66	153	67
rect	152	69	153	70
rect	152	72	153	73
rect	152	73	153	74
rect	152	75	153	76
rect	152	78	153	79
rect	152	81	153	82
rect	152	83	153	84
rect	152	84	153	85
rect	152	87	153	88
rect	152	90	153	91
rect	152	94	153	95
rect	152	97	153	98
rect	152	100	153	101
rect	152	106	153	107
rect	152	110	153	111
rect	152	113	153	114
rect	152	119	153	120
rect	152	126	153	127
rect	152	129	153	130
rect	152	135	153	136
rect	152	138	153	139
rect	152	145	153	146
rect	152	148	153	149
rect	152	151	153	152
rect	152	154	153	155
rect	152	157	153	158
rect	152	161	153	162
rect	152	164	153	165
rect	152	170	153	171
rect	152	173	153	174
rect	152	176	153	177
rect	152	179	153	180
rect	152	182	153	183
rect	152	186	153	187
rect	152	193	153	194
rect	153	1	154	2
rect	153	4	154	5
rect	153	7	154	8
rect	153	10	154	11
rect	153	13	154	14
rect	153	16	154	17
rect	153	17	154	18
rect	153	19	154	20
rect	153	20	154	21
rect	153	22	154	23
rect	153	23	154	24
rect	153	25	154	26
rect	153	26	154	27
rect	153	28	154	29
rect	153	31	154	32
rect	153	35	154	36
rect	153	41	154	42
rect	153	44	154	45
rect	153	47	154	48
rect	153	53	154	54
rect	153	54	154	55
rect	153	56	154	57
rect	153	58	154	59
rect	153	59	154	60
rect	153	60	154	61
rect	153	66	154	67
rect	153	69	154	70
rect	153	72	154	73
rect	153	73	154	74
rect	153	75	154	76
rect	153	78	154	79
rect	153	81	154	82
rect	153	83	154	84
rect	153	87	154	88
rect	153	90	154	91
rect	153	94	154	95
rect	153	97	154	98
rect	153	106	154	107
rect	153	110	154	111
rect	153	113	154	114
rect	153	119	154	120
rect	153	126	154	127
rect	153	129	154	130
rect	153	135	154	136
rect	153	138	154	139
rect	153	145	154	146
rect	153	148	154	149
rect	153	151	154	152
rect	153	154	154	155
rect	153	157	154	158
rect	153	161	154	162
rect	153	164	154	165
rect	153	170	154	171
rect	153	173	154	174
rect	153	176	154	177
rect	153	179	154	180
rect	153	186	154	187
rect	153	193	154	194
rect	154	1	155	2
rect	154	4	155	5
rect	154	7	155	8
rect	154	10	155	11
rect	154	13	155	14
rect	154	16	155	17
rect	154	17	155	18
rect	154	19	155	20
rect	154	20	155	21
rect	154	22	155	23
rect	154	23	155	24
rect	154	25	155	26
rect	154	26	155	27
rect	154	28	155	29
rect	154	31	155	32
rect	154	35	155	36
rect	154	41	155	42
rect	154	44	155	45
rect	154	47	155	48
rect	154	53	155	54
rect	154	54	155	55
rect	154	56	155	57
rect	154	58	155	59
rect	154	59	155	60
rect	154	60	155	61
rect	154	62	155	63
rect	154	66	155	67
rect	154	69	155	70
rect	154	72	155	73
rect	154	73	155	74
rect	154	75	155	76
rect	154	78	155	79
rect	154	81	155	82
rect	154	83	155	84
rect	154	84	155	85
rect	154	87	155	88
rect	154	90	155	91
rect	154	94	155	95
rect	154	97	155	98
rect	154	106	155	107
rect	154	110	155	111
rect	154	113	155	114
rect	154	116	155	117
rect	154	119	155	120
rect	154	126	155	127
rect	154	129	155	130
rect	154	135	155	136
rect	154	138	155	139
rect	154	145	155	146
rect	154	148	155	149
rect	154	151	155	152
rect	154	154	155	155
rect	154	157	155	158
rect	154	161	155	162
rect	154	164	155	165
rect	154	167	155	168
rect	154	170	155	171
rect	154	173	155	174
rect	154	176	155	177
rect	154	179	155	180
rect	154	186	155	187
rect	154	193	155	194
rect	155	1	156	2
rect	155	4	156	5
rect	155	7	156	8
rect	155	10	156	11
rect	155	13	156	14
rect	155	16	156	17
rect	155	17	156	18
rect	155	19	156	20
rect	155	20	156	21
rect	155	22	156	23
rect	155	23	156	24
rect	155	25	156	26
rect	155	26	156	27
rect	155	28	156	29
rect	155	31	156	32
rect	155	35	156	36
rect	155	44	156	45
rect	155	47	156	48
rect	155	53	156	54
rect	155	54	156	55
rect	155	56	156	57
rect	155	58	156	59
rect	155	59	156	60
rect	155	60	156	61
rect	155	62	156	63
rect	155	66	156	67
rect	155	69	156	70
rect	155	73	156	74
rect	155	75	156	76
rect	155	78	156	79
rect	155	81	156	82
rect	155	83	156	84
rect	155	84	156	85
rect	155	87	156	88
rect	155	90	156	91
rect	155	97	156	98
rect	155	106	156	107
rect	155	110	156	111
rect	155	113	156	114
rect	155	116	156	117
rect	155	119	156	120
rect	155	126	156	127
rect	155	129	156	130
rect	155	138	156	139
rect	155	151	156	152
rect	155	154	156	155
rect	155	157	156	158
rect	155	161	156	162
rect	155	164	156	165
rect	155	167	156	168
rect	155	170	156	171
rect	155	173	156	174
rect	155	179	156	180
rect	155	186	156	187
rect	155	193	156	194
rect	156	1	157	2
rect	156	4	157	5
rect	156	7	157	8
rect	156	10	157	11
rect	156	13	157	14
rect	156	16	157	17
rect	156	17	157	18
rect	156	19	157	20
rect	156	20	157	21
rect	156	22	157	23
rect	156	23	157	24
rect	156	25	157	26
rect	156	26	157	27
rect	156	28	157	29
rect	156	31	157	32
rect	156	35	157	36
rect	156	44	157	45
rect	156	47	157	48
rect	156	53	157	54
rect	156	54	157	55
rect	156	56	157	57
rect	156	58	157	59
rect	156	59	157	60
rect	156	60	157	61
rect	156	62	157	63
rect	156	66	157	67
rect	156	69	157	70
rect	156	72	157	73
rect	156	73	157	74
rect	156	75	157	76
rect	156	78	157	79
rect	156	81	157	82
rect	156	83	157	84
rect	156	84	157	85
rect	156	87	157	88
rect	156	90	157	91
rect	156	97	157	98
rect	156	100	157	101
rect	156	106	157	107
rect	156	110	157	111
rect	156	113	157	114
rect	156	116	157	117
rect	156	119	157	120
rect	156	126	157	127
rect	156	129	157	130
rect	156	132	157	133
rect	156	138	157	139
rect	156	151	157	152
rect	156	154	157	155
rect	156	157	157	158
rect	156	161	157	162
rect	156	164	157	165
rect	156	167	157	168
rect	156	170	157	171
rect	156	173	157	174
rect	156	179	157	180
rect	156	183	157	184
rect	156	186	157	187
rect	156	193	157	194
rect	157	1	158	2
rect	157	4	158	5
rect	157	10	158	11
rect	157	13	158	14
rect	157	16	158	17
rect	157	17	158	18
rect	157	19	158	20
rect	157	20	158	21
rect	157	22	158	23
rect	157	23	158	24
rect	157	25	158	26
rect	157	26	158	27
rect	157	28	158	29
rect	157	31	158	32
rect	157	35	158	36
rect	157	44	158	45
rect	157	53	158	54
rect	157	54	158	55
rect	157	56	158	57
rect	157	58	158	59
rect	157	59	158	60
rect	157	60	158	61
rect	157	62	158	63
rect	157	66	158	67
rect	157	72	158	73
rect	157	73	158	74
rect	157	75	158	76
rect	157	78	158	79
rect	157	81	158	82
rect	157	83	158	84
rect	157	87	158	88
rect	157	90	158	91
rect	157	97	158	98
rect	157	100	158	101
rect	157	106	158	107
rect	157	110	158	111
rect	157	113	158	114
rect	157	116	158	117
rect	157	119	158	120
rect	157	126	158	127
rect	157	129	158	130
rect	157	132	158	133
rect	157	138	158	139
rect	157	151	158	152
rect	157	154	158	155
rect	157	157	158	158
rect	157	161	158	162
rect	157	164	158	165
rect	157	167	158	168
rect	157	170	158	171
rect	157	173	158	174
rect	157	179	158	180
rect	157	183	158	184
rect	157	186	158	187
rect	157	193	158	194
rect	158	1	159	2
rect	158	4	159	5
rect	158	10	159	11
rect	158	13	159	14
rect	158	16	159	17
rect	158	17	159	18
rect	158	19	159	20
rect	158	20	159	21
rect	158	22	159	23
rect	158	23	159	24
rect	158	25	159	26
rect	158	26	159	27
rect	158	28	159	29
rect	158	31	159	32
rect	158	35	159	36
rect	158	38	159	39
rect	158	44	159	45
rect	158	50	159	51
rect	158	53	159	54
rect	158	54	159	55
rect	158	56	159	57
rect	158	58	159	59
rect	158	59	159	60
rect	158	60	159	61
rect	158	62	159	63
rect	158	66	159	67
rect	158	72	159	73
rect	158	73	159	74
rect	158	75	159	76
rect	158	78	159	79
rect	158	81	159	82
rect	158	83	159	84
rect	158	84	159	85
rect	158	87	159	88
rect	158	90	159	91
rect	158	97	159	98
rect	158	100	159	101
rect	158	106	159	107
rect	158	110	159	111
rect	158	113	159	114
rect	158	116	159	117
rect	158	119	159	120
rect	158	126	159	127
rect	158	129	159	130
rect	158	132	159	133
rect	158	138	159	139
rect	158	151	159	152
rect	158	154	159	155
rect	158	157	159	158
rect	158	161	159	162
rect	158	164	159	165
rect	158	167	159	168
rect	158	170	159	171
rect	158	173	159	174
rect	158	177	159	178
rect	158	179	159	180
rect	158	183	159	184
rect	158	186	159	187
rect	158	193	159	194
rect	159	1	160	2
rect	159	4	160	5
rect	159	10	160	11
rect	159	13	160	14
rect	159	16	160	17
rect	159	17	160	18
rect	159	19	160	20
rect	159	20	160	21
rect	159	22	160	23
rect	159	23	160	24
rect	159	25	160	26
rect	159	26	160	27
rect	159	28	160	29
rect	159	35	160	36
rect	159	38	160	39
rect	159	44	160	45
rect	159	50	160	51
rect	159	53	160	54
rect	159	54	160	55
rect	159	56	160	57
rect	159	58	160	59
rect	159	59	160	60
rect	159	62	160	63
rect	159	66	160	67
rect	159	72	160	73
rect	159	73	160	74
rect	159	75	160	76
rect	159	78	160	79
rect	159	83	160	84
rect	159	84	160	85
rect	159	87	160	88
rect	159	90	160	91
rect	159	97	160	98
rect	159	100	160	101
rect	159	106	160	107
rect	159	110	160	111
rect	159	113	160	114
rect	159	116	160	117
rect	159	119	160	120
rect	159	126	160	127
rect	159	129	160	130
rect	159	132	160	133
rect	159	138	160	139
rect	159	151	160	152
rect	159	154	160	155
rect	159	157	160	158
rect	159	164	160	165
rect	159	167	160	168
rect	159	170	160	171
rect	159	173	160	174
rect	159	177	160	178
rect	159	179	160	180
rect	159	183	160	184
rect	159	186	160	187
rect	159	193	160	194
rect	160	1	161	2
rect	160	4	161	5
rect	160	7	161	8
rect	160	10	161	11
rect	160	13	161	14
rect	160	16	161	17
rect	160	17	161	18
rect	160	19	161	20
rect	160	20	161	21
rect	160	22	161	23
rect	160	23	161	24
rect	160	25	161	26
rect	160	26	161	27
rect	160	28	161	29
rect	160	35	161	36
rect	160	38	161	39
rect	160	41	161	42
rect	160	44	161	45
rect	160	47	161	48
rect	160	50	161	51
rect	160	53	161	54
rect	160	54	161	55
rect	160	56	161	57
rect	160	58	161	59
rect	160	59	161	60
rect	160	62	161	63
rect	160	66	161	67
rect	160	72	161	73
rect	160	73	161	74
rect	160	75	161	76
rect	160	78	161	79
rect	160	83	161	84
rect	160	84	161	85
rect	160	87	161	88
rect	160	90	161	91
rect	160	97	161	98
rect	160	100	161	101
rect	160	106	161	107
rect	160	110	161	111
rect	160	113	161	114
rect	160	116	161	117
rect	160	119	161	120
rect	160	126	161	127
rect	160	129	161	130
rect	160	132	161	133
rect	160	138	161	139
rect	160	151	161	152
rect	160	154	161	155
rect	160	157	161	158
rect	160	164	161	165
rect	160	167	161	168
rect	160	170	161	171
rect	160	173	161	174
rect	160	177	161	178
rect	160	179	161	180
rect	160	183	161	184
rect	160	186	161	187
rect	160	193	161	194
rect	161	1	162	2
rect	161	7	162	8
rect	161	16	162	17
rect	161	17	162	18
rect	161	19	162	20
rect	161	20	162	21
rect	161	22	162	23
rect	161	23	162	24
rect	161	25	162	26
rect	161	26	162	27
rect	161	28	162	29
rect	161	35	162	36
rect	161	38	162	39
rect	161	41	162	42
rect	161	44	162	45
rect	161	47	162	48
rect	161	50	162	51
rect	161	53	162	54
rect	161	54	162	55
rect	161	56	162	57
rect	161	58	162	59
rect	161	59	162	60
rect	161	62	162	63
rect	161	66	162	67
rect	161	72	162	73
rect	161	73	162	74
rect	161	75	162	76
rect	161	78	162	79
rect	161	83	162	84
rect	161	84	162	85
rect	161	87	162	88
rect	161	90	162	91
rect	161	97	162	98
rect	161	100	162	101
rect	161	106	162	107
rect	161	110	162	111
rect	161	113	162	114
rect	161	116	162	117
rect	161	119	162	120
rect	161	126	162	127
rect	161	129	162	130
rect	161	132	162	133
rect	161	154	162	155
rect	161	157	162	158
rect	161	164	162	165
rect	161	167	162	168
rect	161	170	162	171
rect	161	173	162	174
rect	161	177	162	178
rect	161	179	162	180
rect	161	183	162	184
rect	161	186	162	187
rect	161	193	162	194
rect	162	1	163	2
rect	162	7	163	8
rect	162	16	163	17
rect	162	17	163	18
rect	162	19	163	20
rect	162	20	163	21
rect	162	22	163	23
rect	162	23	163	24
rect	162	25	163	26
rect	162	26	163	27
rect	162	28	163	29
rect	162	32	163	33
rect	162	35	163	36
rect	162	38	163	39
rect	162	41	163	42
rect	162	44	163	45
rect	162	47	163	48
rect	162	50	163	51
rect	162	53	163	54
rect	162	54	163	55
rect	162	56	163	57
rect	162	58	163	59
rect	162	59	163	60
rect	162	62	163	63
rect	162	66	163	67
rect	162	72	163	73
rect	162	73	163	74
rect	162	75	163	76
rect	162	78	163	79
rect	162	83	163	84
rect	162	84	163	85
rect	162	87	163	88
rect	162	90	163	91
rect	162	97	163	98
rect	162	100	163	101
rect	162	103	163	104
rect	162	106	163	107
rect	162	110	163	111
rect	162	113	163	114
rect	162	116	163	117
rect	162	119	163	120
rect	162	126	163	127
rect	162	129	163	130
rect	162	132	163	133
rect	162	135	163	136
rect	162	148	163	149
rect	162	154	163	155
rect	162	157	163	158
rect	162	164	163	165
rect	162	167	163	168
rect	162	170	163	171
rect	162	173	163	174
rect	162	177	163	178
rect	162	179	163	180
rect	162	183	163	184
rect	162	186	163	187
rect	162	193	163	194
rect	163	1	164	2
rect	163	7	164	8
rect	163	16	164	17
rect	163	17	164	18
rect	163	19	164	20
rect	163	20	164	21
rect	163	22	164	23
rect	163	23	164	24
rect	163	25	164	26
rect	163	26	164	27
rect	163	32	164	33
rect	163	35	164	36
rect	163	38	164	39
rect	163	41	164	42
rect	163	44	164	45
rect	163	47	164	48
rect	163	50	164	51
rect	163	53	164	54
rect	163	54	164	55
rect	163	56	164	57
rect	163	58	164	59
rect	163	59	164	60
rect	163	62	164	63
rect	163	72	164	73
rect	163	73	164	74
rect	163	75	164	76
rect	163	78	164	79
rect	163	83	164	84
rect	163	84	164	85
rect	163	87	164	88
rect	163	90	164	91
rect	163	97	164	98
rect	163	100	164	101
rect	163	103	164	104
rect	163	106	164	107
rect	163	110	164	111
rect	163	113	164	114
rect	163	116	164	117
rect	163	119	164	120
rect	163	126	164	127
rect	163	129	164	130
rect	163	132	164	133
rect	163	135	164	136
rect	163	148	164	149
rect	163	154	164	155
rect	163	157	164	158
rect	163	164	164	165
rect	163	167	164	168
rect	163	170	164	171
rect	163	173	164	174
rect	163	177	164	178
rect	163	179	164	180
rect	163	183	164	184
rect	163	186	164	187
rect	164	1	165	2
rect	164	7	165	8
rect	164	10	165	11
rect	164	16	165	17
rect	164	17	165	18
rect	164	19	165	20
rect	164	20	165	21
rect	164	22	165	23
rect	164	23	165	24
rect	164	25	165	26
rect	164	26	165	27
rect	164	32	165	33
rect	164	35	165	36
rect	164	38	165	39
rect	164	41	165	42
rect	164	44	165	45
rect	164	47	165	48
rect	164	50	165	51
rect	164	53	165	54
rect	164	54	165	55
rect	164	56	165	57
rect	164	58	165	59
rect	164	59	165	60
rect	164	62	165	63
rect	164	72	165	73
rect	164	73	165	74
rect	164	75	165	76
rect	164	78	165	79
rect	164	81	165	82
rect	164	83	165	84
rect	164	84	165	85
rect	164	87	165	88
rect	164	90	165	91
rect	164	97	165	98
rect	164	100	165	101
rect	164	103	165	104
rect	164	106	165	107
rect	164	110	165	111
rect	164	113	165	114
rect	164	116	165	117
rect	164	119	165	120
rect	164	126	165	127
rect	164	129	165	130
rect	164	132	165	133
rect	164	135	165	136
rect	164	148	165	149
rect	164	154	165	155
rect	164	157	165	158
rect	164	164	165	165
rect	164	167	165	168
rect	164	170	165	171
rect	164	173	165	174
rect	164	177	165	178
rect	164	179	165	180
rect	164	183	165	184
rect	164	186	165	187
rect	165	1	166	2
rect	165	7	166	8
rect	165	10	166	11
rect	165	16	166	17
rect	165	17	166	18
rect	165	19	166	20
rect	165	20	166	21
rect	165	22	166	23
rect	165	23	166	24
rect	165	25	166	26
rect	165	26	166	27
rect	165	32	166	33
rect	165	35	166	36
rect	165	38	166	39
rect	165	41	166	42
rect	165	44	166	45
rect	165	47	166	48
rect	165	50	166	51
rect	165	53	166	54
rect	165	54	166	55
rect	165	56	166	57
rect	165	58	166	59
rect	165	59	166	60
rect	165	62	166	63
rect	165	72	166	73
rect	165	73	166	74
rect	165	75	166	76
rect	165	78	166	79
rect	165	81	166	82
rect	165	83	166	84
rect	165	84	166	85
rect	165	87	166	88
rect	165	90	166	91
rect	165	97	166	98
rect	165	100	166	101
rect	165	103	166	104
rect	165	106	166	107
rect	165	110	166	111
rect	165	113	166	114
rect	165	116	166	117
rect	165	119	166	120
rect	165	126	166	127
rect	165	129	166	130
rect	165	132	166	133
rect	165	135	166	136
rect	165	148	166	149
rect	165	157	166	158
rect	165	167	166	168
rect	165	173	166	174
rect	165	177	166	178
rect	165	179	166	180
rect	165	183	166	184
rect	166	1	167	2
rect	166	4	167	5
rect	166	7	167	8
rect	166	10	167	11
rect	166	16	167	17
rect	166	17	167	18
rect	166	19	167	20
rect	166	20	167	21
rect	166	22	167	23
rect	166	23	167	24
rect	166	25	167	26
rect	166	26	167	27
rect	166	32	167	33
rect	166	35	167	36
rect	166	38	167	39
rect	166	41	167	42
rect	166	44	167	45
rect	166	47	167	48
rect	166	50	167	51
rect	166	53	167	54
rect	166	54	167	55
rect	166	56	167	57
rect	166	58	167	59
rect	166	59	167	60
rect	166	62	167	63
rect	166	72	167	73
rect	166	73	167	74
rect	166	75	167	76
rect	166	78	167	79
rect	166	81	167	82
rect	166	83	167	84
rect	166	84	167	85
rect	166	87	167	88
rect	166	90	167	91
rect	166	97	167	98
rect	166	100	167	101
rect	166	103	167	104
rect	166	106	167	107
rect	166	110	167	111
rect	166	113	167	114
rect	166	116	167	117
rect	166	119	167	120
rect	166	126	167	127
rect	166	129	167	130
rect	166	132	167	133
rect	166	135	167	136
rect	166	148	167	149
rect	166	151	167	152
rect	166	157	167	158
rect	166	167	167	168
rect	166	173	167	174
rect	166	177	167	178
rect	166	179	167	180
rect	166	183	167	184
rect	167	4	168	5
rect	167	7	168	8
rect	167	10	168	11
rect	167	16	168	17
rect	167	17	168	18
rect	167	19	168	20
rect	167	20	168	21
rect	167	22	168	23
rect	167	23	168	24
rect	167	25	168	26
rect	167	26	168	27
rect	167	32	168	33
rect	167	35	168	36
rect	167	38	168	39
rect	167	41	168	42
rect	167	44	168	45
rect	167	47	168	48
rect	167	50	168	51
rect	167	53	168	54
rect	167	54	168	55
rect	167	56	168	57
rect	167	58	168	59
rect	167	59	168	60
rect	167	62	168	63
rect	167	72	168	73
rect	167	73	168	74
rect	167	75	168	76
rect	167	78	168	79
rect	167	81	168	82
rect	167	83	168	84
rect	167	84	168	85
rect	167	87	168	88
rect	167	90	168	91
rect	167	97	168	98
rect	167	100	168	101
rect	167	103	168	104
rect	167	106	168	107
rect	167	113	168	114
rect	167	116	168	117
rect	167	119	168	120
rect	167	129	168	130
rect	167	132	168	133
rect	167	135	168	136
rect	167	148	168	149
rect	167	151	168	152
rect	167	157	168	158
rect	167	167	168	168
rect	167	173	168	174
rect	167	177	168	178
rect	167	183	168	184
rect	168	4	169	5
rect	168	7	169	8
rect	168	10	169	11
rect	168	16	169	17
rect	168	17	169	18
rect	168	19	169	20
rect	168	20	169	21
rect	168	22	169	23
rect	168	23	169	24
rect	168	25	169	26
rect	168	26	169	27
rect	168	32	169	33
rect	168	35	169	36
rect	168	38	169	39
rect	168	41	169	42
rect	168	44	169	45
rect	168	47	169	48
rect	168	50	169	51
rect	168	53	169	54
rect	168	54	169	55
rect	168	56	169	57
rect	168	58	169	59
rect	168	59	169	60
rect	168	62	169	63
rect	168	72	169	73
rect	168	73	169	74
rect	168	75	169	76
rect	168	78	169	79
rect	168	81	169	82
rect	168	83	169	84
rect	168	84	169	85
rect	168	87	169	88
rect	168	90	169	91
rect	168	97	169	98
rect	168	100	169	101
rect	168	103	169	104
rect	168	106	169	107
rect	168	113	169	114
rect	168	116	169	117
rect	168	119	169	120
rect	168	129	169	130
rect	168	132	169	133
rect	168	135	169	136
rect	168	145	169	146
rect	168	148	169	149
rect	168	151	169	152
rect	168	154	169	155
rect	168	157	169	158
rect	168	167	169	168
rect	168	173	169	174
rect	168	177	169	178
rect	168	183	169	184
rect	169	4	170	5
rect	169	7	170	8
rect	169	10	170	11
rect	169	16	170	17
rect	169	17	170	18
rect	169	19	170	20
rect	169	20	170	21
rect	169	23	170	24
rect	169	25	170	26
rect	169	26	170	27
rect	169	32	170	33
rect	169	35	170	36
rect	169	38	170	39
rect	169	41	170	42
rect	169	44	170	45
rect	169	47	170	48
rect	169	50	170	51
rect	169	53	170	54
rect	169	54	170	55
rect	169	56	170	57
rect	169	58	170	59
rect	169	59	170	60
rect	169	62	170	63
rect	169	72	170	73
rect	169	73	170	74
rect	169	75	170	76
rect	169	78	170	79
rect	169	81	170	82
rect	169	83	170	84
rect	169	84	170	85
rect	169	87	170	88
rect	169	90	170	91
rect	169	97	170	98
rect	169	100	170	101
rect	169	103	170	104
rect	169	106	170	107
rect	169	113	170	114
rect	169	116	170	117
rect	169	119	170	120
rect	169	129	170	130
rect	169	132	170	133
rect	169	135	170	136
rect	169	145	170	146
rect	169	148	170	149
rect	169	151	170	152
rect	169	154	170	155
rect	169	157	170	158
rect	169	167	170	168
rect	169	177	170	178
rect	169	183	170	184
rect	170	1	171	2
rect	170	4	171	5
rect	170	7	171	8
rect	170	10	171	11
rect	170	13	171	14
rect	170	16	171	17
rect	170	17	171	18
rect	170	19	171	20
rect	170	20	171	21
rect	170	22	171	23
rect	170	23	171	24
rect	170	25	171	26
rect	170	26	171	27
rect	170	32	171	33
rect	170	35	171	36
rect	170	38	171	39
rect	170	41	171	42
rect	170	44	171	45
rect	170	47	171	48
rect	170	50	171	51
rect	170	53	171	54
rect	170	54	171	55
rect	170	56	171	57
rect	170	58	171	59
rect	170	59	171	60
rect	170	62	171	63
rect	170	72	171	73
rect	170	73	171	74
rect	170	75	171	76
rect	170	78	171	79
rect	170	81	171	82
rect	170	83	171	84
rect	170	84	171	85
rect	170	87	171	88
rect	170	90	171	91
rect	170	97	171	98
rect	170	100	171	101
rect	170	103	171	104
rect	170	106	171	107
rect	170	113	171	114
rect	170	116	171	117
rect	170	119	171	120
rect	170	123	171	124
rect	170	126	171	127
rect	170	129	171	130
rect	170	132	171	133
rect	170	135	171	136
rect	170	145	171	146
rect	170	148	171	149
rect	170	151	171	152
rect	170	154	171	155
rect	170	157	171	158
rect	170	167	171	168
rect	170	170	171	171
rect	170	177	171	178
rect	170	180	171	181
rect	170	183	171	184
rect	171	16	172	17
rect	171	17	172	18
rect	171	19	172	20
rect	171	20	172	21
rect	171	22	172	23
rect	171	23	172	24
rect	171	26	172	27
rect	171	53	172	54
rect	171	54	172	55
rect	171	58	172	59
rect	171	59	172	60
rect	171	72	172	73
rect	171	73	172	74
rect	171	83	172	84
rect	171	84	172	85
rect	172	16	173	17
rect	172	17	173	18
rect	172	19	173	20
rect	172	20	173	21
rect	172	22	173	23
rect	172	23	173	24
rect	172	26	173	27
rect	172	53	173	54
rect	172	54	173	55
rect	172	58	173	59
rect	172	59	173	60
rect	172	72	173	73
rect	172	73	173	74
rect	172	83	173	84
rect	172	84	173	85
rect	173	16	174	17
rect	173	17	174	18
rect	173	19	174	20
rect	173	20	174	21
rect	173	22	174	23
rect	173	23	174	24
rect	173	26	174	27
rect	173	53	174	54
rect	173	54	174	55
rect	173	58	174	59
rect	173	59	174	60
rect	173	72	174	73
rect	173	73	174	74
rect	173	83	174	84
rect	173	84	174	85
rect	174	16	175	17
rect	174	17	175	18
rect	174	19	175	20
rect	174	20	175	21
rect	174	22	175	23
rect	174	23	175	24
rect	174	26	175	27
rect	174	53	175	54
rect	174	54	175	55
rect	174	58	175	59
rect	174	59	175	60
rect	174	72	175	73
rect	174	73	175	74
rect	174	83	175	84
rect	174	84	175	85
rect	175	16	176	17
rect	175	17	176	18
rect	175	19	176	20
rect	175	20	176	21
rect	175	22	176	23
rect	175	23	176	24
rect	175	26	176	27
rect	175	53	176	54
rect	175	54	176	55
rect	175	58	176	59
rect	175	59	176	60
rect	175	72	176	73
rect	175	73	176	74
rect	175	83	176	84
rect	175	84	176	85
rect	176	17	177	18
rect	176	20	177	21
rect	176	23	177	24
rect	176	26	177	27
rect	176	54	177	55
rect	176	58	177	59
rect	176	73	177	74
rect	176	83	177	84
rect	177	1	178	2
rect	177	7	178	8
rect	177	10	178	11
rect	177	13	178	14
rect	177	17	178	18
rect	177	20	178	21
rect	177	23	178	24
rect	177	25	178	26
rect	177	26	178	27
rect	177	29	178	30
rect	177	32	178	33
rect	177	35	178	36
rect	177	38	178	39
rect	177	41	178	42
rect	177	44	178	45
rect	177	47	178	48
rect	177	50	178	51
rect	177	54	178	55
rect	177	56	178	57
rect	177	58	178	59
rect	177	62	178	63
rect	177	69	178	70
rect	177	73	178	74
rect	177	75	178	76
rect	177	78	178	79
rect	177	81	178	82
rect	177	83	178	84
rect	177	87	178	88
rect	177	90	178	91
rect	177	94	178	95
rect	177	100	178	101
rect	177	103	178	104
rect	177	106	178	107
rect	177	116	178	117
rect	177	119	178	120
rect	177	123	178	124
rect	177	129	178	130
rect	177	132	178	133
rect	177	135	178	136
rect	177	145	178	146
rect	177	148	178	149
rect	177	151	178	152
rect	177	154	178	155
rect	177	157	178	158
rect	177	164	178	165
rect	177	167	178	168
rect	177	170	178	171
rect	177	180	178	181
rect	177	183	178	184
rect	177	187	178	188
rect	177	190	178	191
rect	178	1	179	2
rect	178	7	179	8
rect	178	10	179	11
rect	178	13	179	14
rect	178	17	179	18
rect	178	20	179	21
rect	178	23	179	24
rect	178	25	179	26
rect	178	26	179	27
rect	178	29	179	30
rect	178	32	179	33
rect	178	35	179	36
rect	178	38	179	39
rect	178	41	179	42
rect	178	44	179	45
rect	178	47	179	48
rect	178	50	179	51
rect	178	54	179	55
rect	178	56	179	57
rect	178	58	179	59
rect	178	62	179	63
rect	178	69	179	70
rect	178	73	179	74
rect	178	75	179	76
rect	178	78	179	79
rect	178	81	179	82
rect	178	83	179	84
rect	178	87	179	88
rect	178	90	179	91
rect	178	94	179	95
rect	178	100	179	101
rect	178	103	179	104
rect	178	106	179	107
rect	178	116	179	117
rect	178	119	179	120
rect	178	123	179	124
rect	178	129	179	130
rect	178	132	179	133
rect	178	135	179	136
rect	178	145	179	146
rect	178	148	179	149
rect	178	151	179	152
rect	178	154	179	155
rect	178	157	179	158
rect	178	164	179	165
rect	178	167	179	168
rect	178	170	179	171
rect	178	180	179	181
rect	178	183	179	184
rect	178	187	179	188
rect	178	190	179	191
rect	179	1	180	2
rect	179	7	180	8
rect	179	10	180	11
rect	179	13	180	14
rect	179	17	180	18
rect	179	20	180	21
rect	179	23	180	24
rect	179	25	180	26
rect	179	26	180	27
rect	179	29	180	30
rect	179	32	180	33
rect	179	35	180	36
rect	179	38	180	39
rect	179	41	180	42
rect	179	44	180	45
rect	179	47	180	48
rect	179	50	180	51
rect	179	54	180	55
rect	179	56	180	57
rect	179	58	180	59
rect	179	62	180	63
rect	179	69	180	70
rect	179	73	180	74
rect	179	75	180	76
rect	179	78	180	79
rect	179	81	180	82
rect	179	83	180	84
rect	179	87	180	88
rect	179	90	180	91
rect	179	94	180	95
rect	179	100	180	101
rect	179	103	180	104
rect	179	106	180	107
rect	179	116	180	117
rect	179	119	180	120
rect	179	123	180	124
rect	179	129	180	130
rect	179	132	180	133
rect	179	135	180	136
rect	179	145	180	146
rect	179	148	180	149
rect	179	151	180	152
rect	179	154	180	155
rect	179	157	180	158
rect	179	164	180	165
rect	179	167	180	168
rect	179	170	180	171
rect	179	180	180	181
rect	179	183	180	184
rect	179	187	180	188
rect	179	190	180	191
rect	180	1	181	2
rect	180	7	181	8
rect	180	10	181	11
rect	180	13	181	14
rect	180	17	181	18
rect	180	20	181	21
rect	180	23	181	24
rect	180	25	181	26
rect	180	26	181	27
rect	180	29	181	30
rect	180	32	181	33
rect	180	35	181	36
rect	180	38	181	39
rect	180	41	181	42
rect	180	44	181	45
rect	180	47	181	48
rect	180	50	181	51
rect	180	54	181	55
rect	180	56	181	57
rect	180	58	181	59
rect	180	62	181	63
rect	180	69	181	70
rect	180	73	181	74
rect	180	75	181	76
rect	180	78	181	79
rect	180	81	181	82
rect	180	83	181	84
rect	180	87	181	88
rect	180	90	181	91
rect	180	94	181	95
rect	180	100	181	101
rect	180	103	181	104
rect	180	106	181	107
rect	180	116	181	117
rect	180	119	181	120
rect	180	123	181	124
rect	180	129	181	130
rect	180	132	181	133
rect	180	135	181	136
rect	180	145	181	146
rect	180	148	181	149
rect	180	151	181	152
rect	180	154	181	155
rect	180	157	181	158
rect	180	164	181	165
rect	180	167	181	168
rect	180	170	181	171
rect	180	180	181	181
rect	180	183	181	184
rect	180	187	181	188
rect	180	190	181	191
rect	181	1	182	2
rect	181	7	182	8
rect	181	10	182	11
rect	181	13	182	14
rect	181	17	182	18
rect	181	20	182	21
rect	181	23	182	24
rect	181	25	182	26
rect	181	26	182	27
rect	181	29	182	30
rect	181	32	182	33
rect	181	35	182	36
rect	181	38	182	39
rect	181	41	182	42
rect	181	44	182	45
rect	181	47	182	48
rect	181	50	182	51
rect	181	54	182	55
rect	181	56	182	57
rect	181	58	182	59
rect	181	62	182	63
rect	181	69	182	70
rect	181	73	182	74
rect	181	75	182	76
rect	181	78	182	79
rect	181	81	182	82
rect	181	83	182	84
rect	181	87	182	88
rect	181	90	182	91
rect	181	94	182	95
rect	181	100	182	101
rect	181	103	182	104
rect	181	106	182	107
rect	181	116	182	117
rect	181	119	182	120
rect	181	123	182	124
rect	181	129	182	130
rect	181	132	182	133
rect	181	135	182	136
rect	181	145	182	146
rect	181	148	182	149
rect	181	151	182	152
rect	181	154	182	155
rect	181	157	182	158
rect	181	164	182	165
rect	181	167	182	168
rect	181	170	182	171
rect	181	180	182	181
rect	181	183	182	184
rect	181	187	182	188
rect	181	190	182	191
rect	182	1	183	2
rect	182	7	183	8
rect	182	10	183	11
rect	182	13	183	14
rect	182	17	183	18
rect	182	20	183	21
rect	182	23	183	24
rect	182	25	183	26
rect	182	26	183	27
rect	182	29	183	30
rect	182	32	183	33
rect	182	35	183	36
rect	182	38	183	39
rect	182	41	183	42
rect	182	44	183	45
rect	182	47	183	48
rect	182	50	183	51
rect	182	54	183	55
rect	182	56	183	57
rect	182	58	183	59
rect	182	62	183	63
rect	182	69	183	70
rect	182	73	183	74
rect	182	75	183	76
rect	182	78	183	79
rect	182	81	183	82
rect	182	83	183	84
rect	182	87	183	88
rect	182	90	183	91
rect	182	94	183	95
rect	182	100	183	101
rect	182	103	183	104
rect	182	106	183	107
rect	182	116	183	117
rect	182	119	183	120
rect	182	123	183	124
rect	182	129	183	130
rect	182	132	183	133
rect	182	135	183	136
rect	182	145	183	146
rect	182	148	183	149
rect	182	151	183	152
rect	182	154	183	155
rect	182	157	183	158
rect	182	164	183	165
rect	182	167	183	168
rect	182	170	183	171
rect	182	180	183	181
rect	182	183	183	184
rect	182	187	183	188
rect	182	190	183	191
rect	183	1	184	2
rect	183	7	184	8
rect	183	10	184	11
rect	183	13	184	14
rect	183	17	184	18
rect	183	20	184	21
rect	183	23	184	24
rect	183	25	184	26
rect	183	26	184	27
rect	183	29	184	30
rect	183	32	184	33
rect	183	35	184	36
rect	183	38	184	39
rect	183	41	184	42
rect	183	44	184	45
rect	183	47	184	48
rect	183	50	184	51
rect	183	54	184	55
rect	183	56	184	57
rect	183	58	184	59
rect	183	62	184	63
rect	183	69	184	70
rect	183	73	184	74
rect	183	75	184	76
rect	183	78	184	79
rect	183	81	184	82
rect	183	83	184	84
rect	183	87	184	88
rect	183	90	184	91
rect	183	94	184	95
rect	183	100	184	101
rect	183	103	184	104
rect	183	106	184	107
rect	183	116	184	117
rect	183	119	184	120
rect	183	123	184	124
rect	183	129	184	130
rect	183	132	184	133
rect	183	135	184	136
rect	183	145	184	146
rect	183	148	184	149
rect	183	151	184	152
rect	183	154	184	155
rect	183	157	184	158
rect	183	164	184	165
rect	183	167	184	168
rect	183	170	184	171
rect	183	180	184	181
rect	183	183	184	184
rect	183	187	184	188
rect	183	190	184	191
rect	184	1	185	2
rect	184	7	185	8
rect	184	10	185	11
rect	184	13	185	14
rect	184	17	185	18
rect	184	20	185	21
rect	184	23	185	24
rect	184	25	185	26
rect	184	26	185	27
rect	184	29	185	30
rect	184	32	185	33
rect	184	35	185	36
rect	184	38	185	39
rect	184	41	185	42
rect	184	44	185	45
rect	184	47	185	48
rect	184	50	185	51
rect	184	54	185	55
rect	184	56	185	57
rect	184	58	185	59
rect	184	62	185	63
rect	184	69	185	70
rect	184	73	185	74
rect	184	75	185	76
rect	184	78	185	79
rect	184	81	185	82
rect	184	83	185	84
rect	184	87	185	88
rect	184	90	185	91
rect	184	94	185	95
rect	184	100	185	101
rect	184	103	185	104
rect	184	106	185	107
rect	184	116	185	117
rect	184	119	185	120
rect	184	123	185	124
rect	184	129	185	130
rect	184	132	185	133
rect	184	135	185	136
rect	184	145	185	146
rect	184	148	185	149
rect	184	151	185	152
rect	184	154	185	155
rect	184	157	185	158
rect	184	164	185	165
rect	184	167	185	168
rect	184	170	185	171
rect	184	180	185	181
rect	184	183	185	184
rect	184	187	185	188
rect	184	190	185	191
rect	185	1	186	2
rect	185	7	186	8
rect	185	10	186	11
rect	185	13	186	14
rect	185	17	186	18
rect	185	20	186	21
rect	185	23	186	24
rect	185	25	186	26
rect	185	26	186	27
rect	185	29	186	30
rect	185	32	186	33
rect	185	35	186	36
rect	185	38	186	39
rect	185	41	186	42
rect	185	44	186	45
rect	185	47	186	48
rect	185	50	186	51
rect	185	54	186	55
rect	185	56	186	57
rect	185	58	186	59
rect	185	62	186	63
rect	185	69	186	70
rect	185	73	186	74
rect	185	75	186	76
rect	185	78	186	79
rect	185	81	186	82
rect	185	83	186	84
rect	185	87	186	88
rect	185	90	186	91
rect	185	94	186	95
rect	185	100	186	101
rect	185	103	186	104
rect	185	106	186	107
rect	185	116	186	117
rect	185	119	186	120
rect	185	123	186	124
rect	185	129	186	130
rect	185	132	186	133
rect	185	135	186	136
rect	185	145	186	146
rect	185	148	186	149
rect	185	151	186	152
rect	185	154	186	155
rect	185	157	186	158
rect	185	164	186	165
rect	185	167	186	168
rect	185	170	186	171
rect	185	180	186	181
rect	185	183	186	184
rect	185	187	186	188
rect	185	190	186	191
rect	186	1	187	2
rect	186	7	187	8
rect	186	10	187	11
rect	186	13	187	14
rect	186	17	187	18
rect	186	20	187	21
rect	186	23	187	24
rect	186	25	187	26
rect	186	26	187	27
rect	186	29	187	30
rect	186	32	187	33
rect	186	35	187	36
rect	186	38	187	39
rect	186	41	187	42
rect	186	44	187	45
rect	186	47	187	48
rect	186	50	187	51
rect	186	54	187	55
rect	186	56	187	57
rect	186	58	187	59
rect	186	62	187	63
rect	186	69	187	70
rect	186	73	187	74
rect	186	75	187	76
rect	186	78	187	79
rect	186	81	187	82
rect	186	83	187	84
rect	186	87	187	88
rect	186	90	187	91
rect	186	94	187	95
rect	186	100	187	101
rect	186	103	187	104
rect	186	106	187	107
rect	186	116	187	117
rect	186	119	187	120
rect	186	123	187	124
rect	186	129	187	130
rect	186	132	187	133
rect	186	135	187	136
rect	186	145	187	146
rect	186	148	187	149
rect	186	151	187	152
rect	186	154	187	155
rect	186	157	187	158
rect	186	164	187	165
rect	186	167	187	168
rect	186	170	187	171
rect	186	180	187	181
rect	186	183	187	184
rect	186	187	187	188
rect	186	190	187	191
rect	187	1	188	2
rect	187	7	188	8
rect	187	10	188	11
rect	187	13	188	14
rect	187	17	188	18
rect	187	20	188	21
rect	187	23	188	24
rect	187	25	188	26
rect	187	26	188	27
rect	187	29	188	30
rect	187	32	188	33
rect	187	35	188	36
rect	187	38	188	39
rect	187	41	188	42
rect	187	44	188	45
rect	187	47	188	48
rect	187	50	188	51
rect	187	54	188	55
rect	187	56	188	57
rect	187	58	188	59
rect	187	62	188	63
rect	187	69	188	70
rect	187	73	188	74
rect	187	75	188	76
rect	187	78	188	79
rect	187	81	188	82
rect	187	83	188	84
rect	187	87	188	88
rect	187	90	188	91
rect	187	94	188	95
rect	187	100	188	101
rect	187	103	188	104
rect	187	106	188	107
rect	187	116	188	117
rect	187	119	188	120
rect	187	123	188	124
rect	187	129	188	130
rect	187	132	188	133
rect	187	135	188	136
rect	187	145	188	146
rect	187	148	188	149
rect	187	151	188	152
rect	187	154	188	155
rect	187	157	188	158
rect	187	164	188	165
rect	187	167	188	168
rect	187	170	188	171
rect	187	180	188	181
rect	187	183	188	184
rect	187	187	188	188
rect	187	190	188	191
rect	188	1	189	2
rect	188	7	189	8
rect	188	10	189	11
rect	188	13	189	14
rect	188	17	189	18
rect	188	20	189	21
rect	188	23	189	24
rect	188	25	189	26
rect	188	26	189	27
rect	188	29	189	30
rect	188	32	189	33
rect	188	35	189	36
rect	188	38	189	39
rect	188	41	189	42
rect	188	44	189	45
rect	188	47	189	48
rect	188	50	189	51
rect	188	54	189	55
rect	188	56	189	57
rect	188	58	189	59
rect	188	62	189	63
rect	188	69	189	70
rect	188	73	189	74
rect	188	75	189	76
rect	188	78	189	79
rect	188	81	189	82
rect	188	83	189	84
rect	188	87	189	88
rect	188	90	189	91
rect	188	94	189	95
rect	188	100	189	101
rect	188	103	189	104
rect	188	106	189	107
rect	188	116	189	117
rect	188	119	189	120
rect	188	123	189	124
rect	188	129	189	130
rect	188	132	189	133
rect	188	135	189	136
rect	188	145	189	146
rect	188	148	189	149
rect	188	151	189	152
rect	188	154	189	155
rect	188	157	189	158
rect	188	164	189	165
rect	188	167	189	168
rect	188	170	189	171
rect	188	180	189	181
rect	188	183	189	184
rect	188	187	189	188
rect	188	190	189	191
rect	189	1	190	2
rect	189	7	190	8
rect	189	10	190	11
rect	189	13	190	14
rect	189	17	190	18
rect	189	20	190	21
rect	189	23	190	24
rect	189	25	190	26
rect	189	26	190	27
rect	189	29	190	30
rect	189	32	190	33
rect	189	35	190	36
rect	189	38	190	39
rect	189	41	190	42
rect	189	44	190	45
rect	189	47	190	48
rect	189	50	190	51
rect	189	54	190	55
rect	189	56	190	57
rect	189	58	190	59
rect	189	62	190	63
rect	189	69	190	70
rect	189	73	190	74
rect	189	75	190	76
rect	189	78	190	79
rect	189	81	190	82
rect	189	83	190	84
rect	189	87	190	88
rect	189	90	190	91
rect	189	94	190	95
rect	189	100	190	101
rect	189	103	190	104
rect	189	106	190	107
rect	189	116	190	117
rect	189	119	190	120
rect	189	123	190	124
rect	189	129	190	130
rect	189	132	190	133
rect	189	135	190	136
rect	189	145	190	146
rect	189	148	190	149
rect	189	151	190	152
rect	189	154	190	155
rect	189	157	190	158
rect	189	164	190	165
rect	189	167	190	168
rect	189	170	190	171
rect	189	180	190	181
rect	189	183	190	184
rect	189	187	190	188
rect	189	190	190	191
rect	190	1	191	2
rect	190	7	191	8
rect	190	10	191	11
rect	190	13	191	14
rect	190	17	191	18
rect	190	20	191	21
rect	190	23	191	24
rect	190	25	191	26
rect	190	26	191	27
rect	190	29	191	30
rect	190	32	191	33
rect	190	35	191	36
rect	190	38	191	39
rect	190	41	191	42
rect	190	44	191	45
rect	190	47	191	48
rect	190	50	191	51
rect	190	54	191	55
rect	190	56	191	57
rect	190	58	191	59
rect	190	62	191	63
rect	190	69	191	70
rect	190	73	191	74
rect	190	75	191	76
rect	190	78	191	79
rect	190	81	191	82
rect	190	83	191	84
rect	190	87	191	88
rect	190	90	191	91
rect	190	94	191	95
rect	190	100	191	101
rect	190	103	191	104
rect	190	106	191	107
rect	190	116	191	117
rect	190	119	191	120
rect	190	123	191	124
rect	190	129	191	130
rect	190	132	191	133
rect	190	135	191	136
rect	190	145	191	146
rect	190	148	191	149
rect	190	151	191	152
rect	190	154	191	155
rect	190	157	191	158
rect	190	164	191	165
rect	190	167	191	168
rect	190	170	191	171
rect	190	180	191	181
rect	190	183	191	184
rect	190	187	191	188
rect	190	190	191	191
rect	191	1	192	2
rect	191	7	192	8
rect	191	10	192	11
rect	191	13	192	14
rect	191	17	192	18
rect	191	20	192	21
rect	191	23	192	24
rect	191	25	192	26
rect	191	26	192	27
rect	191	29	192	30
rect	191	32	192	33
rect	191	35	192	36
rect	191	38	192	39
rect	191	41	192	42
rect	191	44	192	45
rect	191	47	192	48
rect	191	50	192	51
rect	191	54	192	55
rect	191	56	192	57
rect	191	58	192	59
rect	191	62	192	63
rect	191	69	192	70
rect	191	73	192	74
rect	191	75	192	76
rect	191	78	192	79
rect	191	81	192	82
rect	191	83	192	84
rect	191	87	192	88
rect	191	90	192	91
rect	191	94	192	95
rect	191	100	192	101
rect	191	103	192	104
rect	191	106	192	107
rect	191	116	192	117
rect	191	119	192	120
rect	191	123	192	124
rect	191	129	192	130
rect	191	132	192	133
rect	191	135	192	136
rect	191	145	192	146
rect	191	148	192	149
rect	191	151	192	152
rect	191	154	192	155
rect	191	157	192	158
rect	191	164	192	165
rect	191	167	192	168
rect	191	170	192	171
rect	191	180	192	181
rect	191	183	192	184
rect	191	187	192	188
rect	191	190	192	191
rect	192	1	193	2
rect	192	7	193	8
rect	192	10	193	11
rect	192	13	193	14
rect	192	17	193	18
rect	192	20	193	21
rect	192	23	193	24
rect	192	25	193	26
rect	192	26	193	27
rect	192	29	193	30
rect	192	32	193	33
rect	192	35	193	36
rect	192	38	193	39
rect	192	41	193	42
rect	192	44	193	45
rect	192	47	193	48
rect	192	50	193	51
rect	192	54	193	55
rect	192	56	193	57
rect	192	58	193	59
rect	192	62	193	63
rect	192	69	193	70
rect	192	73	193	74
rect	192	75	193	76
rect	192	78	193	79
rect	192	81	193	82
rect	192	83	193	84
rect	192	87	193	88
rect	192	90	193	91
rect	192	94	193	95
rect	192	100	193	101
rect	192	103	193	104
rect	192	106	193	107
rect	192	116	193	117
rect	192	119	193	120
rect	192	123	193	124
rect	192	129	193	130
rect	192	132	193	133
rect	192	135	193	136
rect	192	145	193	146
rect	192	148	193	149
rect	192	151	193	152
rect	192	154	193	155
rect	192	157	193	158
rect	192	164	193	165
rect	192	167	193	168
rect	192	170	193	171
rect	192	180	193	181
rect	192	183	193	184
rect	192	187	193	188
rect	192	190	193	191
rect	193	1	194	2
rect	193	7	194	8
rect	193	10	194	11
rect	193	13	194	14
rect	193	17	194	18
rect	193	20	194	21
rect	193	23	194	24
rect	193	25	194	26
rect	193	26	194	27
rect	193	29	194	30
rect	193	32	194	33
rect	193	35	194	36
rect	193	38	194	39
rect	193	41	194	42
rect	193	44	194	45
rect	193	47	194	48
rect	193	50	194	51
rect	193	54	194	55
rect	193	56	194	57
rect	193	58	194	59
rect	193	62	194	63
rect	193	69	194	70
rect	193	73	194	74
rect	193	75	194	76
rect	193	78	194	79
rect	193	81	194	82
rect	193	83	194	84
rect	193	87	194	88
rect	193	90	194	91
rect	193	94	194	95
rect	193	100	194	101
rect	193	103	194	104
rect	193	106	194	107
rect	193	116	194	117
rect	193	119	194	120
rect	193	123	194	124
rect	193	129	194	130
rect	193	132	194	133
rect	193	135	194	136
rect	193	145	194	146
rect	193	148	194	149
rect	193	151	194	152
rect	193	154	194	155
rect	193	157	194	158
rect	193	164	194	165
rect	193	167	194	168
rect	193	170	194	171
rect	193	180	194	181
rect	193	183	194	184
rect	193	187	194	188
rect	193	190	194	191
rect	194	1	195	2
rect	194	7	195	8
rect	194	10	195	11
rect	194	13	195	14
rect	194	17	195	18
rect	194	20	195	21
rect	194	23	195	24
rect	194	25	195	26
rect	194	26	195	27
rect	194	29	195	30
rect	194	32	195	33
rect	194	35	195	36
rect	194	38	195	39
rect	194	41	195	42
rect	194	44	195	45
rect	194	47	195	48
rect	194	50	195	51
rect	194	54	195	55
rect	194	56	195	57
rect	194	58	195	59
rect	194	62	195	63
rect	194	69	195	70
rect	194	73	195	74
rect	194	78	195	79
rect	194	81	195	82
rect	194	83	195	84
rect	194	87	195	88
rect	194	90	195	91
rect	194	94	195	95
rect	194	100	195	101
rect	194	103	195	104
rect	194	106	195	107
rect	194	116	195	117
rect	194	119	195	120
rect	194	123	195	124
rect	194	129	195	130
rect	194	132	195	133
rect	194	135	195	136
rect	194	145	195	146
rect	194	148	195	149
rect	194	151	195	152
rect	194	154	195	155
rect	194	157	195	158
rect	194	164	195	165
rect	194	167	195	168
rect	194	170	195	171
rect	194	180	195	181
rect	194	183	195	184
rect	194	187	195	188
rect	194	190	195	191
rect	195	1	196	2
rect	195	7	196	8
rect	195	10	196	11
rect	195	13	196	14
rect	195	17	196	18
rect	195	20	196	21
rect	195	23	196	24
rect	195	25	196	26
rect	195	26	196	27
rect	195	29	196	30
rect	195	32	196	33
rect	195	35	196	36
rect	195	38	196	39
rect	195	41	196	42
rect	195	44	196	45
rect	195	47	196	48
rect	195	50	196	51
rect	195	54	196	55
rect	195	56	196	57
rect	195	58	196	59
rect	195	62	196	63
rect	195	64	196	65
rect	195	69	196	70
rect	195	73	196	74
rect	195	78	196	79
rect	195	81	196	82
rect	195	83	196	84
rect	195	87	196	88
rect	195	90	196	91
rect	195	94	196	95
rect	195	100	196	101
rect	195	103	196	104
rect	195	106	196	107
rect	195	116	196	117
rect	195	119	196	120
rect	195	123	196	124
rect	195	129	196	130
rect	195	132	196	133
rect	195	135	196	136
rect	195	145	196	146
rect	195	148	196	149
rect	195	151	196	152
rect	195	154	196	155
rect	195	157	196	158
rect	195	164	196	165
rect	195	167	196	168
rect	195	170	196	171
rect	195	180	196	181
rect	195	183	196	184
rect	195	187	196	188
rect	195	190	196	191
rect	196	1	197	2
rect	196	7	197	8
rect	196	10	197	11
rect	196	13	197	14
rect	196	17	197	18
rect	196	20	197	21
rect	196	23	197	24
rect	196	25	197	26
rect	196	26	197	27
rect	196	29	197	30
rect	196	32	197	33
rect	196	35	197	36
rect	196	38	197	39
rect	196	41	197	42
rect	196	44	197	45
rect	196	47	197	48
rect	196	50	197	51
rect	196	54	197	55
rect	196	56	197	57
rect	196	58	197	59
rect	196	62	197	63
rect	196	64	197	65
rect	196	69	197	70
rect	196	73	197	74
rect	196	78	197	79
rect	196	81	197	82
rect	196	83	197	84
rect	196	87	197	88
rect	196	94	197	95
rect	196	100	197	101
rect	196	103	197	104
rect	196	106	197	107
rect	196	116	197	117
rect	196	119	197	120
rect	196	123	197	124
rect	196	129	197	130
rect	196	132	197	133
rect	196	135	197	136
rect	196	145	197	146
rect	196	148	197	149
rect	196	151	197	152
rect	196	154	197	155
rect	196	157	197	158
rect	196	164	197	165
rect	196	167	197	168
rect	196	170	197	171
rect	196	180	197	181
rect	196	183	197	184
rect	196	187	197	188
rect	196	190	197	191
rect	197	1	198	2
rect	197	7	198	8
rect	197	10	198	11
rect	197	13	198	14
rect	197	17	198	18
rect	197	20	198	21
rect	197	23	198	24
rect	197	25	198	26
rect	197	26	198	27
rect	197	29	198	30
rect	197	32	198	33
rect	197	35	198	36
rect	197	38	198	39
rect	197	41	198	42
rect	197	44	198	45
rect	197	47	198	48
rect	197	50	198	51
rect	197	54	198	55
rect	197	56	198	57
rect	197	58	198	59
rect	197	62	198	63
rect	197	64	198	65
rect	197	69	198	70
rect	197	73	198	74
rect	197	76	198	77
rect	197	78	198	79
rect	197	81	198	82
rect	197	83	198	84
rect	197	87	198	88
rect	197	94	198	95
rect	197	100	198	101
rect	197	103	198	104
rect	197	106	198	107
rect	197	116	198	117
rect	197	119	198	120
rect	197	123	198	124
rect	197	129	198	130
rect	197	132	198	133
rect	197	135	198	136
rect	197	145	198	146
rect	197	148	198	149
rect	197	151	198	152
rect	197	154	198	155
rect	197	157	198	158
rect	197	164	198	165
rect	197	167	198	168
rect	197	170	198	171
rect	197	180	198	181
rect	197	183	198	184
rect	197	187	198	188
rect	197	190	198	191
rect	198	1	199	2
rect	198	7	199	8
rect	198	10	199	11
rect	198	13	199	14
rect	198	17	199	18
rect	198	20	199	21
rect	198	23	199	24
rect	198	25	199	26
rect	198	26	199	27
rect	198	29	199	30
rect	198	32	199	33
rect	198	35	199	36
rect	198	38	199	39
rect	198	41	199	42
rect	198	44	199	45
rect	198	47	199	48
rect	198	50	199	51
rect	198	54	199	55
rect	198	56	199	57
rect	198	58	199	59
rect	198	62	199	63
rect	198	64	199	65
rect	198	69	199	70
rect	198	73	199	74
rect	198	76	199	77
rect	198	81	199	82
rect	198	83	199	84
rect	198	87	199	88
rect	198	103	199	104
rect	198	106	199	107
rect	198	116	199	117
rect	198	119	199	120
rect	198	123	199	124
rect	198	129	199	130
rect	198	132	199	133
rect	198	135	199	136
rect	198	145	199	146
rect	198	148	199	149
rect	198	151	199	152
rect	198	154	199	155
rect	198	157	199	158
rect	198	164	199	165
rect	198	167	199	168
rect	198	170	199	171
rect	198	180	199	181
rect	198	183	199	184
rect	198	187	199	188
rect	198	190	199	191
rect	199	1	200	2
rect	199	7	200	8
rect	199	10	200	11
rect	199	13	200	14
rect	199	17	200	18
rect	199	20	200	21
rect	199	23	200	24
rect	199	25	200	26
rect	199	26	200	27
rect	199	29	200	30
rect	199	32	200	33
rect	199	35	200	36
rect	199	38	200	39
rect	199	41	200	42
rect	199	44	200	45
rect	199	47	200	48
rect	199	50	200	51
rect	199	54	200	55
rect	199	56	200	57
rect	199	58	200	59
rect	199	62	200	63
rect	199	64	200	65
rect	199	67	200	68
rect	199	69	200	70
rect	199	73	200	74
rect	199	76	200	77
rect	199	81	200	82
rect	199	83	200	84
rect	199	87	200	88
rect	199	103	200	104
rect	199	106	200	107
rect	199	116	200	117
rect	199	119	200	120
rect	199	123	200	124
rect	199	129	200	130
rect	199	132	200	133
rect	199	135	200	136
rect	199	145	200	146
rect	199	148	200	149
rect	199	151	200	152
rect	199	154	200	155
rect	199	157	200	158
rect	199	164	200	165
rect	199	167	200	168
rect	199	170	200	171
rect	199	180	200	181
rect	199	183	200	184
rect	199	187	200	188
rect	199	190	200	191
rect	200	1	201	2
rect	200	7	201	8
rect	200	10	201	11
rect	200	13	201	14
rect	200	17	201	18
rect	200	20	201	21
rect	200	23	201	24
rect	200	25	201	26
rect	200	26	201	27
rect	200	29	201	30
rect	200	32	201	33
rect	200	35	201	36
rect	200	38	201	39
rect	200	41	201	42
rect	200	44	201	45
rect	200	47	201	48
rect	200	50	201	51
rect	200	54	201	55
rect	200	56	201	57
rect	200	58	201	59
rect	200	64	201	65
rect	200	67	201	68
rect	200	69	201	70
rect	200	73	201	74
rect	200	76	201	77
rect	200	81	201	82
rect	200	83	201	84
rect	200	87	201	88
rect	200	103	201	104
rect	200	116	201	117
rect	200	119	201	120
rect	200	123	201	124
rect	200	129	201	130
rect	200	132	201	133
rect	200	135	201	136
rect	200	145	201	146
rect	200	148	201	149
rect	200	151	201	152
rect	200	154	201	155
rect	200	157	201	158
rect	200	164	201	165
rect	200	167	201	168
rect	200	170	201	171
rect	200	180	201	181
rect	200	183	201	184
rect	200	187	201	188
rect	200	190	201	191
rect	201	1	202	2
rect	201	7	202	8
rect	201	10	202	11
rect	201	13	202	14
rect	201	17	202	18
rect	201	20	202	21
rect	201	23	202	24
rect	201	25	202	26
rect	201	26	202	27
rect	201	29	202	30
rect	201	32	202	33
rect	201	35	202	36
rect	201	38	202	39
rect	201	41	202	42
rect	201	44	202	45
rect	201	47	202	48
rect	201	50	202	51
rect	201	54	202	55
rect	201	56	202	57
rect	201	58	202	59
rect	201	64	202	65
rect	201	67	202	68
rect	201	69	202	70
rect	201	73	202	74
rect	201	76	202	77
rect	201	79	202	80
rect	201	81	202	82
rect	201	83	202	84
rect	201	87	202	88
rect	201	92	202	93
rect	201	103	202	104
rect	201	116	202	117
rect	201	119	202	120
rect	201	123	202	124
rect	201	129	202	130
rect	201	132	202	133
rect	201	135	202	136
rect	201	145	202	146
rect	201	148	202	149
rect	201	151	202	152
rect	201	154	202	155
rect	201	157	202	158
rect	201	164	202	165
rect	201	167	202	168
rect	201	170	202	171
rect	201	180	202	181
rect	201	183	202	184
rect	201	187	202	188
rect	201	190	202	191
rect	202	1	203	2
rect	202	7	203	8
rect	202	10	203	11
rect	202	13	203	14
rect	202	17	203	18
rect	202	20	203	21
rect	202	23	203	24
rect	202	25	203	26
rect	202	26	203	27
rect	202	29	203	30
rect	202	32	203	33
rect	202	35	203	36
rect	202	38	203	39
rect	202	41	203	42
rect	202	44	203	45
rect	202	47	203	48
rect	202	50	203	51
rect	202	54	203	55
rect	202	56	203	57
rect	202	58	203	59
rect	202	64	203	65
rect	202	67	203	68
rect	202	69	203	70
rect	202	73	203	74
rect	202	76	203	77
rect	202	79	203	80
rect	202	81	203	82
rect	202	83	203	84
rect	202	87	203	88
rect	202	92	203	93
rect	202	103	203	104
rect	202	119	203	120
rect	202	123	203	124
rect	202	129	203	130
rect	202	135	203	136
rect	202	145	203	146
rect	202	148	203	149
rect	202	151	203	152
rect	202	154	203	155
rect	202	157	203	158
rect	202	164	203	165
rect	202	167	203	168
rect	202	170	203	171
rect	202	180	203	181
rect	202	183	203	184
rect	202	187	203	188
rect	202	190	203	191
rect	203	1	204	2
rect	203	7	204	8
rect	203	10	204	11
rect	203	13	204	14
rect	203	17	204	18
rect	203	20	204	21
rect	203	23	204	24
rect	203	25	204	26
rect	203	26	204	27
rect	203	29	204	30
rect	203	32	204	33
rect	203	35	204	36
rect	203	38	204	39
rect	203	41	204	42
rect	203	44	204	45
rect	203	47	204	48
rect	203	50	204	51
rect	203	54	204	55
rect	203	56	204	57
rect	203	58	204	59
rect	203	61	204	62
rect	203	64	204	65
rect	203	67	204	68
rect	203	69	204	70
rect	203	73	204	74
rect	203	76	204	77
rect	203	79	204	80
rect	203	81	204	82
rect	203	83	204	84
rect	203	87	204	88
rect	203	92	204	93
rect	203	103	204	104
rect	203	119	204	120
rect	203	121	204	122
rect	203	123	204	124
rect	203	129	204	130
rect	203	135	204	136
rect	203	145	204	146
rect	203	148	204	149
rect	203	151	204	152
rect	203	154	204	155
rect	203	157	204	158
rect	203	164	204	165
rect	203	167	204	168
rect	203	170	204	171
rect	203	180	204	181
rect	203	183	204	184
rect	203	187	204	188
rect	203	190	204	191
rect	204	1	205	2
rect	204	7	205	8
rect	204	10	205	11
rect	204	13	205	14
rect	204	17	205	18
rect	204	20	205	21
rect	204	23	205	24
rect	204	25	205	26
rect	204	26	205	27
rect	204	32	205	33
rect	204	35	205	36
rect	204	41	205	42
rect	204	47	205	48
rect	204	50	205	51
rect	204	54	205	55
rect	204	56	205	57
rect	204	58	205	59
rect	204	61	205	62
rect	204	64	205	65
rect	204	67	205	68
rect	204	69	205	70
rect	204	73	205	74
rect	204	76	205	77
rect	204	79	205	80
rect	204	81	205	82
rect	204	83	205	84
rect	204	87	205	88
rect	204	92	205	93
rect	204	103	205	104
rect	204	119	205	120
rect	204	121	205	122
rect	204	123	205	124
rect	204	129	205	130
rect	204	135	205	136
rect	204	148	205	149
rect	204	151	205	152
rect	204	154	205	155
rect	204	157	205	158
rect	204	167	205	168
rect	204	170	205	171
rect	204	180	205	181
rect	204	183	205	184
rect	204	187	205	188
rect	204	190	205	191
rect	205	1	206	2
rect	205	7	206	8
rect	205	10	206	11
rect	205	13	206	14
rect	205	17	206	18
rect	205	20	206	21
rect	205	23	206	24
rect	205	25	206	26
rect	205	26	206	27
rect	205	32	206	33
rect	205	35	206	36
rect	205	41	206	42
rect	205	47	206	48
rect	205	50	206	51
rect	205	54	206	55
rect	205	56	206	57
rect	205	58	206	59
rect	205	61	206	62
rect	205	64	206	65
rect	205	67	206	68
rect	205	69	206	70
rect	205	73	206	74
rect	205	76	206	77
rect	205	79	206	80
rect	205	81	206	82
rect	205	83	206	84
rect	205	87	206	88
rect	205	92	206	93
rect	205	103	206	104
rect	205	119	206	120
rect	205	121	206	122
rect	205	123	206	124
rect	205	129	206	130
rect	205	131	206	132
rect	205	135	206	136
rect	205	148	206	149
rect	205	151	206	152
rect	205	154	206	155
rect	205	157	206	158
rect	205	167	206	168
rect	205	170	206	171
rect	205	180	206	181
rect	205	183	206	184
rect	205	187	206	188
rect	205	190	206	191
rect	206	1	207	2
rect	206	7	207	8
rect	206	10	207	11
rect	206	13	207	14
rect	206	17	207	18
rect	206	20	207	21
rect	206	23	207	24
rect	206	25	207	26
rect	206	26	207	27
rect	206	32	207	33
rect	206	35	207	36
rect	206	47	207	48
rect	206	54	207	55
rect	206	56	207	57
rect	206	58	207	59
rect	206	61	207	62
rect	206	64	207	65
rect	206	67	207	68
rect	206	73	207	74
rect	206	76	207	77
rect	206	79	207	80
rect	206	81	207	82
rect	206	83	207	84
rect	206	87	207	88
rect	206	92	207	93
rect	206	103	207	104
rect	206	119	207	120
rect	206	121	207	122
rect	206	123	207	124
rect	206	129	207	130
rect	206	131	207	132
rect	206	135	207	136
rect	206	148	207	149
rect	206	151	207	152
rect	206	154	207	155
rect	206	167	207	168
rect	206	170	207	171
rect	206	180	207	181
rect	206	183	207	184
rect	206	187	207	188
rect	206	190	207	191
rect	207	1	208	2
rect	207	7	208	8
rect	207	10	208	11
rect	207	13	208	14
rect	207	17	208	18
rect	207	20	208	21
rect	207	23	208	24
rect	207	25	208	26
rect	207	26	208	27
rect	207	32	208	33
rect	207	35	208	36
rect	207	39	208	40
rect	207	45	208	46
rect	207	47	208	48
rect	207	54	208	55
rect	207	56	208	57
rect	207	58	208	59
rect	207	61	208	62
rect	207	64	208	65
rect	207	67	208	68
rect	207	73	208	74
rect	207	76	208	77
rect	207	79	208	80
rect	207	81	208	82
rect	207	83	208	84
rect	207	87	208	88
rect	207	92	208	93
rect	207	99	208	100
rect	207	103	208	104
rect	207	105	208	106
rect	207	115	208	116
rect	207	119	208	120
rect	207	121	208	122
rect	207	123	208	124
rect	207	129	208	130
rect	207	131	208	132
rect	207	135	208	136
rect	207	146	208	147
rect	207	148	208	149
rect	207	151	208	152
rect	207	154	208	155
rect	207	167	208	168
rect	207	170	208	171
rect	207	180	208	181
rect	207	183	208	184
rect	207	187	208	188
rect	207	190	208	191
rect	208	1	209	2
rect	208	7	209	8
rect	208	10	209	11
rect	208	13	209	14
rect	208	17	209	18
rect	208	20	209	21
rect	208	23	209	24
rect	208	25	209	26
rect	208	26	209	27
rect	208	39	209	40
rect	208	45	209	46
rect	208	47	209	48
rect	208	54	209	55
rect	208	56	209	57
rect	208	58	209	59
rect	208	61	209	62
rect	208	64	209	65
rect	208	67	209	68
rect	208	73	209	74
rect	208	76	209	77
rect	208	79	209	80
rect	208	81	209	82
rect	208	83	209	84
rect	208	87	209	88
rect	208	92	209	93
rect	208	99	209	100
rect	208	103	209	104
rect	208	105	209	106
rect	208	115	209	116
rect	208	119	209	120
rect	208	121	209	122
rect	208	129	209	130
rect	208	131	209	132
rect	208	146	209	147
rect	208	148	209	149
rect	208	151	209	152
rect	208	167	209	168
rect	208	170	209	171
rect	208	180	209	181
rect	208	183	209	184
rect	208	187	209	188
rect	208	190	209	191
rect	209	1	210	2
rect	209	7	210	8
rect	209	10	210	11
rect	209	13	210	14
rect	209	17	210	18
rect	209	20	210	21
rect	209	23	210	24
rect	209	25	210	26
rect	209	26	210	27
rect	209	39	210	40
rect	209	42	210	43
rect	209	45	210	46
rect	209	47	210	48
rect	209	54	210	55
rect	209	56	210	57
rect	209	58	210	59
rect	209	61	210	62
rect	209	64	210	65
rect	209	67	210	68
rect	209	73	210	74
rect	209	76	210	77
rect	209	79	210	80
rect	209	81	210	82
rect	209	83	210	84
rect	209	87	210	88
rect	209	92	210	93
rect	209	99	210	100
rect	209	103	210	104
rect	209	105	210	106
rect	209	115	210	116
rect	209	119	210	120
rect	209	121	210	122
rect	209	127	210	128
rect	209	129	210	130
rect	209	131	210	132
rect	209	143	210	144
rect	209	146	210	147
rect	209	148	210	149
rect	209	151	210	152
rect	209	167	210	168
rect	209	170	210	171
rect	209	180	210	181
rect	209	183	210	184
rect	209	187	210	188
rect	209	190	210	191
rect	210	1	211	2
rect	210	7	211	8
rect	210	10	211	11
rect	210	13	211	14
rect	210	17	211	18
rect	210	20	211	21
rect	210	23	211	24
rect	210	25	211	26
rect	210	26	211	27
rect	210	39	211	40
rect	210	42	211	43
rect	210	45	211	46
rect	210	54	211	55
rect	210	58	211	59
rect	210	61	211	62
rect	210	64	211	65
rect	210	67	211	68
rect	210	73	211	74
rect	210	76	211	77
rect	210	79	211	80
rect	210	83	211	84
rect	210	87	211	88
rect	210	92	211	93
rect	210	99	211	100
rect	210	105	211	106
rect	210	115	211	116
rect	210	121	211	122
rect	210	127	211	128
rect	210	129	211	130
rect	210	131	211	132
rect	210	143	211	144
rect	210	146	211	147
rect	210	151	211	152
rect	210	167	211	168
rect	210	170	211	171
rect	210	180	211	181
rect	210	183	211	184
rect	210	187	211	188
rect	210	190	211	191
rect	211	1	212	2
rect	211	7	212	8
rect	211	10	212	11
rect	211	13	212	14
rect	211	17	212	18
rect	211	20	212	21
rect	211	23	212	24
rect	211	25	212	26
rect	211	26	212	27
rect	211	29	212	30
rect	211	39	212	40
rect	211	42	212	43
rect	211	45	212	46
rect	211	51	212	52
rect	211	54	212	55
rect	211	58	212	59
rect	211	61	212	62
rect	211	64	212	65
rect	211	67	212	68
rect	211	70	212	71
rect	211	73	212	74
rect	211	76	212	77
rect	211	79	212	80
rect	211	83	212	84
rect	211	87	212	88
rect	211	89	212	90
rect	211	92	212	93
rect	211	99	212	100
rect	211	105	212	106
rect	211	108	212	109
rect	211	115	212	116
rect	211	121	212	122
rect	211	124	212	125
rect	211	127	212	128
rect	211	129	212	130
rect	211	131	212	132
rect	211	143	212	144
rect	211	146	212	147
rect	211	151	212	152
rect	211	153	212	154
rect	211	159	212	160
rect	211	167	212	168
rect	211	170	212	171
rect	211	180	212	181
rect	211	183	212	184
rect	211	187	212	188
rect	211	190	212	191
rect	212	1	213	2
rect	212	10	213	11
rect	212	13	213	14
rect	212	17	213	18
rect	212	20	213	21
rect	212	23	213	24
rect	212	26	213	27
rect	212	29	213	30
rect	212	39	213	40
rect	212	42	213	43
rect	212	45	213	46
rect	212	51	213	52
rect	212	54	213	55
rect	212	58	213	59
rect	212	61	213	62
rect	212	64	213	65
rect	212	67	213	68
rect	212	70	213	71
rect	212	73	213	74
rect	212	76	213	77
rect	212	79	213	80
rect	212	83	213	84
rect	212	89	213	90
rect	212	92	213	93
rect	212	99	213	100
rect	212	105	213	106
rect	212	108	213	109
rect	212	115	213	116
rect	212	121	213	122
rect	212	124	213	125
rect	212	127	213	128
rect	212	129	213	130
rect	212	131	213	132
rect	212	143	213	144
rect	212	146	213	147
rect	212	153	213	154
rect	212	159	213	160
rect	212	167	213	168
rect	212	180	213	181
rect	212	183	213	184
rect	212	187	213	188
rect	212	190	213	191
rect	213	1	214	2
rect	213	4	214	5
rect	213	10	214	11
rect	213	13	214	14
rect	213	17	214	18
rect	213	20	214	21
rect	213	23	214	24
rect	213	26	214	27
rect	213	29	214	30
rect	213	33	214	34
rect	213	39	214	40
rect	213	42	214	43
rect	213	45	214	46
rect	213	48	214	49
rect	213	51	214	52
rect	213	54	214	55
rect	213	58	214	59
rect	213	61	214	62
rect	213	64	214	65
rect	213	67	214	68
rect	213	70	214	71
rect	213	73	214	74
rect	213	76	214	77
rect	213	79	214	80
rect	213	83	214	84
rect	213	89	214	90
rect	213	92	214	93
rect	213	95	214	96
rect	213	99	214	100
rect	213	105	214	106
rect	213	108	214	109
rect	213	115	214	116
rect	213	121	214	122
rect	213	124	214	125
rect	213	127	214	128
rect	213	129	214	130
rect	213	131	214	132
rect	213	134	214	135
rect	213	140	214	141
rect	213	143	214	144
rect	213	146	214	147
rect	213	153	214	154
rect	213	159	214	160
rect	213	162	214	163
rect	213	167	214	168
rect	213	180	214	181
rect	213	183	214	184
rect	213	187	214	188
rect	213	190	214	191
rect	214	1	215	2
rect	214	4	215	5
rect	214	10	215	11
rect	214	13	215	14
rect	214	17	215	18
rect	214	20	215	21
rect	214	23	215	24
rect	214	26	215	27
rect	214	29	215	30
rect	214	33	215	34
rect	214	39	215	40
rect	214	42	215	43
rect	214	45	215	46
rect	214	48	215	49
rect	214	51	215	52
rect	214	54	215	55
rect	214	58	215	59
rect	214	61	215	62
rect	214	64	215	65
rect	214	67	215	68
rect	214	70	215	71
rect	214	73	215	74
rect	214	76	215	77
rect	214	79	215	80
rect	214	83	215	84
rect	214	89	215	90
rect	214	92	215	93
rect	214	95	215	96
rect	214	99	215	100
rect	214	105	215	106
rect	214	108	215	109
rect	214	115	215	116
rect	214	121	215	122
rect	214	124	215	125
rect	214	127	215	128
rect	214	129	215	130
rect	214	131	215	132
rect	214	134	215	135
rect	214	140	215	141
rect	214	143	215	144
rect	214	146	215	147
rect	214	153	215	154
rect	214	159	215	160
rect	214	162	215	163
rect	214	167	215	168
rect	214	180	215	181
rect	214	183	215	184
rect	214	187	215	188
rect	214	190	215	191
rect	215	1	216	2
rect	215	4	216	5
rect	215	8	216	9
rect	215	10	216	11
rect	215	13	216	14
rect	215	17	216	18
rect	215	20	216	21
rect	215	23	216	24
rect	215	26	216	27
rect	215	29	216	30
rect	215	33	216	34
rect	215	39	216	40
rect	215	42	216	43
rect	215	45	216	46
rect	215	48	216	49
rect	215	51	216	52
rect	215	54	216	55
rect	215	58	216	59
rect	215	61	216	62
rect	215	64	216	65
rect	215	67	216	68
rect	215	70	216	71
rect	215	73	216	74
rect	215	76	216	77
rect	215	79	216	80
rect	215	83	216	84
rect	215	89	216	90
rect	215	92	216	93
rect	215	95	216	96
rect	215	99	216	100
rect	215	105	216	106
rect	215	108	216	109
rect	215	115	216	116
rect	215	121	216	122
rect	215	124	216	125
rect	215	127	216	128
rect	215	129	216	130
rect	215	131	216	132
rect	215	134	216	135
rect	215	140	216	141
rect	215	143	216	144
rect	215	146	216	147
rect	215	153	216	154
rect	215	159	216	160
rect	215	162	216	163
rect	215	167	216	168
rect	215	169	216	170
rect	215	180	216	181
rect	215	183	216	184
rect	215	187	216	188
rect	215	190	216	191
rect	216	4	217	5
rect	216	8	217	9
rect	216	10	217	11
rect	216	13	217	14
rect	216	17	217	18
rect	216	20	217	21
rect	216	23	217	24
rect	216	26	217	27
rect	216	29	217	30
rect	216	33	217	34
rect	216	39	217	40
rect	216	42	217	43
rect	216	45	217	46
rect	216	48	217	49
rect	216	51	217	52
rect	216	54	217	55
rect	216	58	217	59
rect	216	61	217	62
rect	216	64	217	65
rect	216	67	217	68
rect	216	70	217	71
rect	216	73	217	74
rect	216	76	217	77
rect	216	79	217	80
rect	216	83	217	84
rect	216	89	217	90
rect	216	92	217	93
rect	216	95	217	96
rect	216	99	217	100
rect	216	105	217	106
rect	216	108	217	109
rect	216	115	217	116
rect	216	121	217	122
rect	216	124	217	125
rect	216	127	217	128
rect	216	129	217	130
rect	216	131	217	132
rect	216	134	217	135
rect	216	140	217	141
rect	216	143	217	144
rect	216	146	217	147
rect	216	153	217	154
rect	216	159	217	160
rect	216	162	217	163
rect	216	167	217	168
rect	216	169	217	170
rect	216	180	217	181
rect	216	187	217	188
rect	217	4	218	5
rect	217	8	218	9
rect	217	10	218	11
rect	217	13	218	14
rect	217	17	218	18
rect	217	20	218	21
rect	217	23	218	24
rect	217	26	218	27
rect	217	29	218	30
rect	217	33	218	34
rect	217	39	218	40
rect	217	42	218	43
rect	217	45	218	46
rect	217	48	218	49
rect	217	51	218	52
rect	217	54	218	55
rect	217	58	218	59
rect	217	61	218	62
rect	217	64	218	65
rect	217	67	218	68
rect	217	70	218	71
rect	217	73	218	74
rect	217	76	218	77
rect	217	79	218	80
rect	217	83	218	84
rect	217	89	218	90
rect	217	92	218	93
rect	217	95	218	96
rect	217	99	218	100
rect	217	105	218	106
rect	217	108	218	109
rect	217	115	218	116
rect	217	121	218	122
rect	217	124	218	125
rect	217	127	218	128
rect	217	129	218	130
rect	217	131	218	132
rect	217	134	218	135
rect	217	140	218	141
rect	217	143	218	144
rect	217	146	218	147
rect	217	153	218	154
rect	217	156	218	157
rect	217	159	218	160
rect	217	162	218	163
rect	217	167	218	168
rect	217	169	218	170
rect	217	180	218	181
rect	217	187	218	188
rect	218	4	219	5
rect	218	8	219	9
rect	218	17	219	18
rect	218	20	219	21
rect	218	23	219	24
rect	218	29	219	30
rect	218	33	219	34
rect	218	39	219	40
rect	218	42	219	43
rect	218	45	219	46
rect	218	48	219	49
rect	218	51	219	52
rect	218	54	219	55
rect	218	58	219	59
rect	218	61	219	62
rect	218	64	219	65
rect	218	67	219	68
rect	218	70	219	71
rect	218	73	219	74
rect	218	76	219	77
rect	218	79	219	80
rect	218	83	219	84
rect	218	89	219	90
rect	218	92	219	93
rect	218	95	219	96
rect	218	99	219	100
rect	218	105	219	106
rect	218	108	219	109
rect	218	115	219	116
rect	218	121	219	122
rect	218	124	219	125
rect	218	127	219	128
rect	218	131	219	132
rect	218	134	219	135
rect	218	140	219	141
rect	218	143	219	144
rect	218	146	219	147
rect	218	153	219	154
rect	218	156	219	157
rect	218	159	219	160
rect	218	162	219	163
rect	218	169	219	170
rect	219	1	220	2
rect	219	4	220	5
rect	219	8	220	9
rect	219	14	220	15
rect	219	17	220	18
rect	219	20	220	21
rect	219	23	220	24
rect	219	26	220	27
rect	219	29	220	30
rect	219	33	220	34
rect	219	39	220	40
rect	219	42	220	43
rect	219	45	220	46
rect	219	48	220	49
rect	219	51	220	52
rect	219	54	220	55
rect	219	58	220	59
rect	219	61	220	62
rect	219	64	220	65
rect	219	67	220	68
rect	219	70	220	71
rect	219	73	220	74
rect	219	76	220	77
rect	219	79	220	80
rect	219	83	220	84
rect	219	89	220	90
rect	219	92	220	93
rect	219	95	220	96
rect	219	99	220	100
rect	219	105	220	106
rect	219	108	220	109
rect	219	112	220	113
rect	219	115	220	116
rect	219	118	220	119
rect	219	121	220	122
rect	219	124	220	125
rect	219	127	220	128
rect	219	131	220	132
rect	219	134	220	135
rect	219	137	220	138
rect	219	140	220	141
rect	219	143	220	144
rect	219	146	220	147
rect	219	153	220	154
rect	219	156	220	157
rect	219	159	220	160
rect	219	162	220	163
rect	219	169	220	170
rect	220	23	221	24
rect	220	26	221	27
rect	221	23	222	24
rect	221	26	222	27
rect	222	23	223	24
rect	222	26	223	27
rect	223	23	224	24
rect	223	26	224	27
rect	224	23	225	24
rect	224	26	225	27
rect	225	23	226	24
rect	225	26	226	27
rect	226	4	227	5
rect	226	14	227	15
rect	226	17	227	18
rect	226	20	227	21
rect	226	23	227	24
rect	226	26	227	27
rect	226	29	227	30
rect	226	33	227	34
rect	226	39	227	40
rect	226	42	227	43
rect	226	45	227	46
rect	226	48	227	49
rect	226	51	227	52
rect	226	54	227	55
rect	226	58	227	59
rect	226	61	227	62
rect	226	64	227	65
rect	226	67	227	68
rect	226	70	227	71
rect	226	73	227	74
rect	226	76	227	77
rect	226	79	227	80
rect	226	86	227	87
rect	226	89	227	90
rect	226	92	227	93
rect	226	95	227	96
rect	226	99	227	100
rect	226	102	227	103
rect	226	105	227	106
rect	226	108	227	109
rect	226	112	227	113
rect	226	115	227	116
rect	226	118	227	119
rect	226	121	227	122
rect	226	124	227	125
rect	226	127	227	128
rect	226	131	227	132
rect	226	134	227	135
rect	226	137	227	138
rect	226	140	227	141
rect	226	143	227	144
rect	226	146	227	147
rect	226	156	227	157
rect	226	159	227	160
rect	226	162	227	163
rect	226	166	227	167
rect	227	4	228	5
rect	227	14	228	15
rect	227	17	228	18
rect	227	20	228	21
rect	227	23	228	24
rect	227	26	228	27
rect	227	29	228	30
rect	227	33	228	34
rect	227	39	228	40
rect	227	42	228	43
rect	227	45	228	46
rect	227	48	228	49
rect	227	51	228	52
rect	227	54	228	55
rect	227	58	228	59
rect	227	61	228	62
rect	227	64	228	65
rect	227	67	228	68
rect	227	70	228	71
rect	227	73	228	74
rect	227	76	228	77
rect	227	79	228	80
rect	227	86	228	87
rect	227	89	228	90
rect	227	92	228	93
rect	227	95	228	96
rect	227	99	228	100
rect	227	102	228	103
rect	227	105	228	106
rect	227	108	228	109
rect	227	112	228	113
rect	227	115	228	116
rect	227	118	228	119
rect	227	121	228	122
rect	227	124	228	125
rect	227	127	228	128
rect	227	131	228	132
rect	227	134	228	135
rect	227	137	228	138
rect	227	140	228	141
rect	227	143	228	144
rect	227	146	228	147
rect	227	156	228	157
rect	227	159	228	160
rect	227	162	228	163
rect	227	166	228	167
rect	228	4	229	5
rect	228	14	229	15
rect	228	17	229	18
rect	228	20	229	21
rect	228	23	229	24
rect	228	26	229	27
rect	228	29	229	30
rect	228	33	229	34
rect	228	39	229	40
rect	228	42	229	43
rect	228	45	229	46
rect	228	48	229	49
rect	228	51	229	52
rect	228	54	229	55
rect	228	58	229	59
rect	228	61	229	62
rect	228	64	229	65
rect	228	67	229	68
rect	228	70	229	71
rect	228	73	229	74
rect	228	76	229	77
rect	228	79	229	80
rect	228	86	229	87
rect	228	89	229	90
rect	228	92	229	93
rect	228	95	229	96
rect	228	99	229	100
rect	228	102	229	103
rect	228	105	229	106
rect	228	108	229	109
rect	228	112	229	113
rect	228	115	229	116
rect	228	118	229	119
rect	228	121	229	122
rect	228	124	229	125
rect	228	127	229	128
rect	228	131	229	132
rect	228	134	229	135
rect	228	137	229	138
rect	228	140	229	141
rect	228	143	229	144
rect	228	146	229	147
rect	228	156	229	157
rect	228	159	229	160
rect	228	162	229	163
rect	228	166	229	167
rect	229	4	230	5
rect	229	14	230	15
rect	229	17	230	18
rect	229	20	230	21
rect	229	23	230	24
rect	229	26	230	27
rect	229	29	230	30
rect	229	33	230	34
rect	229	39	230	40
rect	229	42	230	43
rect	229	45	230	46
rect	229	48	230	49
rect	229	51	230	52
rect	229	54	230	55
rect	229	58	230	59
rect	229	61	230	62
rect	229	64	230	65
rect	229	67	230	68
rect	229	70	230	71
rect	229	73	230	74
rect	229	76	230	77
rect	229	79	230	80
rect	229	86	230	87
rect	229	89	230	90
rect	229	92	230	93
rect	229	95	230	96
rect	229	99	230	100
rect	229	102	230	103
rect	229	105	230	106
rect	229	108	230	109
rect	229	112	230	113
rect	229	115	230	116
rect	229	118	230	119
rect	229	121	230	122
rect	229	124	230	125
rect	229	127	230	128
rect	229	131	230	132
rect	229	134	230	135
rect	229	137	230	138
rect	229	140	230	141
rect	229	143	230	144
rect	229	146	230	147
rect	229	156	230	157
rect	229	159	230	160
rect	229	162	230	163
rect	229	166	230	167
rect	230	4	231	5
rect	230	14	231	15
rect	230	17	231	18
rect	230	20	231	21
rect	230	23	231	24
rect	230	26	231	27
rect	230	29	231	30
rect	230	33	231	34
rect	230	39	231	40
rect	230	42	231	43
rect	230	45	231	46
rect	230	48	231	49
rect	230	51	231	52
rect	230	54	231	55
rect	230	58	231	59
rect	230	61	231	62
rect	230	64	231	65
rect	230	67	231	68
rect	230	70	231	71
rect	230	73	231	74
rect	230	76	231	77
rect	230	79	231	80
rect	230	86	231	87
rect	230	89	231	90
rect	230	92	231	93
rect	230	95	231	96
rect	230	99	231	100
rect	230	102	231	103
rect	230	105	231	106
rect	230	108	231	109
rect	230	112	231	113
rect	230	115	231	116
rect	230	118	231	119
rect	230	121	231	122
rect	230	124	231	125
rect	230	127	231	128
rect	230	131	231	132
rect	230	134	231	135
rect	230	137	231	138
rect	230	140	231	141
rect	230	143	231	144
rect	230	146	231	147
rect	230	156	231	157
rect	230	159	231	160
rect	230	162	231	163
rect	230	166	231	167
rect	231	4	232	5
rect	231	14	232	15
rect	231	17	232	18
rect	231	20	232	21
rect	231	23	232	24
rect	231	26	232	27
rect	231	29	232	30
rect	231	33	232	34
rect	231	39	232	40
rect	231	42	232	43
rect	231	45	232	46
rect	231	48	232	49
rect	231	51	232	52
rect	231	54	232	55
rect	231	58	232	59
rect	231	61	232	62
rect	231	64	232	65
rect	231	67	232	68
rect	231	70	232	71
rect	231	73	232	74
rect	231	76	232	77
rect	231	79	232	80
rect	231	86	232	87
rect	231	89	232	90
rect	231	92	232	93
rect	231	95	232	96
rect	231	99	232	100
rect	231	102	232	103
rect	231	105	232	106
rect	231	108	232	109
rect	231	112	232	113
rect	231	115	232	116
rect	231	118	232	119
rect	231	121	232	122
rect	231	124	232	125
rect	231	127	232	128
rect	231	131	232	132
rect	231	134	232	135
rect	231	137	232	138
rect	231	140	232	141
rect	231	143	232	144
rect	231	146	232	147
rect	231	156	232	157
rect	231	159	232	160
rect	231	162	232	163
rect	231	166	232	167
rect	232	4	233	5
rect	232	14	233	15
rect	232	17	233	18
rect	232	20	233	21
rect	232	23	233	24
rect	232	26	233	27
rect	232	29	233	30
rect	232	33	233	34
rect	232	39	233	40
rect	232	42	233	43
rect	232	45	233	46
rect	232	48	233	49
rect	232	51	233	52
rect	232	54	233	55
rect	232	58	233	59
rect	232	61	233	62
rect	232	64	233	65
rect	232	67	233	68
rect	232	70	233	71
rect	232	73	233	74
rect	232	76	233	77
rect	232	79	233	80
rect	232	86	233	87
rect	232	89	233	90
rect	232	92	233	93
rect	232	95	233	96
rect	232	99	233	100
rect	232	102	233	103
rect	232	105	233	106
rect	232	108	233	109
rect	232	112	233	113
rect	232	115	233	116
rect	232	118	233	119
rect	232	121	233	122
rect	232	124	233	125
rect	232	127	233	128
rect	232	131	233	132
rect	232	134	233	135
rect	232	137	233	138
rect	232	140	233	141
rect	232	143	233	144
rect	232	146	233	147
rect	232	156	233	157
rect	232	159	233	160
rect	232	162	233	163
rect	232	166	233	167
rect	233	4	234	5
rect	233	14	234	15
rect	233	17	234	18
rect	233	20	234	21
rect	233	23	234	24
rect	233	26	234	27
rect	233	29	234	30
rect	233	39	234	40
rect	233	42	234	43
rect	233	45	234	46
rect	233	48	234	49
rect	233	51	234	52
rect	233	54	234	55
rect	233	58	234	59
rect	233	61	234	62
rect	233	64	234	65
rect	233	67	234	68
rect	233	70	234	71
rect	233	73	234	74
rect	233	76	234	77
rect	233	79	234	80
rect	233	86	234	87
rect	233	89	234	90
rect	233	92	234	93
rect	233	95	234	96
rect	233	99	234	100
rect	233	102	234	103
rect	233	108	234	109
rect	233	112	234	113
rect	233	115	234	116
rect	233	118	234	119
rect	233	121	234	122
rect	233	124	234	125
rect	233	127	234	128
rect	233	131	234	132
rect	233	134	234	135
rect	233	137	234	138
rect	233	140	234	141
rect	233	143	234	144
rect	233	146	234	147
rect	233	156	234	157
rect	233	159	234	160
rect	233	162	234	163
rect	233	166	234	167
rect	234	4	235	5
rect	234	14	235	15
rect	234	17	235	18
rect	234	20	235	21
rect	234	23	235	24
rect	234	26	235	27
rect	234	29	235	30
rect	234	39	235	40
rect	234	42	235	43
rect	234	45	235	46
rect	234	48	235	49
rect	234	51	235	52
rect	234	54	235	55
rect	234	58	235	59
rect	234	61	235	62
rect	234	64	235	65
rect	234	67	235	68
rect	234	70	235	71
rect	234	73	235	74
rect	234	76	235	77
rect	234	79	235	80
rect	234	86	235	87
rect	234	89	235	90
rect	234	92	235	93
rect	234	95	235	96
rect	234	99	235	100
rect	234	102	235	103
rect	234	108	235	109
rect	234	112	235	113
rect	234	115	235	116
rect	234	118	235	119
rect	234	121	235	122
rect	234	124	235	125
rect	234	127	235	128
rect	234	131	235	132
rect	234	134	235	135
rect	234	137	235	138
rect	234	140	235	141
rect	234	143	235	144
rect	234	146	235	147
rect	234	156	235	157
rect	234	159	235	160
rect	234	162	235	163
rect	234	166	235	167
rect	235	4	236	5
rect	235	14	236	15
rect	235	17	236	18
rect	235	20	236	21
rect	235	23	236	24
rect	235	26	236	27
rect	235	29	236	30
rect	235	39	236	40
rect	235	45	236	46
rect	235	48	236	49
rect	235	51	236	52
rect	235	54	236	55
rect	235	58	236	59
rect	235	61	236	62
rect	235	64	236	65
rect	235	67	236	68
rect	235	70	236	71
rect	235	73	236	74
rect	235	76	236	77
rect	235	79	236	80
rect	235	86	236	87
rect	235	89	236	90
rect	235	92	236	93
rect	235	95	236	96
rect	235	99	236	100
rect	235	102	236	103
rect	235	108	236	109
rect	235	112	236	113
rect	235	115	236	116
rect	235	118	236	119
rect	235	121	236	122
rect	235	124	236	125
rect	235	127	236	128
rect	235	131	236	132
rect	235	134	236	135
rect	235	137	236	138
rect	235	140	236	141
rect	235	143	236	144
rect	235	146	236	147
rect	235	156	236	157
rect	235	159	236	160
rect	235	162	236	163
rect	235	166	236	167
rect	236	4	237	5
rect	236	14	237	15
rect	236	17	237	18
rect	236	20	237	21
rect	236	23	237	24
rect	236	26	237	27
rect	236	29	237	30
rect	236	33	237	34
rect	236	39	237	40
rect	236	45	237	46
rect	236	48	237	49
rect	236	51	237	52
rect	236	54	237	55
rect	236	58	237	59
rect	236	61	237	62
rect	236	64	237	65
rect	236	67	237	68
rect	236	70	237	71
rect	236	73	237	74
rect	236	76	237	77
rect	236	79	237	80
rect	236	86	237	87
rect	236	89	237	90
rect	236	92	237	93
rect	236	95	237	96
rect	236	99	237	100
rect	236	102	237	103
rect	236	108	237	109
rect	236	112	237	113
rect	236	115	237	116
rect	236	118	237	119
rect	236	121	237	122
rect	236	124	237	125
rect	236	127	237	128
rect	236	131	237	132
rect	236	134	237	135
rect	236	137	237	138
rect	236	140	237	141
rect	236	143	237	144
rect	236	146	237	147
rect	236	156	237	157
rect	236	159	237	160
rect	236	162	237	163
rect	236	166	237	167
rect	237	4	238	5
rect	237	14	238	15
rect	237	17	238	18
rect	237	20	238	21
rect	237	23	238	24
rect	237	26	238	27
rect	237	29	238	30
rect	237	33	238	34
rect	237	39	238	40
rect	237	45	238	46
rect	237	48	238	49
rect	237	51	238	52
rect	237	54	238	55
rect	237	58	238	59
rect	237	61	238	62
rect	237	64	238	65
rect	237	67	238	68
rect	237	70	238	71
rect	237	76	238	77
rect	237	79	238	80
rect	237	86	238	87
rect	237	89	238	90
rect	237	92	238	93
rect	237	95	238	96
rect	237	99	238	100
rect	237	102	238	103
rect	237	108	238	109
rect	237	112	238	113
rect	237	115	238	116
rect	237	118	238	119
rect	237	121	238	122
rect	237	124	238	125
rect	237	127	238	128
rect	237	131	238	132
rect	237	134	238	135
rect	237	137	238	138
rect	237	140	238	141
rect	237	143	238	144
rect	237	146	238	147
rect	237	156	238	157
rect	237	159	238	160
rect	237	162	238	163
rect	237	166	238	167
rect	238	4	239	5
rect	238	14	239	15
rect	238	17	239	18
rect	238	20	239	21
rect	238	23	239	24
rect	238	26	239	27
rect	238	29	239	30
rect	238	33	239	34
rect	238	39	239	40
rect	238	42	239	43
rect	238	45	239	46
rect	238	48	239	49
rect	238	51	239	52
rect	238	54	239	55
rect	238	58	239	59
rect	238	61	239	62
rect	238	64	239	65
rect	238	67	239	68
rect	238	70	239	71
rect	238	76	239	77
rect	238	79	239	80
rect	238	86	239	87
rect	238	89	239	90
rect	238	92	239	93
rect	238	95	239	96
rect	238	99	239	100
rect	238	102	239	103
rect	238	108	239	109
rect	238	112	239	113
rect	238	115	239	116
rect	238	118	239	119
rect	238	121	239	122
rect	238	124	239	125
rect	238	127	239	128
rect	238	131	239	132
rect	238	134	239	135
rect	238	137	239	138
rect	238	140	239	141
rect	238	143	239	144
rect	238	146	239	147
rect	238	156	239	157
rect	238	159	239	160
rect	238	162	239	163
rect	238	166	239	167
rect	239	4	240	5
rect	239	14	240	15
rect	239	17	240	18
rect	239	20	240	21
rect	239	23	240	24
rect	239	26	240	27
rect	239	29	240	30
rect	239	33	240	34
rect	239	39	240	40
rect	239	42	240	43
rect	239	45	240	46
rect	239	48	240	49
rect	239	51	240	52
rect	239	61	240	62
rect	239	64	240	65
rect	239	67	240	68
rect	239	70	240	71
rect	239	76	240	77
rect	239	79	240	80
rect	239	89	240	90
rect	239	92	240	93
rect	239	95	240	96
rect	239	99	240	100
rect	239	102	240	103
rect	239	108	240	109
rect	239	112	240	113
rect	239	115	240	116
rect	239	118	240	119
rect	239	121	240	122
rect	239	124	240	125
rect	239	127	240	128
rect	239	131	240	132
rect	239	134	240	135
rect	239	137	240	138
rect	239	140	240	141
rect	239	143	240	144
rect	239	146	240	147
rect	239	156	240	157
rect	239	159	240	160
rect	239	162	240	163
rect	239	166	240	167
rect	240	4	241	5
rect	240	14	241	15
rect	240	17	241	18
rect	240	20	241	21
rect	240	23	241	24
rect	240	26	241	27
rect	240	29	241	30
rect	240	33	241	34
rect	240	39	241	40
rect	240	42	241	43
rect	240	45	241	46
rect	240	48	241	49
rect	240	51	241	52
rect	240	61	241	62
rect	240	64	241	65
rect	240	67	241	68
rect	240	70	241	71
rect	240	73	241	74
rect	240	76	241	77
rect	240	79	241	80
rect	240	89	241	90
rect	240	92	241	93
rect	240	95	241	96
rect	240	99	241	100
rect	240	102	241	103
rect	240	108	241	109
rect	240	112	241	113
rect	240	115	241	116
rect	240	118	241	119
rect	240	121	241	122
rect	240	124	241	125
rect	240	127	241	128
rect	240	131	241	132
rect	240	134	241	135
rect	240	137	241	138
rect	240	140	241	141
rect	240	143	241	144
rect	240	146	241	147
rect	240	156	241	157
rect	240	159	241	160
rect	240	162	241	163
rect	240	166	241	167
rect	241	4	242	5
rect	241	14	242	15
rect	241	17	242	18
rect	241	23	242	24
rect	241	26	242	27
rect	241	29	242	30
rect	241	33	242	34
rect	241	39	242	40
rect	241	42	242	43
rect	241	45	242	46
rect	241	48	242	49
rect	241	51	242	52
rect	241	67	242	68
rect	241	70	242	71
rect	241	73	242	74
rect	241	76	242	77
rect	241	79	242	80
rect	241	89	242	90
rect	241	92	242	93
rect	241	95	242	96
rect	241	99	242	100
rect	241	102	242	103
rect	241	108	242	109
rect	241	112	242	113
rect	241	115	242	116
rect	241	118	242	119
rect	241	121	242	122
rect	241	124	242	125
rect	241	127	242	128
rect	241	131	242	132
rect	241	134	242	135
rect	241	137	242	138
rect	241	140	242	141
rect	241	143	242	144
rect	241	146	242	147
rect	241	156	242	157
rect	241	159	242	160
rect	241	162	242	163
rect	241	166	242	167
rect	242	4	243	5
rect	242	14	243	15
rect	242	17	243	18
rect	242	23	243	24
rect	242	26	243	27
rect	242	29	243	30
rect	242	33	243	34
rect	242	39	243	40
rect	242	42	243	43
rect	242	45	243	46
rect	242	48	243	49
rect	242	51	243	52
rect	242	67	243	68
rect	242	70	243	71
rect	242	73	243	74
rect	242	76	243	77
rect	242	79	243	80
rect	242	83	243	84
rect	242	89	243	90
rect	242	92	243	93
rect	242	95	243	96
rect	242	99	243	100
rect	242	102	243	103
rect	242	108	243	109
rect	242	112	243	113
rect	242	115	243	116
rect	242	118	243	119
rect	242	121	243	122
rect	242	124	243	125
rect	242	127	243	128
rect	242	131	243	132
rect	242	134	243	135
rect	242	137	243	138
rect	242	140	243	141
rect	242	143	243	144
rect	242	146	243	147
rect	242	156	243	157
rect	242	159	243	160
rect	242	162	243	163
rect	242	166	243	167
rect	243	4	244	5
rect	243	14	244	15
rect	243	17	244	18
rect	243	23	244	24
rect	243	26	244	27
rect	243	29	244	30
rect	243	33	244	34
rect	243	39	244	40
rect	243	42	244	43
rect	243	45	244	46
rect	243	48	244	49
rect	243	67	244	68
rect	243	70	244	71
rect	243	73	244	74
rect	243	76	244	77
rect	243	79	244	80
rect	243	83	244	84
rect	243	89	244	90
rect	243	92	244	93
rect	243	95	244	96
rect	243	99	244	100
rect	243	102	244	103
rect	243	108	244	109
rect	243	112	244	113
rect	243	115	244	116
rect	243	118	244	119
rect	243	121	244	122
rect	243	124	244	125
rect	243	127	244	128
rect	243	131	244	132
rect	243	137	244	138
rect	243	140	244	141
rect	243	143	244	144
rect	243	146	244	147
rect	243	156	244	157
rect	243	159	244	160
rect	243	162	244	163
rect	243	166	244	167
rect	244	4	245	5
rect	244	14	245	15
rect	244	17	245	18
rect	244	20	245	21
rect	244	23	245	24
rect	244	26	245	27
rect	244	29	245	30
rect	244	33	245	34
rect	244	39	245	40
rect	244	42	245	43
rect	244	45	245	46
rect	244	48	245	49
rect	244	54	245	55
rect	244	67	245	68
rect	244	70	245	71
rect	244	73	245	74
rect	244	76	245	77
rect	244	79	245	80
rect	244	83	245	84
rect	244	89	245	90
rect	244	92	245	93
rect	244	95	245	96
rect	244	99	245	100
rect	244	102	245	103
rect	244	108	245	109
rect	244	112	245	113
rect	244	115	245	116
rect	244	118	245	119
rect	244	121	245	122
rect	244	124	245	125
rect	244	127	245	128
rect	244	131	245	132
rect	244	137	245	138
rect	244	140	245	141
rect	244	143	245	144
rect	244	146	245	147
rect	244	156	245	157
rect	244	159	245	160
rect	244	162	245	163
rect	244	166	245	167
rect	245	4	246	5
rect	245	14	246	15
rect	245	17	246	18
rect	245	20	246	21
rect	245	23	246	24
rect	245	26	246	27
rect	245	29	246	30
rect	245	33	246	34
rect	245	39	246	40
rect	245	42	246	43
rect	245	45	246	46
rect	245	48	246	49
rect	245	54	246	55
rect	245	67	246	68
rect	245	70	246	71
rect	245	73	246	74
rect	245	79	246	80
rect	245	83	246	84
rect	245	89	246	90
rect	245	92	246	93
rect	245	95	246	96
rect	245	99	246	100
rect	245	102	246	103
rect	245	108	246	109
rect	245	112	246	113
rect	245	115	246	116
rect	245	118	246	119
rect	245	121	246	122
rect	245	124	246	125
rect	245	127	246	128
rect	245	131	246	132
rect	245	137	246	138
rect	245	140	246	141
rect	245	143	246	144
rect	245	146	246	147
rect	245	156	246	157
rect	245	159	246	160
rect	245	162	246	163
rect	245	166	246	167
rect	246	4	247	5
rect	246	14	247	15
rect	246	17	247	18
rect	246	20	247	21
rect	246	23	247	24
rect	246	26	247	27
rect	246	29	247	30
rect	246	33	247	34
rect	246	39	247	40
rect	246	42	247	43
rect	246	45	247	46
rect	246	48	247	49
rect	246	51	247	52
rect	246	54	247	55
rect	246	67	247	68
rect	246	70	247	71
rect	246	73	247	74
rect	246	79	247	80
rect	246	83	247	84
rect	246	89	247	90
rect	246	92	247	93
rect	246	95	247	96
rect	246	99	247	100
rect	246	102	247	103
rect	246	108	247	109
rect	246	112	247	113
rect	246	115	247	116
rect	246	118	247	119
rect	246	121	247	122
rect	246	124	247	125
rect	246	127	247	128
rect	246	131	247	132
rect	246	137	247	138
rect	246	140	247	141
rect	246	143	247	144
rect	246	146	247	147
rect	246	156	247	157
rect	246	159	247	160
rect	246	162	247	163
rect	246	166	247	167
rect	247	4	248	5
rect	247	14	248	15
rect	247	17	248	18
rect	247	20	248	21
rect	247	23	248	24
rect	247	26	248	27
rect	247	29	248	30
rect	247	33	248	34
rect	247	42	248	43
rect	247	45	248	46
rect	247	48	248	49
rect	247	51	248	52
rect	247	54	248	55
rect	247	67	248	68
rect	247	70	248	71
rect	247	73	248	74
rect	247	79	248	80
rect	247	83	248	84
rect	247	89	248	90
rect	247	92	248	93
rect	247	95	248	96
rect	247	99	248	100
rect	247	108	248	109
rect	247	112	248	113
rect	247	115	248	116
rect	247	118	248	119
rect	247	121	248	122
rect	247	124	248	125
rect	247	127	248	128
rect	247	131	248	132
rect	247	137	248	138
rect	247	140	248	141
rect	247	143	248	144
rect	247	146	248	147
rect	247	156	248	157
rect	247	162	248	163
rect	247	166	248	167
rect	248	4	249	5
rect	248	14	249	15
rect	248	17	249	18
rect	248	20	249	21
rect	248	23	249	24
rect	248	26	249	27
rect	248	29	249	30
rect	248	33	249	34
rect	248	42	249	43
rect	248	45	249	46
rect	248	48	249	49
rect	248	51	249	52
rect	248	54	249	55
rect	248	64	249	65
rect	248	67	249	68
rect	248	70	249	71
rect	248	73	249	74
rect	248	79	249	80
rect	248	83	249	84
rect	248	86	249	87
rect	248	89	249	90
rect	248	92	249	93
rect	248	95	249	96
rect	248	99	249	100
rect	248	108	249	109
rect	248	112	249	113
rect	248	115	249	116
rect	248	118	249	119
rect	248	121	249	122
rect	248	124	249	125
rect	248	127	249	128
rect	248	129	249	130
rect	248	131	249	132
rect	248	137	249	138
rect	248	140	249	141
rect	248	143	249	144
rect	248	146	249	147
rect	248	156	249	157
rect	248	162	249	163
rect	248	166	249	167
rect	249	4	250	5
rect	249	14	250	15
rect	249	17	250	18
rect	249	20	250	21
rect	249	23	250	24
rect	249	26	250	27
rect	249	29	250	30
rect	249	33	250	34
rect	249	42	250	43
rect	249	45	250	46
rect	249	48	250	49
rect	249	51	250	52
rect	249	54	250	55
rect	249	64	250	65
rect	249	67	250	68
rect	249	73	250	74
rect	249	79	250	80
rect	249	83	250	84
rect	249	86	250	87
rect	249	89	250	90
rect	249	92	250	93
rect	249	99	250	100
rect	249	108	250	109
rect	249	112	250	113
rect	249	115	250	116
rect	249	118	250	119
rect	249	121	250	122
rect	249	124	250	125
rect	249	129	250	130
rect	249	131	250	132
rect	249	137	250	138
rect	249	140	250	141
rect	249	143	250	144
rect	249	146	250	147
rect	249	156	250	157
rect	249	162	250	163
rect	249	166	250	167
rect	250	4	251	5
rect	250	14	251	15
rect	250	17	251	18
rect	250	20	251	21
rect	250	23	251	24
rect	250	26	251	27
rect	250	29	251	30
rect	250	33	251	34
rect	250	39	251	40
rect	250	42	251	43
rect	250	45	251	46
rect	250	48	251	49
rect	250	51	251	52
rect	250	54	251	55
rect	250	64	251	65
rect	250	67	251	68
rect	250	73	251	74
rect	250	76	251	77
rect	250	79	251	80
rect	250	83	251	84
rect	250	86	251	87
rect	250	89	251	90
rect	250	92	251	93
rect	250	99	251	100
rect	250	108	251	109
rect	250	112	251	113
rect	250	115	251	116
rect	250	118	251	119
rect	250	121	251	122
rect	250	124	251	125
rect	250	129	251	130
rect	250	131	251	132
rect	250	133	251	134
rect	250	137	251	138
rect	250	140	251	141
rect	250	143	251	144
rect	250	146	251	147
rect	250	156	251	157
rect	250	162	251	163
rect	250	166	251	167
rect	251	4	252	5
rect	251	14	252	15
rect	251	20	252	21
rect	251	23	252	24
rect	251	26	252	27
rect	251	29	252	30
rect	251	33	252	34
rect	251	39	252	40
rect	251	42	252	43
rect	251	45	252	46
rect	251	48	252	49
rect	251	51	252	52
rect	251	54	252	55
rect	251	64	252	65
rect	251	73	252	74
rect	251	76	252	77
rect	251	79	252	80
rect	251	83	252	84
rect	251	86	252	87
rect	251	89	252	90
rect	251	99	252	100
rect	251	108	252	109
rect	251	112	252	113
rect	251	115	252	116
rect	251	121	252	122
rect	251	124	252	125
rect	251	129	252	130
rect	251	131	252	132
rect	251	133	252	134
rect	251	137	252	138
rect	251	140	252	141
rect	251	146	252	147
rect	251	156	252	157
rect	251	162	252	163
rect	251	166	252	167
rect	252	4	253	5
rect	252	7	253	8
rect	252	14	253	15
rect	252	20	253	21
rect	252	23	253	24
rect	252	26	253	27
rect	252	29	253	30
rect	252	33	253	34
rect	252	36	253	37
rect	252	39	253	40
rect	252	42	253	43
rect	252	45	253	46
rect	252	48	253	49
rect	252	51	253	52
rect	252	54	253	55
rect	252	64	253	65
rect	252	70	253	71
rect	252	73	253	74
rect	252	76	253	77
rect	252	79	253	80
rect	252	83	253	84
rect	252	86	253	87
rect	252	89	253	90
rect	252	99	253	100
rect	252	106	253	107
rect	252	108	253	109
rect	252	112	253	113
rect	252	115	253	116
rect	252	121	253	122
rect	252	124	253	125
rect	252	126	253	127
rect	252	129	253	130
rect	252	131	253	132
rect	252	133	253	134
rect	252	137	253	138
rect	252	140	253	141
rect	252	146	253	147
rect	252	156	253	157
rect	252	162	253	163
rect	252	166	253	167
rect	253	4	254	5
rect	253	7	254	8
rect	253	14	254	15
rect	253	20	254	21
rect	253	23	254	24
rect	253	26	254	27
rect	253	29	254	30
rect	253	33	254	34
rect	253	36	254	37
rect	253	39	254	40
rect	253	42	254	43
rect	253	45	254	46
rect	253	48	254	49
rect	253	51	254	52
rect	253	54	254	55
rect	253	64	254	65
rect	253	70	254	71
rect	253	73	254	74
rect	253	76	254	77
rect	253	79	254	80
rect	253	83	254	84
rect	253	86	254	87
rect	253	89	254	90
rect	253	106	254	107
rect	253	108	254	109
rect	253	112	254	113
rect	253	115	254	116
rect	253	121	254	122
rect	253	124	254	125
rect	253	126	254	127
rect	253	129	254	130
rect	253	131	254	132
rect	253	133	254	134
rect	253	137	254	138
rect	253	146	254	147
rect	253	156	254	157
rect	253	162	254	163
rect	253	166	254	167
rect	254	4	255	5
rect	254	7	255	8
rect	254	14	255	15
rect	254	17	255	18
rect	254	20	255	21
rect	254	23	255	24
rect	254	26	255	27
rect	254	29	255	30
rect	254	33	255	34
rect	254	36	255	37
rect	254	39	255	40
rect	254	42	255	43
rect	254	45	255	46
rect	254	48	255	49
rect	254	51	255	52
rect	254	54	255	55
rect	254	64	255	65
rect	254	70	255	71
rect	254	73	255	74
rect	254	76	255	77
rect	254	79	255	80
rect	254	83	255	84
rect	254	86	255	87
rect	254	89	255	90
rect	254	102	255	103
rect	254	106	255	107
rect	254	108	255	109
rect	254	112	255	113
rect	254	115	255	116
rect	254	121	255	122
rect	254	124	255	125
rect	254	126	255	127
rect	254	129	255	130
rect	254	131	255	132
rect	254	133	255	134
rect	254	137	255	138
rect	254	146	255	147
rect	254	156	255	157
rect	254	162	255	163
rect	254	166	255	167
rect	255	4	256	5
rect	255	7	256	8
rect	255	14	256	15
rect	255	17	256	18
rect	255	20	256	21
rect	255	23	256	24
rect	255	26	256	27
rect	255	29	256	30
rect	255	33	256	34
rect	255	36	256	37
rect	255	39	256	40
rect	255	42	256	43
rect	255	45	256	46
rect	255	48	256	49
rect	255	51	256	52
rect	255	54	256	55
rect	255	64	256	65
rect	255	70	256	71
rect	255	73	256	74
rect	255	76	256	77
rect	255	79	256	80
rect	255	83	256	84
rect	255	86	256	87
rect	255	102	256	103
rect	255	106	256	107
rect	255	108	256	109
rect	255	112	256	113
rect	255	115	256	116
rect	255	121	256	122
rect	255	124	256	125
rect	255	126	256	127
rect	255	129	256	130
rect	255	131	256	132
rect	255	133	256	134
rect	255	146	256	147
rect	255	156	256	157
rect	255	162	256	163
rect	255	166	256	167
rect	256	4	257	5
rect	256	7	257	8
rect	256	14	257	15
rect	256	17	257	18
rect	256	20	257	21
rect	256	23	257	24
rect	256	26	257	27
rect	256	29	257	30
rect	256	33	257	34
rect	256	36	257	37
rect	256	39	257	40
rect	256	42	257	43
rect	256	45	257	46
rect	256	48	257	49
rect	256	51	257	52
rect	256	54	257	55
rect	256	64	257	65
rect	256	67	257	68
rect	256	70	257	71
rect	256	73	257	74
rect	256	76	257	77
rect	256	79	257	80
rect	256	83	257	84
rect	256	86	257	87
rect	256	99	257	100
rect	256	102	257	103
rect	256	106	257	107
rect	256	108	257	109
rect	256	112	257	113
rect	256	115	257	116
rect	256	121	257	122
rect	256	124	257	125
rect	256	126	257	127
rect	256	129	257	130
rect	256	131	257	132
rect	256	133	257	134
rect	256	146	257	147
rect	256	156	257	157
rect	256	162	257	163
rect	256	166	257	167
rect	257	7	258	8
rect	257	14	258	15
rect	257	17	258	18
rect	257	20	258	21
rect	257	23	258	24
rect	257	26	258	27
rect	257	33	258	34
rect	257	36	258	37
rect	257	39	258	40
rect	257	42	258	43
rect	257	45	258	46
rect	257	48	258	49
rect	257	51	258	52
rect	257	54	258	55
rect	257	64	258	65
rect	257	67	258	68
rect	257	70	258	71
rect	257	73	258	74
rect	257	76	258	77
rect	257	79	258	80
rect	257	83	258	84
rect	257	86	258	87
rect	257	99	258	100
rect	257	102	258	103
rect	257	106	258	107
rect	257	108	258	109
rect	257	126	258	127
rect	257	129	258	130
rect	257	133	258	134
rect	257	162	258	163
rect	258	7	259	8
rect	258	14	259	15
rect	258	17	259	18
rect	258	20	259	21
rect	258	23	259	24
rect	258	26	259	27
rect	258	33	259	34
rect	258	36	259	37
rect	258	39	259	40
rect	258	42	259	43
rect	258	45	259	46
rect	258	48	259	49
rect	258	51	259	52
rect	258	54	259	55
rect	258	57	259	58
rect	258	64	259	65
rect	258	67	259	68
rect	258	70	259	71
rect	258	73	259	74
rect	258	76	259	77
rect	258	79	259	80
rect	258	83	259	84
rect	258	86	259	87
rect	258	99	259	100
rect	258	102	259	103
rect	258	106	259	107
rect	258	108	259	109
rect	258	126	259	127
rect	258	129	259	130
rect	258	133	259	134
rect	258	139	259	140
rect	258	162	259	163
rect	259	7	260	8
rect	259	17	260	18
rect	259	20	260	21
rect	259	23	260	24
rect	259	26	260	27
rect	259	33	260	34
rect	259	36	260	37
rect	259	39	260	40
rect	259	42	260	43
rect	259	45	260	46
rect	259	48	260	49
rect	259	51	260	52
rect	259	54	260	55
rect	259	57	260	58
rect	259	64	260	65
rect	259	67	260	68
rect	259	70	260	71
rect	259	73	260	74
rect	259	76	260	77
rect	259	83	260	84
rect	259	86	260	87
rect	259	99	260	100
rect	259	102	260	103
rect	259	106	260	107
rect	259	126	260	127
rect	259	129	260	130
rect	259	133	260	134
rect	259	139	260	140
rect	260	7	261	8
rect	260	17	261	18
rect	260	20	261	21
rect	260	23	261	24
rect	260	26	261	27
rect	260	30	261	31
rect	260	33	261	34
rect	260	36	261	37
rect	260	39	261	40
rect	260	42	261	43
rect	260	45	261	46
rect	260	48	261	49
rect	260	51	261	52
rect	260	54	261	55
rect	260	57	261	58
rect	260	60	261	61
rect	260	64	261	65
rect	260	67	261	68
rect	260	70	261	71
rect	260	73	261	74
rect	260	76	261	77
rect	260	83	261	84
rect	260	86	261	87
rect	260	89	261	90
rect	260	99	261	100
rect	260	102	261	103
rect	260	106	261	107
rect	260	112	261	113
rect	260	126	261	127
rect	260	129	261	130
rect	260	133	261	134
rect	260	139	261	140
rect	267	4	268	5
rect	267	7	268	8
rect	267	11	268	12
rect	267	17	268	18
rect	267	20	268	21
rect	267	23	268	24
rect	267	26	268	27
rect	267	30	268	31
rect	267	33	268	34
rect	267	36	268	37
rect	267	39	268	40
rect	267	42	268	43
rect	267	45	268	46
rect	267	48	268	49
rect	267	51	268	52
rect	267	54	268	55
rect	267	57	268	58
rect	267	60	268	61
rect	267	64	268	65
rect	267	67	268	68
rect	267	70	268	71
rect	267	73	268	74
rect	267	76	268	77
rect	267	80	268	81
rect	267	83	268	84
rect	267	86	268	87
rect	267	89	268	90
rect	267	99	268	100
rect	267	102	268	103
rect	267	112	268	113
rect	267	116	268	117
rect	267	119	268	120
rect	267	126	268	127
rect	267	129	268	130
rect	267	139	268	140
rect	268	4	269	5
rect	268	7	269	8
rect	268	11	269	12
rect	268	17	269	18
rect	268	20	269	21
rect	268	23	269	24
rect	268	26	269	27
rect	268	30	269	31
rect	268	33	269	34
rect	268	36	269	37
rect	268	39	269	40
rect	268	42	269	43
rect	268	45	269	46
rect	268	48	269	49
rect	268	51	269	52
rect	268	57	269	58
rect	268	60	269	61
rect	268	64	269	65
rect	268	67	269	68
rect	268	70	269	71
rect	268	73	269	74
rect	268	76	269	77
rect	268	80	269	81
rect	268	83	269	84
rect	268	86	269	87
rect	268	89	269	90
rect	268	99	269	100
rect	268	102	269	103
rect	268	112	269	113
rect	268	116	269	117
rect	268	119	269	120
rect	268	126	269	127
rect	268	129	269	130
rect	268	139	269	140
rect	269	4	270	5
rect	269	7	270	8
rect	269	11	270	12
rect	269	17	270	18
rect	269	20	270	21
rect	269	23	270	24
rect	269	26	270	27
rect	269	28	270	29
rect	269	30	270	31
rect	269	33	270	34
rect	269	36	270	37
rect	269	39	270	40
rect	269	42	270	43
rect	269	45	270	46
rect	269	48	270	49
rect	269	51	270	52
rect	269	57	270	58
rect	269	60	270	61
rect	269	64	270	65
rect	269	67	270	68
rect	269	70	270	71
rect	269	73	270	74
rect	269	76	270	77
rect	269	80	270	81
rect	269	83	270	84
rect	269	86	270	87
rect	269	89	270	90
rect	269	99	270	100
rect	269	102	270	103
rect	269	112	270	113
rect	269	116	270	117
rect	269	119	270	120
rect	269	126	270	127
rect	269	129	270	130
rect	269	139	270	140
rect	270	4	271	5
rect	270	7	271	8
rect	270	11	271	12
rect	270	17	271	18
rect	270	20	271	21
rect	270	23	271	24
rect	270	26	271	27
rect	270	28	271	29
rect	270	30	271	31
rect	270	36	271	37
rect	270	39	271	40
rect	270	42	271	43
rect	270	45	271	46
rect	270	48	271	49
rect	270	57	271	58
rect	270	64	271	65
rect	270	67	271	68
rect	270	70	271	71
rect	270	73	271	74
rect	270	76	271	77
rect	270	80	271	81
rect	270	83	271	84
rect	270	86	271	87
rect	270	89	271	90
rect	270	99	271	100
rect	270	102	271	103
rect	270	112	271	113
rect	270	116	271	117
rect	270	119	271	120
rect	270	126	271	127
rect	270	129	271	130
rect	270	139	271	140
rect	271	4	272	5
rect	271	7	272	8
rect	271	11	272	12
rect	271	17	272	18
rect	271	20	272	21
rect	271	23	272	24
rect	271	26	272	27
rect	271	28	272	29
rect	271	30	272	31
rect	271	36	272	37
rect	271	39	272	40
rect	271	42	272	43
rect	271	45	272	46
rect	271	48	272	49
rect	271	55	272	56
rect	271	57	272	58
rect	271	64	272	65
rect	271	67	272	68
rect	271	70	272	71
rect	271	73	272	74
rect	271	76	272	77
rect	271	80	272	81
rect	271	83	272	84
rect	271	86	272	87
rect	271	89	272	90
rect	271	99	272	100
rect	271	102	272	103
rect	271	112	272	113
rect	271	116	272	117
rect	271	119	272	120
rect	271	126	272	127
rect	271	129	272	130
rect	271	139	272	140
rect	272	4	273	5
rect	272	7	273	8
rect	272	11	273	12
rect	272	17	273	18
rect	272	20	273	21
rect	272	23	273	24
rect	272	26	273	27
rect	272	28	273	29
rect	272	30	273	31
rect	272	36	273	37
rect	272	39	273	40
rect	272	42	273	43
rect	272	45	273	46
rect	272	48	273	49
rect	272	55	273	56
rect	272	57	273	58
rect	272	64	273	65
rect	272	67	273	68
rect	272	70	273	71
rect	272	73	273	74
rect	272	80	273	81
rect	272	83	273	84
rect	272	86	273	87
rect	272	89	273	90
rect	272	99	273	100
rect	272	102	273	103
rect	272	112	273	113
rect	272	116	273	117
rect	272	119	273	120
rect	272	126	273	127
rect	272	129	273	130
rect	272	139	273	140
rect	273	4	274	5
rect	273	7	274	8
rect	273	11	274	12
rect	273	17	274	18
rect	273	20	274	21
rect	273	23	274	24
rect	273	26	274	27
rect	273	28	274	29
rect	273	30	274	31
rect	273	36	274	37
rect	273	39	274	40
rect	273	42	274	43
rect	273	45	274	46
rect	273	48	274	49
rect	273	52	274	53
rect	273	55	274	56
rect	273	57	274	58
rect	273	64	274	65
rect	273	67	274	68
rect	273	70	274	71
rect	273	73	274	74
rect	273	80	274	81
rect	273	83	274	84
rect	273	86	274	87
rect	273	89	274	90
rect	273	99	274	100
rect	273	102	274	103
rect	273	112	274	113
rect	273	116	274	117
rect	273	119	274	120
rect	273	126	274	127
rect	273	129	274	130
rect	273	139	274	140
rect	274	4	275	5
rect	274	7	275	8
rect	274	11	275	12
rect	274	17	275	18
rect	274	20	275	21
rect	274	23	275	24
rect	274	26	275	27
rect	274	28	275	29
rect	274	30	275	31
rect	274	36	275	37
rect	274	39	275	40
rect	274	42	275	43
rect	274	45	275	46
rect	274	52	275	53
rect	274	55	275	56
rect	274	57	275	58
rect	274	67	275	68
rect	274	70	275	71
rect	274	73	275	74
rect	274	83	275	84
rect	274	89	275	90
rect	274	99	275	100
rect	274	102	275	103
rect	274	112	275	113
rect	274	116	275	117
rect	274	119	275	120
rect	274	126	275	127
rect	274	129	275	130
rect	274	139	275	140
rect	275	4	276	5
rect	275	7	276	8
rect	275	11	276	12
rect	275	17	276	18
rect	275	20	276	21
rect	275	23	276	24
rect	275	26	276	27
rect	275	28	276	29
rect	275	30	276	31
rect	275	36	276	37
rect	275	39	276	40
rect	275	42	276	43
rect	275	45	276	46
rect	275	52	276	53
rect	275	55	276	56
rect	275	57	276	58
rect	275	67	276	68
rect	275	70	276	71
rect	275	73	276	74
rect	275	83	276	84
rect	275	89	276	90
rect	275	99	276	100
rect	275	102	276	103
rect	275	112	276	113
rect	275	116	276	117
rect	275	119	276	120
rect	275	126	276	127
rect	275	129	276	130
rect	275	139	276	140
rect	276	4	277	5
rect	276	7	277	8
rect	276	17	277	18
rect	276	23	277	24
rect	276	28	277	29
rect	276	30	277	31
rect	276	36	277	37
rect	276	39	277	40
rect	276	42	277	43
rect	276	45	277	46
rect	276	52	277	53
rect	276	55	277	56
rect	276	57	277	58
rect	276	67	277	68
rect	276	70	277	71
rect	276	73	277	74
rect	276	83	277	84
rect	276	89	277	90
rect	276	102	277	103
rect	276	112	277	113
rect	276	116	277	117
rect	276	119	277	120
rect	276	126	277	127
rect	276	129	277	130
rect	276	139	277	140
rect	277	4	278	5
rect	277	7	278	8
rect	277	17	278	18
rect	277	23	278	24
rect	277	25	278	26
rect	277	28	278	29
rect	277	30	278	31
rect	277	36	278	37
rect	277	39	278	40
rect	277	42	278	43
rect	277	45	278	46
rect	277	49	278	50
rect	277	52	278	53
rect	277	55	278	56
rect	277	57	278	58
rect	277	67	278	68
rect	277	70	278	71
rect	277	73	278	74
rect	277	83	278	84
rect	277	89	278	90
rect	277	102	278	103
rect	277	112	278	113
rect	277	116	278	117
rect	277	119	278	120
rect	277	126	278	127
rect	277	129	278	130
rect	277	139	278	140
rect	278	4	279	5
rect	278	7	279	8
rect	278	23	279	24
rect	278	25	279	26
rect	278	28	279	29
rect	278	30	279	31
rect	278	36	279	37
rect	278	42	279	43
rect	278	49	279	50
rect	278	52	279	53
rect	278	55	279	56
rect	278	57	279	58
rect	278	70	279	71
rect	278	89	279	90
rect	278	102	279	103
rect	278	112	279	113
rect	278	116	279	117
rect	278	119	279	120
rect	278	126	279	127
rect	278	129	279	130
rect	278	139	279	140
rect	279	4	280	5
rect	279	7	280	8
rect	279	11	280	12
rect	279	21	280	22
rect	279	23	280	24
rect	279	25	280	26
rect	279	28	280	29
rect	279	30	280	31
rect	279	36	280	37
rect	279	42	280	43
rect	279	49	280	50
rect	279	52	280	53
rect	279	55	280	56
rect	279	57	280	58
rect	279	70	280	71
rect	279	89	280	90
rect	279	102	280	103
rect	279	112	280	113
rect	279	116	280	117
rect	279	119	280	120
rect	279	126	280	127
rect	279	129	280	130
rect	279	139	280	140
rect	280	4	281	5
rect	280	7	281	8
rect	280	11	281	12
rect	280	21	281	22
rect	280	23	281	24
rect	280	25	281	26
rect	280	28	281	29
rect	280	30	281	31
rect	280	42	281	43
rect	280	49	281	50
rect	280	52	281	53
rect	280	55	281	56
rect	280	57	281	58
rect	280	89	281	90
rect	280	112	281	113
rect	280	119	281	120
rect	280	126	281	127
rect	280	139	281	140
rect	281	4	282	5
rect	281	7	282	8
rect	281	11	282	12
rect	281	18	282	19
rect	281	21	282	22
rect	281	23	282	24
rect	281	25	282	26
rect	281	28	282	29
rect	281	30	282	31
rect	281	39	282	40
rect	281	42	282	43
rect	281	49	282	50
rect	281	52	282	53
rect	281	55	282	56
rect	281	57	282	58
rect	281	73	282	74
rect	281	89	282	90
rect	281	112	282	113
rect	281	119	282	120
rect	281	126	282	127
rect	281	139	282	140
rect	282	11	283	12
rect	282	18	283	19
rect	282	21	283	22
rect	282	25	283	26
rect	282	28	283	29
rect	282	39	283	40
rect	282	49	283	50
rect	282	52	283	53
rect	282	55	283	56
rect	282	73	283	74
rect	283	11	284	12
rect	283	14	284	15
rect	283	18	284	19
rect	283	21	284	22
rect	283	25	284	26
rect	283	28	284	29
rect	283	39	284	40
rect	283	45	284	46
rect	283	49	284	50
rect	283	52	284	53
rect	283	55	284	56
rect	283	62	284	63
rect	283	73	284	74
rect	290	8	291	9
rect	290	11	291	12
rect	290	14	291	15
rect	290	39	291	40
rect	290	45	291	46
rect	290	55	291	56
rect	290	59	291	60
rect	290	73	291	74
rect	291	8	292	9
rect	291	73	292	74
rect	292	8	293	9
rect	292	73	293	74
<< via >>
rect	0	40	1	41
rect	0	46	1	47
rect	2	37	3	38
rect	2	43	3	44
rect	2	63	3	64
rect	2	73	3	74
rect	2	83	3	84
rect	2	87	3	88
rect	2	90	3	91
rect	2	93	3	94
rect	4	4	5	5
rect	4	10	5	11
rect	4	33	5	34
rect	4	50	5	51
rect	4	60	5	61
rect	4	66	5	67
rect	4	77	5	78
rect	4	103	5	104
rect	6	1	7	2
rect	6	7	7	8
rect	6	17	7	18
rect	6	20	7	21
rect	6	23	7	24
rect	6	97	7	98
rect	8	16	9	17
rect	8	17	9	18
rect	8	19	9	20
rect	8	20	9	21
rect	8	22	9	23
rect	8	23	9	24
rect	8	25	9	26
rect	8	26	9	27
rect	8	34	9	35
rect	8	35	9	36
rect	8	53	9	54
rect	8	54	9	55
rect	8	58	9	59
rect	8	59	9	60
rect	8	72	9	73
rect	8	73	9	74
rect	8	74	9	75
rect	8	75	9	76
rect	8	80	9	81
rect	8	81	9	82
rect	8	83	9	84
rect	8	84	9	85
rect	15	50	16	51
rect	15	71	16	72
rect	17	43	18	44
rect	17	55	18	56
rect	17	77	18	78
rect	17	115	18	116
rect	19	7	20	8
rect	19	17	20	18
rect	19	39	20	40
rect	19	77	20	78
rect	19	93	20	94
rect	19	112	20	113
rect	21	29	22	30
rect	21	33	22	34
rect	21	37	22	38
rect	21	52	22	53
rect	21	93	22	94
rect	21	139	22	140
rect	23	10	24	11
rect	23	14	24	15
rect	23	27	24	28
rect	23	42	24	43
rect	23	46	24	47
rect	23	58	24	59
rect	23	61	24	62
rect	23	63	24	64
rect	23	68	24	69
rect	23	96	24	97
rect	23	99	24	100
rect	23	100	24	101
rect	23	103	24	104
rect	23	142	24	143
rect	25	14	26	15
rect	25	102	26	103
rect	27	1	28	2
rect	27	4	28	5
rect	27	11	28	12
rect	27	49	28	50
rect	27	64	28	65
rect	27	66	28	67
rect	27	80	28	81
rect	27	83	28	84
rect	27	87	28	88
rect	27	132	28	133
rect	29	4	30	5
rect	29	32	30	33
rect	29	36	30	37
rect	29	80	30	81
rect	29	87	30	88
rect	29	126	30	127
rect	38	58	39	59
rect	38	70	39	71
rect	40	68	41	69
rect	42	55	43	56
rect	42	67	43	68
rect	42	90	43	91
rect	42	93	43	94
rect	42	102	43	103
rect	42	108	43	109
rect	44	10	45	11
rect	44	29	45	30
rect	44	45	45	46
rect	44	61	45	62
rect	44	77	45	78
rect	44	89	45	90
rect	44	99	45	100
rect	44	105	45	106
rect	46	7	47	8
rect	46	29	47	30
rect	46	52	47	53
rect	46	61	47	62
rect	46	64	47	65
rect	46	76	47	77
rect	46	92	47	93
rect	46	96	47	97
rect	46	122	47	123
rect	46	137	47	138
rect	46	142	47	143
rect	46	147	47	148
rect	46	157	47	158
rect	48	7	49	8
rect	48	39	49	40
rect	48	166	49	167
rect	50	32	51	33
rect	50	39	51	40
rect	50	42	51	43
rect	50	64	51	65
rect	50	102	51	103
rect	50	112	51	113
rect	50	124	51	125
rect	50	132	51	133
rect	50	160	51	161
rect	52	14	53	15
rect	52	33	53	34
rect	52	42	53	43
rect	52	49	53	50
rect	52	55	53	56
rect	52	73	53	74
rect	52	83	53	84
rect	52	86	53	87
rect	52	96	53	97
rect	52	99	53	100
rect	52	163	53	164
rect	54	4	55	5
rect	54	13	55	14
rect	54	20	55	21
rect	54	111	55	112
rect	54	115	55	116
rect	54	121	55	122
rect	54	129	55	130
rect	54	134	55	135
rect	54	141	55	142
rect	54	150	55	151
rect	63	166	64	167
rect	63	178	64	179
rect	65	115	66	116
rect	65	166	66	167
rect	67	111	68	112
rect	67	115	68	116
rect	69	108	70	109
rect	69	112	70	113
rect	69	154	70	155
rect	69	208	70	209
rect	71	61	72	62
rect	71	105	72	106
rect	71	109	72	110
rect	71	134	72	135
rect	71	153	72	154
rect	73	76	74	77
rect	73	83	74	84
rect	73	102	74	103
rect	73	134	74	135
rect	75	73	76	74
rect	75	80	76	81
rect	75	92	76	93
rect	75	106	76	107
rect	75	124	76	125
rect	75	140	76	141
rect	75	147	76	148
rect	75	156	76	157
rect	77	70	78	71
rect	77	77	78	78
rect	77	89	78	90
rect	77	103	78	104
rect	77	125	78	126
rect	77	147	78	148
rect	79	67	80	68
rect	79	86	80	87
rect	79	93	80	94
rect	79	97	80	98
rect	79	169	80	170
rect	81	17	82	18
rect	81	29	82	30
rect	81	42	82	43
rect	81	52	82	53
rect	81	64	82	65
rect	81	68	82	69
rect	81	71	82	72
rect	81	128	82	129
rect	83	29	84	30
rect	83	39	84	40
rect	83	49	84	50
rect	83	58	84	59
rect	83	100	84	101
rect	83	121	84	122
rect	83	128	84	129
rect	83	163	84	164
rect	83	172	84	173
rect	85	1	86	2
rect	85	10	86	11
rect	85	13	86	14
rect	85	26	86	27
rect	85	36	86	37
rect	85	39	86	40
rect	85	42	86	43
rect	85	45	86	46
rect	85	55	86	56
rect	85	62	86	63
rect	85	65	86	66
rect	85	163	86	164
rect	87	4	88	5
rect	87	7	88	8
rect	87	11	88	12
rect	87	14	88	15
rect	87	33	88	34
rect	87	131	88	132
rect	87	160	88	161
rect	87	175	88	176
rect	102	39	103	40
rect	102	100	103	101
rect	102	122	103	123
rect	102	128	103	129
rect	104	38	105	39
rect	104	87	105	88
rect	104	90	105	91
rect	104	100	105	101
rect	104	109	105	110
rect	104	129	105	130
rect	106	47	107	48
rect	106	65	107	66
rect	106	68	107	69
rect	106	88	107	89
rect	106	110	107	111
rect	106	125	107	126
rect	108	66	109	67
rect	108	93	109	94
rect	108	126	109	127
rect	108	131	109	132
rect	108	147	109	148
rect	108	150	109	151
rect	110	62	111	63
rect	110	196	111	197
rect	112	31	113	32
rect	112	60	113	61
rect	112	63	113	64
rect	112	71	113	72
rect	112	77	113	78
rect	112	97	113	98
rect	112	103	113	104
rect	112	119	113	120
rect	112	132	113	133
rect	112	156	113	157
rect	114	20	115	21
rect	114	33	115	34
rect	114	42	115	43
rect	114	57	115	58
rect	114	91	115	92
rect	114	97	115	98
rect	114	106	115	107
rect	114	115	115	116
rect	114	116	115	117
rect	114	134	115	135
rect	114	144	115	145
rect	114	148	115	149
rect	114	153	115	154
rect	114	157	115	158
rect	114	175	115	176
rect	116	29	117	30
rect	116	72	117	73
rect	116	83	117	84
rect	116	84	117	85
rect	116	94	117	95
rect	116	104	117	105
rect	116	112	117	113
rect	116	113	117	114
rect	116	135	117	136
rect	116	137	117	138
rect	116	142	117	143
rect	116	151	117	152
rect	116	172	117	173
rect	116	176	117	177
rect	118	14	119	15
rect	118	28	119	29
rect	118	52	119	53
rect	118	120	119	121
rect	118	138	119	139
rect	118	140	119	141
rect	118	154	119	155
rect	118	166	119	167
rect	118	169	119	170
rect	118	173	119	174
rect	120	4	121	5
rect	120	41	121	42
rect	120	44	121	45
rect	120	51	121	52
rect	120	69	121	70
rect	120	78	121	79
rect	120	160	121	161
rect	120	164	121	165
rect	120	170	121	171
rect	120	178	121	179
rect	120	182	121	183
rect	122	1	123	2
rect	122	7	123	8
rect	122	11	123	12
rect	122	13	123	14
rect	122	23	123	24
rect	122	193	123	194
rect	124	1	125	2
rect	124	10	125	11
rect	124	145	125	146
rect	124	161	125	162
rect	124	167	125	168
rect	124	179	125	180
rect	124	208	125	209
rect	139	97	140	98
rect	139	104	140	105
rect	141	57	142	58
rect	141	97	142	98
rect	143	56	144	57
rect	143	78	144	79
rect	145	78	146	79
rect	145	88	146	89
rect	147	75	148	76
rect	147	90	148	91
rect	149	72	150	73
rect	149	87	150	88
rect	149	106	150	107
rect	149	113	150	114
rect	149	116	150	117
rect	149	119	150	120
rect	151	63	152	64
rect	151	75	152	76
rect	151	113	152	114
rect	151	132	152	133
rect	151	167	152	168
rect	151	196	152	197
rect	153	62	154	63
rect	153	84	154	85
rect	153	100	154	101
rect	153	116	154	117
rect	153	167	154	168
rect	153	182	154	183
rect	155	41	156	42
rect	155	72	156	73
rect	155	94	156	95
rect	155	100	156	101
rect	155	132	156	133
rect	155	135	156	136
rect	155	145	156	146
rect	155	148	156	149
rect	155	176	156	177
rect	155	183	156	184
rect	157	7	158	8
rect	157	38	158	39
rect	157	47	158	48
rect	157	50	158	51
rect	157	69	158	70
rect	157	84	158	85
rect	157	177	158	178
rect	159	7	160	8
rect	159	31	160	32
rect	159	41	160	42
rect	159	47	160	48
rect	159	60	160	61
rect	159	81	160	82
rect	159	161	160	162
rect	161	4	162	5
rect	161	10	162	11
rect	161	13	162	14
rect	161	32	162	33
rect	161	103	162	104
rect	161	135	162	136
rect	161	138	162	139
rect	161	148	162	149
rect	161	151	162	152
rect	163	10	164	11
rect	163	28	164	29
rect	163	66	164	67
rect	163	81	164	82
rect	163	193	164	194
rect	165	4	166	5
rect	165	151	166	152
rect	165	154	166	155
rect	165	164	166	165
rect	165	170	166	171
rect	165	186	166	187
rect	167	1	168	2
rect	167	110	168	111
rect	167	126	168	127
rect	167	145	168	146
rect	167	154	168	155
rect	167	179	168	180
rect	169	1	170	2
rect	169	13	170	14
rect	169	22	170	23
rect	169	123	170	124
rect	169	126	170	127
rect	169	170	170	171
rect	169	173	170	174
rect	169	180	170	181
rect	194	64	195	65
rect	194	75	195	76
rect	196	76	197	77
rect	196	90	197	91
rect	198	67	199	68
rect	198	78	199	79
rect	198	94	199	95
rect	198	100	199	101
rect	200	62	201	63
rect	200	79	201	80
rect	200	92	201	93
rect	200	106	201	107
rect	202	61	203	62
rect	202	116	203	117
rect	202	121	203	122
rect	202	132	203	133
rect	204	29	205	30
rect	204	38	205	39
rect	204	44	205	45
rect	204	131	205	132
rect	204	145	205	146
rect	204	164	205	165
rect	206	39	207	40
rect	206	41	207	42
rect	206	45	207	46
rect	206	50	207	51
rect	206	69	207	70
rect	206	99	207	100
rect	206	105	207	106
rect	206	115	207	116
rect	206	146	207	147
rect	206	157	207	158
rect	208	32	209	33
rect	208	35	209	36
rect	208	42	209	43
rect	208	123	209	124
rect	208	127	209	128
rect	208	135	209	136
rect	208	143	209	144
rect	208	154	209	155
rect	210	29	211	30
rect	210	47	211	48
rect	210	51	211	52
rect	210	56	211	57
rect	210	70	211	71
rect	210	81	211	82
rect	210	89	211	90
rect	210	103	211	104
rect	210	108	211	109
rect	210	119	211	120
rect	210	124	211	125
rect	210	148	211	149
rect	210	153	211	154
rect	210	159	211	160
rect	212	4	213	5
rect	212	7	213	8
rect	212	25	213	26
rect	212	33	213	34
rect	212	48	213	49
rect	212	87	213	88
rect	212	95	213	96
rect	212	134	213	135
rect	212	140	213	141
rect	212	151	213	152
rect	212	162	213	163
rect	212	170	213	171
rect	214	8	215	9
rect	214	169	215	170
rect	216	1	217	2
rect	216	156	217	157
rect	216	183	217	184
rect	216	190	217	191
rect	218	1	219	2
rect	218	10	219	11
rect	218	13	219	14
rect	218	14	219	15
rect	218	26	219	27
rect	218	112	219	113
rect	218	118	219	119
rect	218	129	219	130
rect	218	137	219	138
rect	218	167	219	168
rect	218	180	219	181
rect	218	187	219	188
rect	233	33	234	34
rect	233	105	234	106
rect	235	33	236	34
rect	235	42	236	43
rect	237	42	238	43
rect	237	73	238	74
rect	239	54	240	55
rect	239	58	240	59
rect	239	73	240	74
rect	239	86	240	87
rect	241	20	242	21
rect	241	61	242	62
rect	241	64	242	65
rect	241	83	242	84
rect	243	20	244	21
rect	243	51	244	52
rect	243	54	244	55
rect	243	134	244	135
rect	245	51	246	52
rect	245	76	246	77
rect	247	39	248	40
rect	247	64	248	65
rect	247	86	248	87
rect	247	102	248	103
rect	247	129	248	130
rect	247	159	248	160
rect	249	39	250	40
rect	249	70	250	71
rect	249	76	250	77
rect	249	95	250	96
rect	249	127	250	128
rect	249	133	250	134
rect	251	7	252	8
rect	251	17	252	18
rect	251	36	252	37
rect	251	67	252	68
rect	251	70	252	71
rect	251	92	252	93
rect	251	106	252	107
rect	251	118	252	119
rect	251	126	252	127
rect	251	143	252	144
rect	253	17	254	18
rect	253	99	254	100
rect	253	102	254	103
rect	253	140	254	141
rect	255	67	256	68
rect	255	89	256	90
rect	255	99	256	100
rect	255	137	256	138
rect	257	4	258	5
rect	257	29	258	30
rect	257	57	258	58
rect	257	112	258	113
rect	257	115	258	116
rect	257	121	258	122
rect	257	124	258	125
rect	257	131	258	132
rect	257	139	258	140
rect	257	146	258	147
rect	257	156	258	157
rect	257	166	258	167
rect	259	14	260	15
rect	259	30	260	31
rect	259	60	260	61
rect	259	79	260	80
rect	259	89	260	90
rect	259	108	260	109
rect	259	112	260	113
rect	259	162	260	163
rect	268	28	269	29
rect	268	54	269	55
rect	270	33	271	34
rect	270	51	271	52
rect	270	55	271	56
rect	270	60	271	61
rect	272	52	273	53
rect	272	76	273	77
rect	274	48	275	49
rect	274	64	275	65
rect	274	80	275	81
rect	274	86	275	87
rect	276	11	277	12
rect	276	20	277	21
rect	276	25	277	26
rect	276	26	277	27
rect	276	49	277	50
rect	276	99	277	100
rect	278	11	279	12
rect	278	17	279	18
rect	278	21	279	22
rect	278	39	279	40
rect	278	45	279	46
rect	278	67	279	68
rect	278	73	279	74
rect	278	83	279	84
rect	280	18	281	19
rect	280	36	281	37
rect	280	39	281	40
rect	280	70	281	71
rect	280	73	281	74
rect	280	102	281	103
rect	280	116	281	117
rect	280	129	281	130
rect	282	4	283	5
rect	282	7	283	8
rect	282	14	283	15
rect	282	23	283	24
rect	282	30	283	31
rect	282	42	283	43
rect	282	45	283	46
rect	282	57	283	58
rect	282	62	283	63
rect	282	89	283	90
rect	282	112	283	113
rect	282	119	283	120
rect	282	126	283	127
rect	282	139	283	140
rect	291	11	292	12
rect	291	14	292	15
rect	291	39	292	40
rect	291	45	292	46
rect	291	55	292	56
rect	291	59	292	60
rect	293	8	294	9
rect	293	73	294	74
