magic
tech scmos
timestamp
<< pdiffusion >>
rect	0	5	6	11
rect	0	33	6	39
rect	17	5	23	11
rect	56	33	62	39
rect	0	19	6	25
rect	0	49	6	55
rect	29	19	35	25
rect	20	49	26	55
rect	10	5	16	11
rect	31	33	37	39
rect	27	5	33	11
rect	78	33	84	39
rect	13	19	19	25
rect	10	49	16	55
rect	54	19	60	25
rect	27	49	33	55
rect	0	12	6	18
rect	0	40	6	46
rect	17	12	23	18
rect	35	40	41	46
rect	0	26	6	32
rect	3	56	9	62
rect	35	26	41	32
rect	37	5	43	11
rect	94	33	100	39
rect	60	5	66	11
rect	123	33	129	39
rect	82	19	88	25
rect	37	49	43	55
rect	105	19	111	25
rect	51	49	57	55
rect	47	5	53	11
rect	107	33	113	39
rect	73	5	79	11
rect	130	33	136	39
rect	95	19	101	25
rect	44	49	50	55
rect	112	19	118	25
rect	67	49	73	55
rect	46	12	52	18
rect	82	40	88	46
rect	75	12	81	18
rect	105	40	111	46
rect	67	26	73	32
rect	31	56	37	62
rect	65	12	68	18
rect	6	19	9	25
rect	23	12	26	18
rect	111	40	114	46
rect	6	5	9	11
rect	9	19	12	25
rect	55	40	58	46
rect	41	40	44	46
rect	66	5	69	11
rect	57	49	60	55
rect	53	5	56	11
rect	113	33	116	39
rect	101	40	104	46
rect	31	12	34	18
rect	41	26	44	32
rect	60	19	63	25
rect	116	33	119	39
rect	6	33	9	39
rect	19	19	22	25
rect	23	5	26	11
rect	44	26	47	32
rect	16	49	19	55
rect	88	19	91	25
rect	127	26	130	32
rect	26	12	29	18
rect	14	40	17	46
rect	34	12	37	18
rect	37	33	40	39
rect	33	5	36	11
rect	59	40	62	46
rect	28	40	31	46
rect	100	33	103	39
rect	40	33	43	39
rect	0	56	3	62
rect	69	40	72	46
rect	62	40	65	46
rect	9	33	12	39
rect	33	49	36	55
rect	31	40	34	46
rect	56	5	59	11
rect	6	49	9	55
rect	91	19	94	25
rect	63	19	66	25
rect	66	19	69	25
rect	10	26	13	32
rect	22	19	25	25
rect	136	33	139	39
rect	7	12	10	18
rect	13	26	16	32
rect	62	33	65	39
rect	65	33	68	39
rect	68	12	71	18
rect	88	40	91	46
rect	93	40	96	46
rect	119	33	122	39
rect	35	19	38	25
rect	73	26	76	32
rect	117	26	120	32
rect	7	40	10	46
rect	38	19	41	25
rect	23	40	26	46
rect	107	26	110	32
rect	41	19	44	25
rect	12	33	15	39
rect	44	19	47	25
rect	84	33	87	39
rect	15	33	18	39
rect	72	40	75	46
rect	87	33	90	39
rect	16	26	19	32
rect	44	40	47	46
rect	43	33	46	39
rect	60	12	63	18
rect	10	40	13	46
rect	113	26	116	32
rect	88	26	91	32
rect	91	26	94	32
rect	18	33	21	39
rect	47	26	50	32
rect	140	26	143	32
rect	21	33	24	39
rect	76	26	79	32
rect	69	19	72	25
rect	90	33	93	39
rect	91	49	94	55
rect	123	26	126	32
rect	101	19	104	25
rect	24	33	27	39
rect	57	26	60	32
rect	19	26	22	32
rect	79	26	82	32
rect	6	26	9	32
rect	60	49	63	55
rect	46	33	49	39
rect	50	26	53	32
rect	72	19	75	25
rect	27	33	30	39
rect	103	33	106	39
rect	68	33	71	39
rect	71	33	74	39
rect	19	40	22	46
rect	49	33	52	39
rect	75	19	78	25
rect	82	26	85	32
rect	94	26	97	32
rect	127	19	130	25
rect	102	12	105	18
rect	25	26	28	32
rect	52	33	55	39
rect	25	19	28	25
rect	53	26	56	32
rect	78	19	81	25
rect	28	26	31	32
rect	75	40	78	46
rect	78	40	81	46
rect	50	40	53	46
rect	71	12	74	18
rect	74	33	77	39
rect	131	12	134	18
rect	47	19	50	25
rect	82	12	85	18
rect	50	19	53	25
rect	76	49	79	55
rect	79	49	82	55
rect	69	5	72	11
rect	65	40	68	46
rect	52	12	55	18
rect	42	12	45	18
rect	77	56	80	62
rect	63	49	66	55
rect	43	5	46	11
