magic
tech scmos
timestamp
<< pdiffusion >>
rect	6	0	7	1
rect	6	1	7	2
rect	6	2	7	3
rect	6	3	7	4
rect	6	4	7	5
rect	6	5	7	6
rect	6	6	7	7
rect	6	7	7	8
rect	6	8	7	9
rect	6	9	7	10
rect	6	10	7	11
rect	6	11	7	12
rect	6	12	7	13
rect	6	13	7	14
rect	6	14	7	15
rect	6	15	7	16
rect	6	16	7	17
rect	6	17	7	18
rect	6	18	7	19
rect	6	19	7	20
rect	6	20	7	21
rect	6	21	7	22
rect	6	22	7	23
rect	6	23	7	24
rect	6	24	7	25
rect	6	25	7	26
rect	6	26	7	27
rect	6	27	7	28
rect	6	28	7	29
rect	6	29	7	30
rect	6	30	7	31
rect	6	31	7	32
rect	6	32	7	33
rect	6	33	7	34
rect	6	34	7	35
rect	6	35	7	36
rect	6	36	7	37
rect	6	37	7	38
rect	6	38	7	39
rect	6	39	7	40
rect	6	40	7	41
rect	6	41	7	42
rect	6	42	7	43
rect	6	43	7	44
rect	6	44	7	45
rect	6	45	7	46
rect	6	46	7	47
rect	6	47	7	48
rect	6	48	7	49
rect	6	49	7	50
rect	6	50	7	51
rect	6	51	7	52
rect	6	52	7	53
rect	6	53	7	54
rect	6	54	7	55
rect	6	55	7	56
rect	6	56	7	57
rect	6	57	7	58
rect	6	58	7	59
rect	6	59	7	60
rect	6	60	7	61
rect	6	61	7	62
rect	6	62	7	63
rect	6	63	7	64
rect	6	64	7	65
rect	6	65	7	66
rect	6	66	7	67
rect	6	67	7	68
rect	6	68	7	69
rect	6	69	7	70
rect	6	70	7	71
rect	6	71	7	72
rect	6	72	7	73
rect	6	73	7	74
rect	6	74	7	75
rect	6	75	7	76
rect	6	76	7	77
rect	6	77	7	78
rect	6	78	7	79
rect	6	79	7	80
rect	6	80	7	81
rect	6	81	7	82
rect	6	82	7	83
rect	6	83	7	84
rect	6	84	7	85
rect	6	85	7	86
rect	6	86	7	87
rect	6	87	7	88
rect	6	88	7	89
rect	6	89	7	90
rect	6	90	7	91
rect	6	91	7	92
rect	6	92	7	93
rect	6	93	7	94
rect	6	94	7	95
rect	6	95	7	96
rect	6	96	7	97
rect	6	97	7	98
rect	6	98	7	99
rect	6	99	7	100
rect	6	100	7	101
rect	6	101	7	102
rect	6	102	7	103
rect	6	103	7	104
rect	6	104	7	105
rect	6	105	7	106
rect	6	106	7	107
rect	6	107	7	108
rect	6	108	7	109
rect	6	109	7	110
rect	6	110	7	111
rect	6	111	7	112
rect	6	112	7	113
rect	6	113	7	114
rect	6	114	7	115
rect	6	115	7	116
rect	6	116	7	117
rect	6	117	7	118
rect	6	118	7	119
rect	6	119	7	120
rect	6	120	7	121
rect	6	121	7	122
rect	6	122	7	123
rect	6	123	7	124
rect	6	124	7	125
rect	6	125	7	126
rect	6	126	7	127
rect	6	127	7	128
rect	6	128	7	129
rect	6	129	7	130
rect	6	130	7	131
rect	6	131	7	132
rect	6	132	7	133
rect	6	133	7	134
rect	6	134	7	135
rect	6	135	7	136
rect	6	136	7	137
rect	6	137	7	138
rect	6	138	7	139
rect	6	139	7	140
rect	6	140	7	141
rect	6	141	7	142
rect	6	142	7	143
rect	6	143	7	144
rect	6	144	7	145
rect	6	145	7	146
rect	6	146	7	147
rect	6	147	7	148
rect	6	148	7	149
rect	6	149	7	150
rect	6	150	7	151
rect	6	151	7	152
rect	6	152	7	153
rect	6	153	7	154
rect	6	154	7	155
rect	6	155	7	156
rect	6	156	7	157
rect	6	157	7	158
rect	6	158	7	159
rect	6	159	7	160
rect	6	160	7	161
rect	6	161	7	162
rect	6	162	7	163
rect	6	163	7	164
rect	6	164	7	165
rect	6	165	7	166
rect	6	166	7	167
rect	6	167	7	168
rect	6	168	7	169
rect	6	169	7	170
rect	6	170	7	171
rect	6	171	7	172
rect	6	172	7	173
rect	6	173	7	174
rect	7	0	8	1
rect	7	1	8	2
rect	7	2	8	3
rect	7	3	8	4
rect	7	4	8	5
rect	7	5	8	6
rect	7	6	8	7
rect	7	7	8	8
rect	7	8	8	9
rect	7	9	8	10
rect	7	10	8	11
rect	7	11	8	12
rect	7	12	8	13
rect	7	13	8	14
rect	7	14	8	15
rect	7	15	8	16
rect	7	16	8	17
rect	7	17	8	18
rect	7	18	8	19
rect	7	19	8	20
rect	7	20	8	21
rect	7	21	8	22
rect	7	22	8	23
rect	7	23	8	24
rect	7	24	8	25
rect	7	25	8	26
rect	7	26	8	27
rect	7	27	8	28
rect	7	28	8	29
rect	7	29	8	30
rect	7	30	8	31
rect	7	31	8	32
rect	7	32	8	33
rect	7	33	8	34
rect	7	34	8	35
rect	7	35	8	36
rect	7	36	8	37
rect	7	37	8	38
rect	7	38	8	39
rect	7	39	8	40
rect	7	40	8	41
rect	7	41	8	42
rect	7	42	8	43
rect	7	43	8	44
rect	7	44	8	45
rect	7	45	8	46
rect	7	46	8	47
rect	7	47	8	48
rect	7	48	8	49
rect	7	49	8	50
rect	7	50	8	51
rect	7	51	8	52
rect	7	52	8	53
rect	7	53	8	54
rect	7	54	8	55
rect	7	55	8	56
rect	7	56	8	57
rect	7	57	8	58
rect	7	58	8	59
rect	7	59	8	60
rect	7	60	8	61
rect	7	61	8	62
rect	7	62	8	63
rect	7	63	8	64
rect	7	64	8	65
rect	7	65	8	66
rect	7	66	8	67
rect	7	67	8	68
rect	7	68	8	69
rect	7	69	8	70
rect	7	70	8	71
rect	7	71	8	72
rect	7	72	8	73
rect	7	73	8	74
rect	7	74	8	75
rect	7	75	8	76
rect	7	76	8	77
rect	7	77	8	78
rect	7	78	8	79
rect	7	79	8	80
rect	7	80	8	81
rect	7	81	8	82
rect	7	82	8	83
rect	7	83	8	84
rect	7	84	8	85
rect	7	85	8	86
rect	7	86	8	87
rect	7	87	8	88
rect	7	88	8	89
rect	7	89	8	90
rect	7	90	8	91
rect	7	91	8	92
rect	7	92	8	93
rect	7	93	8	94
rect	7	94	8	95
rect	7	95	8	96
rect	7	96	8	97
rect	7	97	8	98
rect	7	98	8	99
rect	7	99	8	100
rect	7	100	8	101
rect	7	101	8	102
rect	7	102	8	103
rect	7	103	8	104
rect	7	104	8	105
rect	7	105	8	106
rect	7	106	8	107
rect	7	107	8	108
rect	7	108	8	109
rect	7	109	8	110
rect	7	110	8	111
rect	7	111	8	112
rect	7	112	8	113
rect	7	113	8	114
rect	7	114	8	115
rect	7	115	8	116
rect	7	116	8	117
rect	7	117	8	118
rect	7	118	8	119
rect	7	119	8	120
rect	7	120	8	121
rect	7	121	8	122
rect	7	122	8	123
rect	7	123	8	124
rect	7	124	8	125
rect	7	125	8	126
rect	7	126	8	127
rect	7	127	8	128
rect	7	128	8	129
rect	7	129	8	130
rect	7	130	8	131
rect	7	131	8	132
rect	7	132	8	133
rect	7	133	8	134
rect	7	134	8	135
rect	7	135	8	136
rect	7	136	8	137
rect	7	137	8	138
rect	7	138	8	139
rect	7	139	8	140
rect	7	140	8	141
rect	7	141	8	142
rect	7	142	8	143
rect	7	143	8	144
rect	7	144	8	145
rect	7	145	8	146
rect	7	146	8	147
rect	7	147	8	148
rect	7	148	8	149
rect	7	149	8	150
rect	7	150	8	151
rect	7	151	8	152
rect	7	152	8	153
rect	7	153	8	154
rect	7	154	8	155
rect	7	155	8	156
rect	7	156	8	157
rect	7	157	8	158
rect	7	158	8	159
rect	7	159	8	160
rect	7	160	8	161
rect	7	161	8	162
rect	7	162	8	163
rect	7	163	8	164
rect	7	164	8	165
rect	7	165	8	166
rect	7	166	8	167
rect	7	167	8	168
rect	7	168	8	169
rect	7	169	8	170
rect	7	170	8	171
rect	7	171	8	172
rect	7	172	8	173
rect	7	173	8	174
rect	8	0	9	1
rect	8	1	9	2
rect	8	2	9	3
rect	8	3	9	4
rect	8	4	9	5
rect	8	5	9	6
rect	8	6	9	7
rect	8	7	9	8
rect	8	8	9	9
rect	8	9	9	10
rect	8	10	9	11
rect	8	11	9	12
rect	8	12	9	13
rect	8	13	9	14
rect	8	14	9	15
rect	8	15	9	16
rect	8	16	9	17
rect	8	17	9	18
rect	8	18	9	19
rect	8	19	9	20
rect	8	20	9	21
rect	8	21	9	22
rect	8	22	9	23
rect	8	23	9	24
rect	8	24	9	25
rect	8	25	9	26
rect	8	26	9	27
rect	8	27	9	28
rect	8	28	9	29
rect	8	29	9	30
rect	8	30	9	31
rect	8	31	9	32
rect	8	32	9	33
rect	8	33	9	34
rect	8	34	9	35
rect	8	35	9	36
rect	8	36	9	37
rect	8	37	9	38
rect	8	38	9	39
rect	8	39	9	40
rect	8	40	9	41
rect	8	41	9	42
rect	8	42	9	43
rect	8	43	9	44
rect	8	44	9	45
rect	8	45	9	46
rect	8	46	9	47
rect	8	47	9	48
rect	8	48	9	49
rect	8	49	9	50
rect	8	50	9	51
rect	8	51	9	52
rect	8	52	9	53
rect	8	53	9	54
rect	8	54	9	55
rect	8	55	9	56
rect	8	56	9	57
rect	8	57	9	58
rect	8	58	9	59
rect	8	59	9	60
rect	8	60	9	61
rect	8	61	9	62
rect	8	62	9	63
rect	8	63	9	64
rect	8	64	9	65
rect	8	65	9	66
rect	8	66	9	67
rect	8	67	9	68
rect	8	68	9	69
rect	8	69	9	70
rect	8	70	9	71
rect	8	71	9	72
rect	8	72	9	73
rect	8	73	9	74
rect	8	74	9	75
rect	8	75	9	76
rect	8	76	9	77
rect	8	77	9	78
rect	8	78	9	79
rect	8	79	9	80
rect	8	80	9	81
rect	8	81	9	82
rect	8	82	9	83
rect	8	83	9	84
rect	8	84	9	85
rect	8	85	9	86
rect	8	86	9	87
rect	8	87	9	88
rect	8	88	9	89
rect	8	89	9	90
rect	8	90	9	91
rect	8	91	9	92
rect	8	92	9	93
rect	8	93	9	94
rect	8	94	9	95
rect	8	95	9	96
rect	8	96	9	97
rect	8	97	9	98
rect	8	98	9	99
rect	8	99	9	100
rect	8	100	9	101
rect	8	101	9	102
rect	8	102	9	103
rect	8	103	9	104
rect	8	104	9	105
rect	8	105	9	106
rect	8	106	9	107
rect	8	107	9	108
rect	8	108	9	109
rect	8	109	9	110
rect	8	110	9	111
rect	8	111	9	112
rect	8	112	9	113
rect	8	113	9	114
rect	8	114	9	115
rect	8	115	9	116
rect	8	116	9	117
rect	8	117	9	118
rect	8	118	9	119
rect	8	119	9	120
rect	8	120	9	121
rect	8	121	9	122
rect	8	122	9	123
rect	8	123	9	124
rect	8	124	9	125
rect	8	125	9	126
rect	8	126	9	127
rect	8	127	9	128
rect	8	128	9	129
rect	8	129	9	130
rect	8	130	9	131
rect	8	131	9	132
rect	8	132	9	133
rect	8	133	9	134
rect	8	134	9	135
rect	8	135	9	136
rect	8	136	9	137
rect	8	137	9	138
rect	8	138	9	139
rect	8	139	9	140
rect	8	140	9	141
rect	8	141	9	142
rect	8	142	9	143
rect	8	143	9	144
rect	8	144	9	145
rect	8	145	9	146
rect	8	146	9	147
rect	8	147	9	148
rect	8	148	9	149
rect	8	149	9	150
rect	8	150	9	151
rect	8	151	9	152
rect	8	152	9	153
rect	8	153	9	154
rect	8	154	9	155
rect	8	155	9	156
rect	8	156	9	157
rect	8	157	9	158
rect	8	158	9	159
rect	8	159	9	160
rect	8	160	9	161
rect	8	161	9	162
rect	8	162	9	163
rect	8	163	9	164
rect	8	164	9	165
rect	8	165	9	166
rect	8	166	9	167
rect	8	167	9	168
rect	8	168	9	169
rect	8	169	9	170
rect	8	170	9	171
rect	8	171	9	172
rect	8	172	9	173
rect	8	173	9	174
rect	9	0	10	1
rect	9	1	10	2
rect	9	2	10	3
rect	9	3	10	4
rect	9	4	10	5
rect	9	5	10	6
rect	9	6	10	7
rect	9	7	10	8
rect	9	8	10	9
rect	9	9	10	10
rect	9	10	10	11
rect	9	11	10	12
rect	9	12	10	13
rect	9	13	10	14
rect	9	14	10	15
rect	9	15	10	16
rect	9	16	10	17
rect	9	17	10	18
rect	9	18	10	19
rect	9	19	10	20
rect	9	20	10	21
rect	9	21	10	22
rect	9	22	10	23
rect	9	23	10	24
rect	9	24	10	25
rect	9	25	10	26
rect	9	26	10	27
rect	9	27	10	28
rect	9	28	10	29
rect	9	29	10	30
rect	9	30	10	31
rect	9	31	10	32
rect	9	32	10	33
rect	9	33	10	34
rect	9	34	10	35
rect	9	35	10	36
rect	9	36	10	37
rect	9	37	10	38
rect	9	38	10	39
rect	9	39	10	40
rect	9	40	10	41
rect	9	41	10	42
rect	9	42	10	43
rect	9	43	10	44
rect	9	44	10	45
rect	9	45	10	46
rect	9	46	10	47
rect	9	47	10	48
rect	9	48	10	49
rect	9	49	10	50
rect	9	50	10	51
rect	9	51	10	52
rect	9	52	10	53
rect	9	53	10	54
rect	9	54	10	55
rect	9	55	10	56
rect	9	56	10	57
rect	9	57	10	58
rect	9	58	10	59
rect	9	59	10	60
rect	9	60	10	61
rect	9	61	10	62
rect	9	62	10	63
rect	9	63	10	64
rect	9	64	10	65
rect	9	65	10	66
rect	9	66	10	67
rect	9	67	10	68
rect	9	68	10	69
rect	9	69	10	70
rect	9	70	10	71
rect	9	71	10	72
rect	9	72	10	73
rect	9	73	10	74
rect	9	74	10	75
rect	9	75	10	76
rect	9	76	10	77
rect	9	77	10	78
rect	9	78	10	79
rect	9	79	10	80
rect	9	80	10	81
rect	9	81	10	82
rect	9	82	10	83
rect	9	83	10	84
rect	9	84	10	85
rect	9	85	10	86
rect	9	86	10	87
rect	9	87	10	88
rect	9	88	10	89
rect	9	89	10	90
rect	9	90	10	91
rect	9	91	10	92
rect	9	92	10	93
rect	9	93	10	94
rect	9	94	10	95
rect	9	95	10	96
rect	9	96	10	97
rect	9	97	10	98
rect	9	98	10	99
rect	9	99	10	100
rect	9	100	10	101
rect	9	101	10	102
rect	9	102	10	103
rect	9	103	10	104
rect	9	104	10	105
rect	9	105	10	106
rect	9	106	10	107
rect	9	107	10	108
rect	9	108	10	109
rect	9	109	10	110
rect	9	110	10	111
rect	9	111	10	112
rect	9	112	10	113
rect	9	113	10	114
rect	9	114	10	115
rect	9	115	10	116
rect	9	116	10	117
rect	9	117	10	118
rect	9	118	10	119
rect	9	119	10	120
rect	9	120	10	121
rect	9	121	10	122
rect	9	122	10	123
rect	9	123	10	124
rect	9	124	10	125
rect	9	125	10	126
rect	9	126	10	127
rect	9	127	10	128
rect	9	128	10	129
rect	9	129	10	130
rect	9	130	10	131
rect	9	131	10	132
rect	9	132	10	133
rect	9	133	10	134
rect	9	134	10	135
rect	9	135	10	136
rect	9	136	10	137
rect	9	137	10	138
rect	9	138	10	139
rect	9	139	10	140
rect	9	140	10	141
rect	9	141	10	142
rect	9	142	10	143
rect	9	143	10	144
rect	9	144	10	145
rect	9	145	10	146
rect	9	146	10	147
rect	9	147	10	148
rect	9	148	10	149
rect	9	149	10	150
rect	9	150	10	151
rect	9	151	10	152
rect	9	152	10	153
rect	9	153	10	154
rect	9	154	10	155
rect	9	155	10	156
rect	9	156	10	157
rect	9	157	10	158
rect	9	158	10	159
rect	9	159	10	160
rect	9	160	10	161
rect	9	161	10	162
rect	9	162	10	163
rect	9	163	10	164
rect	9	164	10	165
rect	9	165	10	166
rect	9	166	10	167
rect	9	167	10	168
rect	9	168	10	169
rect	9	169	10	170
rect	9	170	10	171
rect	9	171	10	172
rect	9	172	10	173
rect	9	173	10	174
rect	10	0	11	1
rect	10	1	11	2
rect	10	2	11	3
rect	10	3	11	4
rect	10	4	11	5
rect	10	5	11	6
rect	10	6	11	7
rect	10	7	11	8
rect	10	8	11	9
rect	10	9	11	10
rect	10	10	11	11
rect	10	11	11	12
rect	10	12	11	13
rect	10	13	11	14
rect	10	14	11	15
rect	10	15	11	16
rect	10	16	11	17
rect	10	17	11	18
rect	10	18	11	19
rect	10	19	11	20
rect	10	20	11	21
rect	10	21	11	22
rect	10	22	11	23
rect	10	23	11	24
rect	10	24	11	25
rect	10	25	11	26
rect	10	26	11	27
rect	10	27	11	28
rect	10	28	11	29
rect	10	29	11	30
rect	10	30	11	31
rect	10	31	11	32
rect	10	32	11	33
rect	10	33	11	34
rect	10	34	11	35
rect	10	35	11	36
rect	10	36	11	37
rect	10	37	11	38
rect	10	38	11	39
rect	10	39	11	40
rect	10	40	11	41
rect	10	41	11	42
rect	10	42	11	43
rect	10	43	11	44
rect	10	44	11	45
rect	10	45	11	46
rect	10	46	11	47
rect	10	47	11	48
rect	10	48	11	49
rect	10	49	11	50
rect	10	50	11	51
rect	10	51	11	52
rect	10	52	11	53
rect	10	53	11	54
rect	10	54	11	55
rect	10	55	11	56
rect	10	56	11	57
rect	10	57	11	58
rect	10	58	11	59
rect	10	59	11	60
rect	10	60	11	61
rect	10	61	11	62
rect	10	62	11	63
rect	10	63	11	64
rect	10	64	11	65
rect	10	65	11	66
rect	10	66	11	67
rect	10	67	11	68
rect	10	68	11	69
rect	10	69	11	70
rect	10	70	11	71
rect	10	71	11	72
rect	10	72	11	73
rect	10	73	11	74
rect	10	74	11	75
rect	10	75	11	76
rect	10	76	11	77
rect	10	77	11	78
rect	10	78	11	79
rect	10	79	11	80
rect	10	80	11	81
rect	10	81	11	82
rect	10	82	11	83
rect	10	83	11	84
rect	10	84	11	85
rect	10	85	11	86
rect	10	86	11	87
rect	10	87	11	88
rect	10	88	11	89
rect	10	89	11	90
rect	10	90	11	91
rect	10	91	11	92
rect	10	92	11	93
rect	10	93	11	94
rect	10	94	11	95
rect	10	95	11	96
rect	10	96	11	97
rect	10	97	11	98
rect	10	98	11	99
rect	10	99	11	100
rect	10	100	11	101
rect	10	101	11	102
rect	10	102	11	103
rect	10	103	11	104
rect	10	104	11	105
rect	10	105	11	106
rect	10	106	11	107
rect	10	107	11	108
rect	10	108	11	109
rect	10	109	11	110
rect	10	110	11	111
rect	10	111	11	112
rect	10	112	11	113
rect	10	113	11	114
rect	10	114	11	115
rect	10	115	11	116
rect	10	116	11	117
rect	10	117	11	118
rect	10	118	11	119
rect	10	119	11	120
rect	10	120	11	121
rect	10	121	11	122
rect	10	122	11	123
rect	10	123	11	124
rect	10	124	11	125
rect	10	125	11	126
rect	10	126	11	127
rect	10	127	11	128
rect	10	128	11	129
rect	10	129	11	130
rect	10	130	11	131
rect	10	131	11	132
rect	10	132	11	133
rect	10	133	11	134
rect	10	134	11	135
rect	10	135	11	136
rect	10	136	11	137
rect	10	137	11	138
rect	10	138	11	139
rect	10	139	11	140
rect	10	140	11	141
rect	10	141	11	142
rect	10	142	11	143
rect	10	143	11	144
rect	10	144	11	145
rect	10	145	11	146
rect	10	146	11	147
rect	10	147	11	148
rect	10	148	11	149
rect	10	149	11	150
rect	10	150	11	151
rect	10	151	11	152
rect	10	152	11	153
rect	10	153	11	154
rect	10	154	11	155
rect	10	155	11	156
rect	10	156	11	157
rect	10	157	11	158
rect	10	158	11	159
rect	10	159	11	160
rect	10	160	11	161
rect	10	161	11	162
rect	10	162	11	163
rect	10	163	11	164
rect	10	164	11	165
rect	10	165	11	166
rect	10	166	11	167
rect	10	167	11	168
rect	10	168	11	169
rect	10	169	11	170
rect	10	170	11	171
rect	10	171	11	172
rect	10	172	11	173
rect	10	173	11	174
rect	11	0	12	1
rect	11	1	12	2
rect	11	2	12	3
rect	11	3	12	4
rect	11	4	12	5
rect	11	5	12	6
rect	11	6	12	7
rect	11	7	12	8
rect	11	8	12	9
rect	11	9	12	10
rect	11	10	12	11
rect	11	11	12	12
rect	11	12	12	13
rect	11	13	12	14
rect	11	14	12	15
rect	11	15	12	16
rect	11	16	12	17
rect	11	17	12	18
rect	11	18	12	19
rect	11	19	12	20
rect	11	20	12	21
rect	11	21	12	22
rect	11	22	12	23
rect	11	23	12	24
rect	11	24	12	25
rect	11	25	12	26
rect	11	26	12	27
rect	11	27	12	28
rect	11	28	12	29
rect	11	29	12	30
rect	11	30	12	31
rect	11	31	12	32
rect	11	32	12	33
rect	11	33	12	34
rect	11	34	12	35
rect	11	35	12	36
rect	11	36	12	37
rect	11	37	12	38
rect	11	38	12	39
rect	11	39	12	40
rect	11	40	12	41
rect	11	41	12	42
rect	11	42	12	43
rect	11	43	12	44
rect	11	44	12	45
rect	11	45	12	46
rect	11	46	12	47
rect	11	47	12	48
rect	11	48	12	49
rect	11	49	12	50
rect	11	50	12	51
rect	11	51	12	52
rect	11	52	12	53
rect	11	53	12	54
rect	11	54	12	55
rect	11	55	12	56
rect	11	56	12	57
rect	11	57	12	58
rect	11	58	12	59
rect	11	59	12	60
rect	11	60	12	61
rect	11	61	12	62
rect	11	62	12	63
rect	11	63	12	64
rect	11	64	12	65
rect	11	65	12	66
rect	11	66	12	67
rect	11	67	12	68
rect	11	68	12	69
rect	11	69	12	70
rect	11	70	12	71
rect	11	71	12	72
rect	11	72	12	73
rect	11	73	12	74
rect	11	74	12	75
rect	11	75	12	76
rect	11	76	12	77
rect	11	77	12	78
rect	11	78	12	79
rect	11	79	12	80
rect	11	80	12	81
rect	11	81	12	82
rect	11	82	12	83
rect	11	83	12	84
rect	11	84	12	85
rect	11	85	12	86
rect	11	86	12	87
rect	11	87	12	88
rect	11	88	12	89
rect	11	89	12	90
rect	11	90	12	91
rect	11	91	12	92
rect	11	92	12	93
rect	11	93	12	94
rect	11	94	12	95
rect	11	95	12	96
rect	11	96	12	97
rect	11	97	12	98
rect	11	98	12	99
rect	11	99	12	100
rect	11	100	12	101
rect	11	101	12	102
rect	11	102	12	103
rect	11	103	12	104
rect	11	104	12	105
rect	11	105	12	106
rect	11	106	12	107
rect	11	107	12	108
rect	11	108	12	109
rect	11	109	12	110
rect	11	110	12	111
rect	11	111	12	112
rect	11	112	12	113
rect	11	113	12	114
rect	11	114	12	115
rect	11	115	12	116
rect	11	116	12	117
rect	11	117	12	118
rect	11	118	12	119
rect	11	119	12	120
rect	11	120	12	121
rect	11	121	12	122
rect	11	122	12	123
rect	11	123	12	124
rect	11	124	12	125
rect	11	125	12	126
rect	11	126	12	127
rect	11	127	12	128
rect	11	128	12	129
rect	11	129	12	130
rect	11	130	12	131
rect	11	131	12	132
rect	11	132	12	133
rect	11	133	12	134
rect	11	134	12	135
rect	11	135	12	136
rect	11	136	12	137
rect	11	137	12	138
rect	11	138	12	139
rect	11	139	12	140
rect	11	140	12	141
rect	11	141	12	142
rect	11	142	12	143
rect	11	143	12	144
rect	11	144	12	145
rect	11	145	12	146
rect	11	146	12	147
rect	11	147	12	148
rect	11	148	12	149
rect	11	149	12	150
rect	11	150	12	151
rect	11	151	12	152
rect	11	152	12	153
rect	11	153	12	154
rect	11	154	12	155
rect	11	155	12	156
rect	11	156	12	157
rect	11	157	12	158
rect	11	158	12	159
rect	11	159	12	160
rect	11	160	12	161
rect	11	161	12	162
rect	11	162	12	163
rect	11	163	12	164
rect	11	164	12	165
rect	11	165	12	166
rect	11	166	12	167
rect	11	167	12	168
rect	11	168	12	169
rect	11	169	12	170
rect	11	170	12	171
rect	11	171	12	172
rect	11	172	12	173
rect	11	173	12	174
rect	27	68	28	69
rect	27	69	28	70
rect	27	70	28	71
rect	27	71	28	72
rect	27	72	28	73
rect	27	73	28	74
rect	27	74	28	75
rect	27	75	28	76
rect	27	77	28	78
rect	27	78	28	79
rect	29	0	30	1
rect	29	1	30	2
rect	29	2	30	3
rect	29	3	30	4
rect	29	4	30	5
rect	29	5	30	6
rect	29	6	30	7
rect	29	7	30	8
rect	29	8	30	9
rect	29	9	30	10
rect	29	10	30	11
rect	29	11	30	12
rect	29	12	30	13
rect	29	13	30	14
rect	29	14	30	15
rect	29	15	30	16
rect	29	16	30	17
rect	29	17	30	18
rect	29	18	30	19
rect	29	19	30	20
rect	29	20	30	21
rect	29	21	30	22
rect	29	22	30	23
rect	29	23	30	24
rect	29	24	30	25
rect	29	25	30	26
rect	29	26	30	27
rect	29	27	30	28
rect	29	28	30	29
rect	29	29	30	30
rect	29	30	30	31
rect	29	31	30	32
rect	29	32	30	33
rect	29	33	30	34
rect	29	34	30	35
rect	29	35	30	36
rect	29	36	30	37
rect	29	37	30	38
rect	29	38	30	39
rect	29	39	30	40
rect	29	40	30	41
rect	29	41	30	42
rect	29	42	30	43
rect	29	43	30	44
rect	29	44	30	45
rect	29	45	30	46
rect	29	46	30	47
rect	29	47	30	48
rect	29	48	30	49
rect	29	49	30	50
rect	29	50	30	51
rect	29	51	30	52
rect	29	52	30	53
rect	29	53	30	54
rect	29	54	30	55
rect	29	55	30	56
rect	29	56	30	57
rect	29	57	30	58
rect	29	58	30	59
rect	29	59	30	60
rect	29	60	30	61
rect	29	61	30	62
rect	29	62	30	63
rect	29	63	30	64
rect	29	64	30	65
rect	29	65	30	66
rect	29	66	30	67
rect	29	67	30	68
rect	29	68	30	69
rect	29	69	30	70
rect	29	70	30	71
rect	29	71	30	72
rect	29	72	30	73
rect	29	73	30	74
rect	29	74	30	75
rect	29	75	30	76
rect	29	76	30	77
rect	29	77	30	78
rect	29	78	30	79
rect	29	79	30	80
rect	29	80	30	81
rect	29	81	30	82
rect	29	82	30	83
rect	29	83	30	84
rect	29	84	30	85
rect	29	85	30	86
rect	29	86	30	87
rect	29	87	30	88
rect	29	88	30	89
rect	29	89	30	90
rect	29	90	30	91
rect	29	91	30	92
rect	29	92	30	93
rect	29	93	30	94
rect	29	94	30	95
rect	29	95	30	96
rect	29	96	30	97
rect	29	97	30	98
rect	29	98	30	99
rect	29	99	30	100
rect	29	100	30	101
rect	29	101	30	102
rect	29	102	30	103
rect	29	103	30	104
rect	29	104	30	105
rect	29	105	30	106
rect	29	106	30	107
rect	29	107	30	108
rect	29	108	30	109
rect	29	109	30	110
rect	29	110	30	111
rect	29	111	30	112
rect	29	112	30	113
rect	29	113	30	114
rect	29	114	30	115
rect	29	115	30	116
rect	29	116	30	117
rect	29	117	30	118
rect	29	118	30	119
rect	29	119	30	120
rect	29	120	30	121
rect	29	121	30	122
rect	29	122	30	123
rect	29	123	30	124
rect	29	124	30	125
rect	29	125	30	126
rect	29	126	30	127
rect	29	127	30	128
rect	29	128	30	129
rect	29	129	30	130
rect	29	130	30	131
rect	29	131	30	132
rect	29	132	30	133
rect	29	133	30	134
rect	29	134	30	135
rect	29	135	30	136
rect	29	136	30	137
rect	29	137	30	138
rect	29	138	30	139
rect	29	139	30	140
rect	29	140	30	141
rect	29	141	30	142
rect	29	142	30	143
rect	29	143	30	144
rect	29	144	30	145
rect	29	145	30	146
rect	29	146	30	147
rect	29	147	30	148
rect	29	148	30	149
rect	29	149	30	150
rect	29	150	30	151
rect	29	151	30	152
rect	29	152	30	153
rect	29	153	30	154
rect	29	154	30	155
rect	29	155	30	156
rect	29	156	30	157
rect	29	157	30	158
rect	29	158	30	159
rect	29	159	30	160
rect	29	160	30	161
rect	29	161	30	162
rect	29	162	30	163
rect	29	163	30	164
rect	29	164	30	165
rect	29	165	30	166
rect	29	166	30	167
rect	29	167	30	168
rect	29	168	30	169
rect	29	169	30	170
rect	29	170	30	171
rect	29	171	30	172
rect	29	172	30	173
rect	29	173	30	174
rect	29	174	30	175
rect	29	175	30	176
rect	29	176	30	177
rect	29	177	30	178
rect	29	178	30	179
rect	29	179	30	180
rect	29	180	30	181
rect	29	181	30	182
rect	29	182	30	183
rect	29	183	30	184
rect	29	184	30	185
rect	29	185	30	186
rect	29	186	30	187
rect	29	187	30	188
rect	29	188	30	189
rect	29	189	30	190
rect	29	190	30	191
rect	29	191	30	192
rect	29	192	30	193
rect	29	193	30	194
rect	29	194	30	195
rect	29	195	30	196
rect	29	196	30	197
rect	29	197	30	198
rect	29	198	30	199
rect	29	199	30	200
rect	29	200	30	201
rect	29	201	30	202
rect	29	202	30	203
rect	29	203	30	204
rect	29	204	30	205
rect	29	205	30	206
rect	29	206	30	207
rect	29	207	30	208
rect	29	208	30	209
rect	29	209	30	210
rect	29	210	30	211
rect	29	211	30	212
rect	29	212	30	213
rect	29	213	30	214
rect	29	214	30	215
rect	29	215	30	216
rect	30	0	31	1
rect	30	1	31	2
rect	30	2	31	3
rect	30	3	31	4
rect	30	4	31	5
rect	30	5	31	6
rect	30	6	31	7
rect	30	7	31	8
rect	30	8	31	9
rect	30	9	31	10
rect	30	10	31	11
rect	30	11	31	12
rect	30	12	31	13
rect	30	13	31	14
rect	30	14	31	15
rect	30	15	31	16
rect	30	16	31	17
rect	30	17	31	18
rect	30	18	31	19
rect	30	19	31	20
rect	30	20	31	21
rect	30	21	31	22
rect	30	22	31	23
rect	30	23	31	24
rect	30	24	31	25
rect	30	25	31	26
rect	30	26	31	27
rect	30	27	31	28
rect	30	28	31	29
rect	30	29	31	30
rect	30	30	31	31
rect	30	31	31	32
rect	30	32	31	33
rect	30	33	31	34
rect	30	34	31	35
rect	30	35	31	36
rect	30	36	31	37
rect	30	37	31	38
rect	30	38	31	39
rect	30	39	31	40
rect	30	40	31	41
rect	30	41	31	42
rect	30	42	31	43
rect	30	43	31	44
rect	30	44	31	45
rect	30	45	31	46
rect	30	46	31	47
rect	30	47	31	48
rect	30	48	31	49
rect	30	49	31	50
rect	30	50	31	51
rect	30	51	31	52
rect	30	52	31	53
rect	30	53	31	54
rect	30	54	31	55
rect	30	55	31	56
rect	30	56	31	57
rect	30	57	31	58
rect	30	58	31	59
rect	30	59	31	60
rect	30	60	31	61
rect	30	61	31	62
rect	30	62	31	63
rect	30	63	31	64
rect	30	64	31	65
rect	30	65	31	66
rect	30	66	31	67
rect	30	67	31	68
rect	30	68	31	69
rect	30	69	31	70
rect	30	70	31	71
rect	30	71	31	72
rect	30	72	31	73
rect	30	73	31	74
rect	30	74	31	75
rect	30	75	31	76
rect	30	76	31	77
rect	30	77	31	78
rect	30	78	31	79
rect	30	79	31	80
rect	30	80	31	81
rect	30	81	31	82
rect	30	82	31	83
rect	30	83	31	84
rect	30	84	31	85
rect	30	85	31	86
rect	30	86	31	87
rect	30	87	31	88
rect	30	88	31	89
rect	30	89	31	90
rect	30	90	31	91
rect	30	91	31	92
rect	30	92	31	93
rect	30	93	31	94
rect	30	94	31	95
rect	30	95	31	96
rect	30	96	31	97
rect	30	97	31	98
rect	30	98	31	99
rect	30	99	31	100
rect	30	100	31	101
rect	30	101	31	102
rect	30	102	31	103
rect	30	103	31	104
rect	30	104	31	105
rect	30	105	31	106
rect	30	106	31	107
rect	30	107	31	108
rect	30	108	31	109
rect	30	109	31	110
rect	30	110	31	111
rect	30	111	31	112
rect	30	112	31	113
rect	30	113	31	114
rect	30	114	31	115
rect	30	115	31	116
rect	30	116	31	117
rect	30	117	31	118
rect	30	118	31	119
rect	30	119	31	120
rect	30	120	31	121
rect	30	121	31	122
rect	30	122	31	123
rect	30	123	31	124
rect	30	124	31	125
rect	30	125	31	126
rect	30	126	31	127
rect	30	127	31	128
rect	30	128	31	129
rect	30	129	31	130
rect	30	130	31	131
rect	30	131	31	132
rect	30	132	31	133
rect	30	133	31	134
rect	30	134	31	135
rect	30	135	31	136
rect	30	136	31	137
rect	30	137	31	138
rect	30	138	31	139
rect	30	139	31	140
rect	30	140	31	141
rect	30	141	31	142
rect	30	142	31	143
rect	30	143	31	144
rect	30	144	31	145
rect	30	145	31	146
rect	30	146	31	147
rect	30	147	31	148
rect	30	148	31	149
rect	30	149	31	150
rect	30	150	31	151
rect	30	151	31	152
rect	30	152	31	153
rect	30	153	31	154
rect	30	154	31	155
rect	30	155	31	156
rect	30	156	31	157
rect	30	157	31	158
rect	30	158	31	159
rect	30	159	31	160
rect	30	160	31	161
rect	30	161	31	162
rect	30	162	31	163
rect	30	163	31	164
rect	30	164	31	165
rect	30	165	31	166
rect	30	166	31	167
rect	30	167	31	168
rect	30	168	31	169
rect	30	169	31	170
rect	30	170	31	171
rect	30	171	31	172
rect	30	172	31	173
rect	30	173	31	174
rect	30	174	31	175
rect	30	175	31	176
rect	30	176	31	177
rect	30	177	31	178
rect	30	178	31	179
rect	30	179	31	180
rect	30	180	31	181
rect	30	181	31	182
rect	30	182	31	183
rect	30	183	31	184
rect	30	184	31	185
rect	30	185	31	186
rect	30	186	31	187
rect	30	187	31	188
rect	30	188	31	189
rect	30	189	31	190
rect	30	190	31	191
rect	30	191	31	192
rect	30	192	31	193
rect	30	193	31	194
rect	30	194	31	195
rect	30	195	31	196
rect	30	196	31	197
rect	30	197	31	198
rect	30	198	31	199
rect	30	199	31	200
rect	30	200	31	201
rect	30	201	31	202
rect	30	202	31	203
rect	30	203	31	204
rect	30	204	31	205
rect	30	205	31	206
rect	30	206	31	207
rect	30	207	31	208
rect	30	208	31	209
rect	30	209	31	210
rect	30	210	31	211
rect	30	211	31	212
rect	30	212	31	213
rect	30	213	31	214
rect	30	214	31	215
rect	30	215	31	216
rect	31	0	32	1
rect	31	1	32	2
rect	31	2	32	3
rect	31	3	32	4
rect	31	4	32	5
rect	31	5	32	6
rect	31	6	32	7
rect	31	7	32	8
rect	31	8	32	9
rect	31	9	32	10
rect	31	10	32	11
rect	31	11	32	12
rect	31	12	32	13
rect	31	13	32	14
rect	31	14	32	15
rect	31	15	32	16
rect	31	16	32	17
rect	31	17	32	18
rect	31	18	32	19
rect	31	19	32	20
rect	31	20	32	21
rect	31	21	32	22
rect	31	22	32	23
rect	31	23	32	24
rect	31	24	32	25
rect	31	25	32	26
rect	31	26	32	27
rect	31	27	32	28
rect	31	28	32	29
rect	31	29	32	30
rect	31	30	32	31
rect	31	31	32	32
rect	31	32	32	33
rect	31	33	32	34
rect	31	34	32	35
rect	31	35	32	36
rect	31	36	32	37
rect	31	37	32	38
rect	31	38	32	39
rect	31	39	32	40
rect	31	40	32	41
rect	31	41	32	42
rect	31	42	32	43
rect	31	43	32	44
rect	31	44	32	45
rect	31	45	32	46
rect	31	46	32	47
rect	31	47	32	48
rect	31	48	32	49
rect	31	49	32	50
rect	31	50	32	51
rect	31	51	32	52
rect	31	52	32	53
rect	31	53	32	54
rect	31	54	32	55
rect	31	55	32	56
rect	31	56	32	57
rect	31	57	32	58
rect	31	58	32	59
rect	31	59	32	60
rect	31	60	32	61
rect	31	61	32	62
rect	31	62	32	63
rect	31	63	32	64
rect	31	64	32	65
rect	31	65	32	66
rect	31	66	32	67
rect	31	67	32	68
rect	31	68	32	69
rect	31	69	32	70
rect	31	70	32	71
rect	31	71	32	72
rect	31	72	32	73
rect	31	73	32	74
rect	31	74	32	75
rect	31	75	32	76
rect	31	76	32	77
rect	31	77	32	78
rect	31	78	32	79
rect	31	79	32	80
rect	31	80	32	81
rect	31	81	32	82
rect	31	82	32	83
rect	31	83	32	84
rect	31	84	32	85
rect	31	85	32	86
rect	31	86	32	87
rect	31	87	32	88
rect	31	88	32	89
rect	31	89	32	90
rect	31	90	32	91
rect	31	91	32	92
rect	31	92	32	93
rect	31	93	32	94
rect	31	94	32	95
rect	31	95	32	96
rect	31	96	32	97
rect	31	97	32	98
rect	31	98	32	99
rect	31	99	32	100
rect	31	100	32	101
rect	31	101	32	102
rect	31	102	32	103
rect	31	103	32	104
rect	31	104	32	105
rect	31	105	32	106
rect	31	106	32	107
rect	31	107	32	108
rect	31	108	32	109
rect	31	109	32	110
rect	31	110	32	111
rect	31	111	32	112
rect	31	112	32	113
rect	31	113	32	114
rect	31	114	32	115
rect	31	115	32	116
rect	31	116	32	117
rect	31	117	32	118
rect	31	118	32	119
rect	31	119	32	120
rect	31	120	32	121
rect	31	121	32	122
rect	31	122	32	123
rect	31	123	32	124
rect	31	124	32	125
rect	31	125	32	126
rect	31	126	32	127
rect	31	127	32	128
rect	31	128	32	129
rect	31	129	32	130
rect	31	130	32	131
rect	31	131	32	132
rect	31	132	32	133
rect	31	133	32	134
rect	31	134	32	135
rect	31	135	32	136
rect	31	136	32	137
rect	31	137	32	138
rect	31	138	32	139
rect	31	139	32	140
rect	31	140	32	141
rect	31	141	32	142
rect	31	142	32	143
rect	31	143	32	144
rect	31	144	32	145
rect	31	145	32	146
rect	31	146	32	147
rect	31	147	32	148
rect	31	148	32	149
rect	31	149	32	150
rect	31	150	32	151
rect	31	151	32	152
rect	31	152	32	153
rect	31	153	32	154
rect	31	154	32	155
rect	31	155	32	156
rect	31	156	32	157
rect	31	157	32	158
rect	31	158	32	159
rect	31	159	32	160
rect	31	160	32	161
rect	31	161	32	162
rect	31	162	32	163
rect	31	163	32	164
rect	31	164	32	165
rect	31	165	32	166
rect	31	166	32	167
rect	31	167	32	168
rect	31	168	32	169
rect	31	169	32	170
rect	31	170	32	171
rect	31	171	32	172
rect	31	172	32	173
rect	31	173	32	174
rect	31	174	32	175
rect	31	175	32	176
rect	31	176	32	177
rect	31	177	32	178
rect	31	178	32	179
rect	31	179	32	180
rect	31	180	32	181
rect	31	181	32	182
rect	31	182	32	183
rect	31	183	32	184
rect	31	184	32	185
rect	31	185	32	186
rect	31	186	32	187
rect	31	187	32	188
rect	31	188	32	189
rect	31	189	32	190
rect	31	190	32	191
rect	31	191	32	192
rect	31	192	32	193
rect	31	193	32	194
rect	31	194	32	195
rect	31	195	32	196
rect	31	196	32	197
rect	31	197	32	198
rect	31	198	32	199
rect	31	199	32	200
rect	31	200	32	201
rect	31	201	32	202
rect	31	202	32	203
rect	31	203	32	204
rect	31	204	32	205
rect	31	205	32	206
rect	31	206	32	207
rect	31	207	32	208
rect	31	208	32	209
rect	31	209	32	210
rect	31	210	32	211
rect	31	211	32	212
rect	31	212	32	213
rect	31	213	32	214
rect	31	214	32	215
rect	31	215	32	216
rect	32	0	33	1
rect	32	1	33	2
rect	32	2	33	3
rect	32	3	33	4
rect	32	4	33	5
rect	32	5	33	6
rect	32	6	33	7
rect	32	7	33	8
rect	32	8	33	9
rect	32	9	33	10
rect	32	10	33	11
rect	32	11	33	12
rect	32	12	33	13
rect	32	13	33	14
rect	32	14	33	15
rect	32	15	33	16
rect	32	16	33	17
rect	32	17	33	18
rect	32	18	33	19
rect	32	19	33	20
rect	32	20	33	21
rect	32	21	33	22
rect	32	22	33	23
rect	32	23	33	24
rect	32	24	33	25
rect	32	25	33	26
rect	32	26	33	27
rect	32	27	33	28
rect	32	28	33	29
rect	32	29	33	30
rect	32	30	33	31
rect	32	31	33	32
rect	32	32	33	33
rect	32	33	33	34
rect	32	34	33	35
rect	32	35	33	36
rect	32	36	33	37
rect	32	37	33	38
rect	32	38	33	39
rect	32	39	33	40
rect	32	40	33	41
rect	32	41	33	42
rect	32	42	33	43
rect	32	43	33	44
rect	32	44	33	45
rect	32	45	33	46
rect	32	46	33	47
rect	32	47	33	48
rect	32	48	33	49
rect	32	49	33	50
rect	32	50	33	51
rect	32	51	33	52
rect	32	52	33	53
rect	32	53	33	54
rect	32	54	33	55
rect	32	55	33	56
rect	32	56	33	57
rect	32	57	33	58
rect	32	58	33	59
rect	32	59	33	60
rect	32	60	33	61
rect	32	61	33	62
rect	32	62	33	63
rect	32	63	33	64
rect	32	64	33	65
rect	32	65	33	66
rect	32	66	33	67
rect	32	67	33	68
rect	32	68	33	69
rect	32	69	33	70
rect	32	70	33	71
rect	32	71	33	72
rect	32	72	33	73
rect	32	73	33	74
rect	32	74	33	75
rect	32	75	33	76
rect	32	76	33	77
rect	32	77	33	78
rect	32	78	33	79
rect	32	79	33	80
rect	32	80	33	81
rect	32	81	33	82
rect	32	82	33	83
rect	32	83	33	84
rect	32	84	33	85
rect	32	85	33	86
rect	32	86	33	87
rect	32	87	33	88
rect	32	88	33	89
rect	32	89	33	90
rect	32	90	33	91
rect	32	91	33	92
rect	32	92	33	93
rect	32	93	33	94
rect	32	94	33	95
rect	32	95	33	96
rect	32	96	33	97
rect	32	97	33	98
rect	32	98	33	99
rect	32	99	33	100
rect	32	100	33	101
rect	32	101	33	102
rect	32	102	33	103
rect	32	103	33	104
rect	32	104	33	105
rect	32	105	33	106
rect	32	106	33	107
rect	32	107	33	108
rect	32	108	33	109
rect	32	109	33	110
rect	32	110	33	111
rect	32	111	33	112
rect	32	112	33	113
rect	32	113	33	114
rect	32	114	33	115
rect	32	115	33	116
rect	32	116	33	117
rect	32	117	33	118
rect	32	118	33	119
rect	32	119	33	120
rect	32	120	33	121
rect	32	121	33	122
rect	32	122	33	123
rect	32	123	33	124
rect	32	124	33	125
rect	32	125	33	126
rect	32	126	33	127
rect	32	127	33	128
rect	32	128	33	129
rect	32	129	33	130
rect	32	130	33	131
rect	32	131	33	132
rect	32	132	33	133
rect	32	133	33	134
rect	32	134	33	135
rect	32	135	33	136
rect	32	136	33	137
rect	32	137	33	138
rect	32	138	33	139
rect	32	139	33	140
rect	32	140	33	141
rect	32	141	33	142
rect	32	142	33	143
rect	32	143	33	144
rect	32	144	33	145
rect	32	145	33	146
rect	32	146	33	147
rect	32	147	33	148
rect	32	148	33	149
rect	32	149	33	150
rect	32	150	33	151
rect	32	151	33	152
rect	32	152	33	153
rect	32	153	33	154
rect	32	154	33	155
rect	32	155	33	156
rect	32	156	33	157
rect	32	157	33	158
rect	32	158	33	159
rect	32	159	33	160
rect	32	160	33	161
rect	32	161	33	162
rect	32	162	33	163
rect	32	163	33	164
rect	32	164	33	165
rect	32	165	33	166
rect	32	166	33	167
rect	32	167	33	168
rect	32	168	33	169
rect	32	169	33	170
rect	32	170	33	171
rect	32	171	33	172
rect	32	172	33	173
rect	32	173	33	174
rect	32	174	33	175
rect	32	175	33	176
rect	32	176	33	177
rect	32	177	33	178
rect	32	178	33	179
rect	32	179	33	180
rect	32	180	33	181
rect	32	181	33	182
rect	32	182	33	183
rect	32	183	33	184
rect	32	184	33	185
rect	32	185	33	186
rect	32	186	33	187
rect	32	187	33	188
rect	32	188	33	189
rect	32	189	33	190
rect	32	190	33	191
rect	32	191	33	192
rect	32	192	33	193
rect	32	193	33	194
rect	32	194	33	195
rect	32	195	33	196
rect	32	196	33	197
rect	32	197	33	198
rect	32	198	33	199
rect	32	199	33	200
rect	32	200	33	201
rect	32	201	33	202
rect	32	202	33	203
rect	32	203	33	204
rect	32	204	33	205
rect	32	205	33	206
rect	32	206	33	207
rect	32	207	33	208
rect	32	208	33	209
rect	32	209	33	210
rect	32	210	33	211
rect	32	211	33	212
rect	32	212	33	213
rect	32	213	33	214
rect	32	214	33	215
rect	32	215	33	216
rect	33	0	34	1
rect	33	1	34	2
rect	33	2	34	3
rect	33	3	34	4
rect	33	4	34	5
rect	33	5	34	6
rect	33	6	34	7
rect	33	7	34	8
rect	33	8	34	9
rect	33	9	34	10
rect	33	10	34	11
rect	33	11	34	12
rect	33	12	34	13
rect	33	13	34	14
rect	33	14	34	15
rect	33	15	34	16
rect	33	16	34	17
rect	33	17	34	18
rect	33	18	34	19
rect	33	19	34	20
rect	33	20	34	21
rect	33	21	34	22
rect	33	22	34	23
rect	33	23	34	24
rect	33	24	34	25
rect	33	25	34	26
rect	33	26	34	27
rect	33	27	34	28
rect	33	28	34	29
rect	33	29	34	30
rect	33	30	34	31
rect	33	31	34	32
rect	33	32	34	33
rect	33	33	34	34
rect	33	34	34	35
rect	33	35	34	36
rect	33	36	34	37
rect	33	37	34	38
rect	33	38	34	39
rect	33	39	34	40
rect	33	40	34	41
rect	33	41	34	42
rect	33	42	34	43
rect	33	43	34	44
rect	33	44	34	45
rect	33	45	34	46
rect	33	46	34	47
rect	33	47	34	48
rect	33	48	34	49
rect	33	49	34	50
rect	33	50	34	51
rect	33	51	34	52
rect	33	52	34	53
rect	33	53	34	54
rect	33	54	34	55
rect	33	55	34	56
rect	33	56	34	57
rect	33	57	34	58
rect	33	58	34	59
rect	33	59	34	60
rect	33	60	34	61
rect	33	61	34	62
rect	33	62	34	63
rect	33	63	34	64
rect	33	64	34	65
rect	33	65	34	66
rect	33	66	34	67
rect	33	67	34	68
rect	33	68	34	69
rect	33	69	34	70
rect	33	70	34	71
rect	33	71	34	72
rect	33	72	34	73
rect	33	73	34	74
rect	33	74	34	75
rect	33	75	34	76
rect	33	76	34	77
rect	33	77	34	78
rect	33	78	34	79
rect	33	79	34	80
rect	33	80	34	81
rect	33	81	34	82
rect	33	82	34	83
rect	33	83	34	84
rect	33	84	34	85
rect	33	85	34	86
rect	33	86	34	87
rect	33	87	34	88
rect	33	88	34	89
rect	33	89	34	90
rect	33	90	34	91
rect	33	91	34	92
rect	33	92	34	93
rect	33	93	34	94
rect	33	94	34	95
rect	33	95	34	96
rect	33	96	34	97
rect	33	97	34	98
rect	33	98	34	99
rect	33	99	34	100
rect	33	100	34	101
rect	33	101	34	102
rect	33	102	34	103
rect	33	103	34	104
rect	33	104	34	105
rect	33	105	34	106
rect	33	106	34	107
rect	33	107	34	108
rect	33	108	34	109
rect	33	109	34	110
rect	33	110	34	111
rect	33	111	34	112
rect	33	112	34	113
rect	33	113	34	114
rect	33	114	34	115
rect	33	115	34	116
rect	33	116	34	117
rect	33	117	34	118
rect	33	118	34	119
rect	33	119	34	120
rect	33	120	34	121
rect	33	121	34	122
rect	33	122	34	123
rect	33	123	34	124
rect	33	124	34	125
rect	33	125	34	126
rect	33	126	34	127
rect	33	127	34	128
rect	33	128	34	129
rect	33	129	34	130
rect	33	130	34	131
rect	33	131	34	132
rect	33	132	34	133
rect	33	133	34	134
rect	33	134	34	135
rect	33	135	34	136
rect	33	136	34	137
rect	33	137	34	138
rect	33	138	34	139
rect	33	139	34	140
rect	33	140	34	141
rect	33	141	34	142
rect	33	142	34	143
rect	33	143	34	144
rect	33	144	34	145
rect	33	145	34	146
rect	33	146	34	147
rect	33	147	34	148
rect	33	148	34	149
rect	33	149	34	150
rect	33	150	34	151
rect	33	151	34	152
rect	33	152	34	153
rect	33	153	34	154
rect	33	154	34	155
rect	33	155	34	156
rect	33	156	34	157
rect	33	157	34	158
rect	33	158	34	159
rect	33	159	34	160
rect	33	160	34	161
rect	33	161	34	162
rect	33	162	34	163
rect	33	163	34	164
rect	33	164	34	165
rect	33	165	34	166
rect	33	166	34	167
rect	33	167	34	168
rect	33	168	34	169
rect	33	169	34	170
rect	33	170	34	171
rect	33	171	34	172
rect	33	172	34	173
rect	33	173	34	174
rect	33	174	34	175
rect	33	175	34	176
rect	33	176	34	177
rect	33	177	34	178
rect	33	178	34	179
rect	33	179	34	180
rect	33	180	34	181
rect	33	181	34	182
rect	33	182	34	183
rect	33	183	34	184
rect	33	184	34	185
rect	33	185	34	186
rect	33	186	34	187
rect	33	187	34	188
rect	33	188	34	189
rect	33	189	34	190
rect	33	190	34	191
rect	33	191	34	192
rect	33	192	34	193
rect	33	193	34	194
rect	33	194	34	195
rect	33	195	34	196
rect	33	196	34	197
rect	33	197	34	198
rect	33	198	34	199
rect	33	199	34	200
rect	33	200	34	201
rect	33	201	34	202
rect	33	202	34	203
rect	33	203	34	204
rect	33	204	34	205
rect	33	205	34	206
rect	33	206	34	207
rect	33	207	34	208
rect	33	208	34	209
rect	33	209	34	210
rect	33	210	34	211
rect	33	211	34	212
rect	33	212	34	213
rect	33	213	34	214
rect	33	214	34	215
rect	33	215	34	216
rect	34	0	35	1
rect	34	1	35	2
rect	34	2	35	3
rect	34	3	35	4
rect	34	4	35	5
rect	34	5	35	6
rect	34	6	35	7
rect	34	7	35	8
rect	34	8	35	9
rect	34	9	35	10
rect	34	10	35	11
rect	34	11	35	12
rect	34	12	35	13
rect	34	13	35	14
rect	34	14	35	15
rect	34	15	35	16
rect	34	16	35	17
rect	34	17	35	18
rect	34	18	35	19
rect	34	19	35	20
rect	34	20	35	21
rect	34	21	35	22
rect	34	22	35	23
rect	34	23	35	24
rect	34	24	35	25
rect	34	25	35	26
rect	34	26	35	27
rect	34	27	35	28
rect	34	28	35	29
rect	34	29	35	30
rect	34	30	35	31
rect	34	31	35	32
rect	34	32	35	33
rect	34	33	35	34
rect	34	34	35	35
rect	34	35	35	36
rect	34	36	35	37
rect	34	37	35	38
rect	34	38	35	39
rect	34	39	35	40
rect	34	40	35	41
rect	34	41	35	42
rect	34	42	35	43
rect	34	43	35	44
rect	34	44	35	45
rect	34	45	35	46
rect	34	46	35	47
rect	34	47	35	48
rect	34	48	35	49
rect	34	49	35	50
rect	34	50	35	51
rect	34	51	35	52
rect	34	52	35	53
rect	34	53	35	54
rect	34	54	35	55
rect	34	55	35	56
rect	34	56	35	57
rect	34	57	35	58
rect	34	58	35	59
rect	34	59	35	60
rect	34	60	35	61
rect	34	61	35	62
rect	34	62	35	63
rect	34	63	35	64
rect	34	64	35	65
rect	34	65	35	66
rect	34	66	35	67
rect	34	67	35	68
rect	34	68	35	69
rect	34	69	35	70
rect	34	70	35	71
rect	34	71	35	72
rect	34	72	35	73
rect	34	73	35	74
rect	34	74	35	75
rect	34	75	35	76
rect	34	76	35	77
rect	34	77	35	78
rect	34	78	35	79
rect	34	79	35	80
rect	34	80	35	81
rect	34	81	35	82
rect	34	82	35	83
rect	34	83	35	84
rect	34	84	35	85
rect	34	85	35	86
rect	34	86	35	87
rect	34	87	35	88
rect	34	88	35	89
rect	34	89	35	90
rect	34	90	35	91
rect	34	91	35	92
rect	34	92	35	93
rect	34	93	35	94
rect	34	94	35	95
rect	34	95	35	96
rect	34	96	35	97
rect	34	97	35	98
rect	34	98	35	99
rect	34	99	35	100
rect	34	100	35	101
rect	34	101	35	102
rect	34	102	35	103
rect	34	103	35	104
rect	34	104	35	105
rect	34	105	35	106
rect	34	106	35	107
rect	34	107	35	108
rect	34	108	35	109
rect	34	109	35	110
rect	34	110	35	111
rect	34	111	35	112
rect	34	112	35	113
rect	34	113	35	114
rect	34	114	35	115
rect	34	115	35	116
rect	34	116	35	117
rect	34	117	35	118
rect	34	118	35	119
rect	34	119	35	120
rect	34	120	35	121
rect	34	121	35	122
rect	34	122	35	123
rect	34	123	35	124
rect	34	124	35	125
rect	34	125	35	126
rect	34	126	35	127
rect	34	127	35	128
rect	34	128	35	129
rect	34	129	35	130
rect	34	130	35	131
rect	34	131	35	132
rect	34	132	35	133
rect	34	133	35	134
rect	34	134	35	135
rect	34	135	35	136
rect	34	136	35	137
rect	34	137	35	138
rect	34	138	35	139
rect	34	139	35	140
rect	34	140	35	141
rect	34	141	35	142
rect	34	142	35	143
rect	34	143	35	144
rect	34	144	35	145
rect	34	145	35	146
rect	34	146	35	147
rect	34	147	35	148
rect	34	148	35	149
rect	34	149	35	150
rect	34	150	35	151
rect	34	151	35	152
rect	34	152	35	153
rect	34	153	35	154
rect	34	154	35	155
rect	34	155	35	156
rect	34	156	35	157
rect	34	157	35	158
rect	34	158	35	159
rect	34	159	35	160
rect	34	160	35	161
rect	34	161	35	162
rect	34	162	35	163
rect	34	163	35	164
rect	34	164	35	165
rect	34	165	35	166
rect	34	166	35	167
rect	34	167	35	168
rect	34	168	35	169
rect	34	169	35	170
rect	34	170	35	171
rect	34	171	35	172
rect	34	172	35	173
rect	34	173	35	174
rect	34	174	35	175
rect	34	175	35	176
rect	34	176	35	177
rect	34	177	35	178
rect	34	178	35	179
rect	34	179	35	180
rect	34	180	35	181
rect	34	181	35	182
rect	34	182	35	183
rect	34	183	35	184
rect	34	184	35	185
rect	34	185	35	186
rect	34	186	35	187
rect	34	187	35	188
rect	34	188	35	189
rect	34	189	35	190
rect	34	190	35	191
rect	34	191	35	192
rect	34	192	35	193
rect	34	193	35	194
rect	34	194	35	195
rect	34	195	35	196
rect	34	196	35	197
rect	34	197	35	198
rect	34	198	35	199
rect	34	199	35	200
rect	34	200	35	201
rect	34	201	35	202
rect	34	202	35	203
rect	34	203	35	204
rect	34	204	35	205
rect	34	205	35	206
rect	34	206	35	207
rect	34	207	35	208
rect	34	208	35	209
rect	34	209	35	210
rect	34	210	35	211
rect	34	211	35	212
rect	34	212	35	213
rect	34	213	35	214
rect	34	214	35	215
rect	34	215	35	216
rect	52	0	53	1
rect	52	1	53	2
rect	52	2	53	3
rect	52	3	53	4
rect	52	4	53	5
rect	52	5	53	6
rect	52	6	53	7
rect	52	7	53	8
rect	52	8	53	9
rect	52	9	53	10
rect	52	10	53	11
rect	52	11	53	12
rect	52	12	53	13
rect	52	13	53	14
rect	52	14	53	15
rect	52	15	53	16
rect	52	16	53	17
rect	52	17	53	18
rect	52	18	53	19
rect	52	19	53	20
rect	52	20	53	21
rect	52	21	53	22
rect	52	22	53	23
rect	52	23	53	24
rect	52	24	53	25
rect	52	25	53	26
rect	52	26	53	27
rect	52	27	53	28
rect	52	28	53	29
rect	52	29	53	30
rect	52	30	53	31
rect	52	31	53	32
rect	52	32	53	33
rect	52	33	53	34
rect	52	34	53	35
rect	52	35	53	36
rect	52	36	53	37
rect	52	37	53	38
rect	52	38	53	39
rect	52	39	53	40
rect	52	40	53	41
rect	52	41	53	42
rect	52	42	53	43
rect	52	43	53	44
rect	52	44	53	45
rect	52	45	53	46
rect	52	46	53	47
rect	52	47	53	48
rect	52	48	53	49
rect	52	49	53	50
rect	52	50	53	51
rect	52	51	53	52
rect	52	52	53	53
rect	52	53	53	54
rect	52	54	53	55
rect	52	55	53	56
rect	52	56	53	57
rect	52	57	53	58
rect	52	58	53	59
rect	52	59	53	60
rect	52	60	53	61
rect	52	61	53	62
rect	52	62	53	63
rect	52	63	53	64
rect	52	64	53	65
rect	52	65	53	66
rect	52	66	53	67
rect	52	67	53	68
rect	52	68	53	69
rect	52	69	53	70
rect	52	70	53	71
rect	52	71	53	72
rect	52	72	53	73
rect	52	73	53	74
rect	52	74	53	75
rect	52	75	53	76
rect	52	76	53	77
rect	52	77	53	78
rect	52	78	53	79
rect	52	79	53	80
rect	52	80	53	81
rect	52	81	53	82
rect	52	82	53	83
rect	52	83	53	84
rect	52	84	53	85
rect	52	85	53	86
rect	52	86	53	87
rect	52	87	53	88
rect	52	88	53	89
rect	52	89	53	90
rect	52	90	53	91
rect	52	91	53	92
rect	52	92	53	93
rect	52	93	53	94
rect	52	94	53	95
rect	52	95	53	96
rect	52	96	53	97
rect	52	97	53	98
rect	52	98	53	99
rect	52	99	53	100
rect	52	100	53	101
rect	52	101	53	102
rect	52	102	53	103
rect	52	103	53	104
rect	52	104	53	105
rect	52	105	53	106
rect	52	106	53	107
rect	52	107	53	108
rect	52	108	53	109
rect	52	109	53	110
rect	52	110	53	111
rect	52	111	53	112
rect	52	112	53	113
rect	52	113	53	114
rect	52	114	53	115
rect	52	115	53	116
rect	52	116	53	117
rect	52	117	53	118
rect	52	118	53	119
rect	52	119	53	120
rect	52	120	53	121
rect	52	121	53	122
rect	52	122	53	123
rect	52	123	53	124
rect	52	124	53	125
rect	52	125	53	126
rect	52	126	53	127
rect	52	127	53	128
rect	52	128	53	129
rect	52	129	53	130
rect	52	130	53	131
rect	52	131	53	132
rect	52	132	53	133
rect	52	133	53	134
rect	52	134	53	135
rect	52	135	53	136
rect	52	136	53	137
rect	52	137	53	138
rect	52	138	53	139
rect	52	139	53	140
rect	52	140	53	141
rect	52	141	53	142
rect	52	142	53	143
rect	52	143	53	144
rect	52	144	53	145
rect	52	145	53	146
rect	52	146	53	147
rect	52	147	53	148
rect	52	148	53	149
rect	52	149	53	150
rect	52	150	53	151
rect	52	151	53	152
rect	52	152	53	153
rect	52	153	53	154
rect	52	154	53	155
rect	52	155	53	156
rect	52	156	53	157
rect	52	157	53	158
rect	52	158	53	159
rect	52	159	53	160
rect	52	160	53	161
rect	52	161	53	162
rect	52	162	53	163
rect	52	163	53	164
rect	52	164	53	165
rect	52	165	53	166
rect	52	166	53	167
rect	52	167	53	168
rect	52	168	53	169
rect	52	169	53	170
rect	52	170	53	171
rect	52	171	53	172
rect	52	172	53	173
rect	52	173	53	174
rect	52	174	53	175
rect	52	175	53	176
rect	52	176	53	177
rect	52	177	53	178
rect	52	178	53	179
rect	52	179	53	180
rect	52	180	53	181
rect	52	181	53	182
rect	52	182	53	183
rect	52	183	53	184
rect	52	184	53	185
rect	52	185	53	186
rect	52	186	53	187
rect	52	187	53	188
rect	52	188	53	189
rect	52	189	53	190
rect	52	190	53	191
rect	52	191	53	192
rect	52	192	53	193
rect	52	193	53	194
rect	52	194	53	195
rect	52	195	53	196
rect	52	196	53	197
rect	52	197	53	198
rect	52	198	53	199
rect	52	199	53	200
rect	52	200	53	201
rect	52	201	53	202
rect	52	202	53	203
rect	52	203	53	204
rect	52	204	53	205
rect	52	205	53	206
rect	52	206	53	207
rect	52	207	53	208
rect	52	208	53	209
rect	52	209	53	210
rect	52	210	53	211
rect	52	211	53	212
rect	52	212	53	213
rect	52	213	53	214
rect	52	214	53	215
rect	52	215	53	216
rect	52	216	53	217
rect	52	217	53	218
rect	52	218	53	219
rect	52	219	53	220
rect	52	220	53	221
rect	52	221	53	222
rect	52	222	53	223
rect	52	223	53	224
rect	52	224	53	225
rect	52	225	53	226
rect	52	226	53	227
rect	52	227	53	228
rect	52	228	53	229
rect	52	229	53	230
rect	52	230	53	231
rect	52	231	53	232
rect	52	232	53	233
rect	52	233	53	234
rect	52	234	53	235
rect	52	235	53	236
rect	52	236	53	237
rect	52	237	53	238
rect	52	238	53	239
rect	52	239	53	240
rect	52	240	53	241
rect	52	241	53	242
rect	52	242	53	243
rect	53	0	54	1
rect	53	1	54	2
rect	53	2	54	3
rect	53	3	54	4
rect	53	4	54	5
rect	53	5	54	6
rect	53	6	54	7
rect	53	7	54	8
rect	53	8	54	9
rect	53	9	54	10
rect	53	10	54	11
rect	53	11	54	12
rect	53	12	54	13
rect	53	13	54	14
rect	53	14	54	15
rect	53	15	54	16
rect	53	16	54	17
rect	53	17	54	18
rect	53	18	54	19
rect	53	19	54	20
rect	53	20	54	21
rect	53	21	54	22
rect	53	22	54	23
rect	53	23	54	24
rect	53	24	54	25
rect	53	25	54	26
rect	53	26	54	27
rect	53	27	54	28
rect	53	28	54	29
rect	53	29	54	30
rect	53	30	54	31
rect	53	31	54	32
rect	53	32	54	33
rect	53	33	54	34
rect	53	34	54	35
rect	53	35	54	36
rect	53	36	54	37
rect	53	37	54	38
rect	53	38	54	39
rect	53	39	54	40
rect	53	40	54	41
rect	53	41	54	42
rect	53	42	54	43
rect	53	43	54	44
rect	53	44	54	45
rect	53	45	54	46
rect	53	46	54	47
rect	53	47	54	48
rect	53	48	54	49
rect	53	49	54	50
rect	53	50	54	51
rect	53	51	54	52
rect	53	52	54	53
rect	53	53	54	54
rect	53	54	54	55
rect	53	55	54	56
rect	53	56	54	57
rect	53	57	54	58
rect	53	58	54	59
rect	53	59	54	60
rect	53	60	54	61
rect	53	61	54	62
rect	53	62	54	63
rect	53	63	54	64
rect	53	64	54	65
rect	53	65	54	66
rect	53	66	54	67
rect	53	67	54	68
rect	53	68	54	69
rect	53	69	54	70
rect	53	70	54	71
rect	53	71	54	72
rect	53	72	54	73
rect	53	73	54	74
rect	53	74	54	75
rect	53	75	54	76
rect	53	76	54	77
rect	53	77	54	78
rect	53	78	54	79
rect	53	79	54	80
rect	53	80	54	81
rect	53	81	54	82
rect	53	82	54	83
rect	53	83	54	84
rect	53	84	54	85
rect	53	85	54	86
rect	53	86	54	87
rect	53	87	54	88
rect	53	88	54	89
rect	53	89	54	90
rect	53	90	54	91
rect	53	91	54	92
rect	53	92	54	93
rect	53	93	54	94
rect	53	94	54	95
rect	53	95	54	96
rect	53	96	54	97
rect	53	97	54	98
rect	53	98	54	99
rect	53	99	54	100
rect	53	100	54	101
rect	53	101	54	102
rect	53	102	54	103
rect	53	103	54	104
rect	53	104	54	105
rect	53	105	54	106
rect	53	106	54	107
rect	53	107	54	108
rect	53	108	54	109
rect	53	109	54	110
rect	53	110	54	111
rect	53	111	54	112
rect	53	112	54	113
rect	53	113	54	114
rect	53	114	54	115
rect	53	115	54	116
rect	53	116	54	117
rect	53	117	54	118
rect	53	118	54	119
rect	53	119	54	120
rect	53	120	54	121
rect	53	121	54	122
rect	53	122	54	123
rect	53	123	54	124
rect	53	124	54	125
rect	53	125	54	126
rect	53	126	54	127
rect	53	127	54	128
rect	53	128	54	129
rect	53	129	54	130
rect	53	130	54	131
rect	53	131	54	132
rect	53	132	54	133
rect	53	133	54	134
rect	53	134	54	135
rect	53	135	54	136
rect	53	136	54	137
rect	53	137	54	138
rect	53	138	54	139
rect	53	139	54	140
rect	53	140	54	141
rect	53	141	54	142
rect	53	142	54	143
rect	53	143	54	144
rect	53	144	54	145
rect	53	145	54	146
rect	53	146	54	147
rect	53	147	54	148
rect	53	148	54	149
rect	53	149	54	150
rect	53	150	54	151
rect	53	151	54	152
rect	53	152	54	153
rect	53	153	54	154
rect	53	154	54	155
rect	53	155	54	156
rect	53	156	54	157
rect	53	157	54	158
rect	53	158	54	159
rect	53	159	54	160
rect	53	160	54	161
rect	53	161	54	162
rect	53	162	54	163
rect	53	163	54	164
rect	53	164	54	165
rect	53	165	54	166
rect	53	166	54	167
rect	53	167	54	168
rect	53	168	54	169
rect	53	169	54	170
rect	53	170	54	171
rect	53	171	54	172
rect	53	172	54	173
rect	53	173	54	174
rect	53	174	54	175
rect	53	175	54	176
rect	53	176	54	177
rect	53	177	54	178
rect	53	178	54	179
rect	53	179	54	180
rect	53	180	54	181
rect	53	181	54	182
rect	53	182	54	183
rect	53	183	54	184
rect	53	184	54	185
rect	53	185	54	186
rect	53	186	54	187
rect	53	187	54	188
rect	53	188	54	189
rect	53	189	54	190
rect	53	190	54	191
rect	53	191	54	192
rect	53	192	54	193
rect	53	193	54	194
rect	53	194	54	195
rect	53	195	54	196
rect	53	196	54	197
rect	53	197	54	198
rect	53	198	54	199
rect	53	199	54	200
rect	53	200	54	201
rect	53	201	54	202
rect	53	202	54	203
rect	53	203	54	204
rect	53	204	54	205
rect	53	205	54	206
rect	53	206	54	207
rect	53	207	54	208
rect	53	208	54	209
rect	53	209	54	210
rect	53	210	54	211
rect	53	211	54	212
rect	53	212	54	213
rect	53	213	54	214
rect	53	214	54	215
rect	53	215	54	216
rect	53	216	54	217
rect	53	217	54	218
rect	53	218	54	219
rect	53	219	54	220
rect	53	220	54	221
rect	53	221	54	222
rect	53	222	54	223
rect	53	223	54	224
rect	53	224	54	225
rect	53	225	54	226
rect	53	226	54	227
rect	53	227	54	228
rect	53	228	54	229
rect	53	229	54	230
rect	53	230	54	231
rect	53	231	54	232
rect	53	232	54	233
rect	53	233	54	234
rect	53	234	54	235
rect	53	235	54	236
rect	53	236	54	237
rect	53	237	54	238
rect	53	238	54	239
rect	53	239	54	240
rect	53	240	54	241
rect	53	241	54	242
rect	53	242	54	243
rect	54	0	55	1
rect	54	1	55	2
rect	54	2	55	3
rect	54	3	55	4
rect	54	4	55	5
rect	54	5	55	6
rect	54	6	55	7
rect	54	7	55	8
rect	54	8	55	9
rect	54	9	55	10
rect	54	10	55	11
rect	54	11	55	12
rect	54	12	55	13
rect	54	13	55	14
rect	54	14	55	15
rect	54	15	55	16
rect	54	16	55	17
rect	54	17	55	18
rect	54	18	55	19
rect	54	19	55	20
rect	54	20	55	21
rect	54	21	55	22
rect	54	22	55	23
rect	54	23	55	24
rect	54	24	55	25
rect	54	25	55	26
rect	54	26	55	27
rect	54	27	55	28
rect	54	28	55	29
rect	54	29	55	30
rect	54	30	55	31
rect	54	31	55	32
rect	54	32	55	33
rect	54	33	55	34
rect	54	34	55	35
rect	54	35	55	36
rect	54	36	55	37
rect	54	37	55	38
rect	54	38	55	39
rect	54	39	55	40
rect	54	40	55	41
rect	54	41	55	42
rect	54	42	55	43
rect	54	43	55	44
rect	54	44	55	45
rect	54	45	55	46
rect	54	46	55	47
rect	54	47	55	48
rect	54	48	55	49
rect	54	49	55	50
rect	54	50	55	51
rect	54	51	55	52
rect	54	52	55	53
rect	54	53	55	54
rect	54	54	55	55
rect	54	55	55	56
rect	54	56	55	57
rect	54	57	55	58
rect	54	58	55	59
rect	54	59	55	60
rect	54	60	55	61
rect	54	61	55	62
rect	54	62	55	63
rect	54	63	55	64
rect	54	64	55	65
rect	54	65	55	66
rect	54	66	55	67
rect	54	67	55	68
rect	54	68	55	69
rect	54	69	55	70
rect	54	70	55	71
rect	54	71	55	72
rect	54	72	55	73
rect	54	73	55	74
rect	54	74	55	75
rect	54	75	55	76
rect	54	76	55	77
rect	54	77	55	78
rect	54	78	55	79
rect	54	79	55	80
rect	54	80	55	81
rect	54	81	55	82
rect	54	82	55	83
rect	54	83	55	84
rect	54	84	55	85
rect	54	85	55	86
rect	54	86	55	87
rect	54	87	55	88
rect	54	88	55	89
rect	54	89	55	90
rect	54	90	55	91
rect	54	91	55	92
rect	54	92	55	93
rect	54	93	55	94
rect	54	94	55	95
rect	54	95	55	96
rect	54	96	55	97
rect	54	97	55	98
rect	54	98	55	99
rect	54	99	55	100
rect	54	100	55	101
rect	54	101	55	102
rect	54	102	55	103
rect	54	103	55	104
rect	54	104	55	105
rect	54	105	55	106
rect	54	106	55	107
rect	54	107	55	108
rect	54	108	55	109
rect	54	109	55	110
rect	54	110	55	111
rect	54	111	55	112
rect	54	112	55	113
rect	54	113	55	114
rect	54	114	55	115
rect	54	115	55	116
rect	54	116	55	117
rect	54	117	55	118
rect	54	118	55	119
rect	54	119	55	120
rect	54	120	55	121
rect	54	121	55	122
rect	54	122	55	123
rect	54	123	55	124
rect	54	124	55	125
rect	54	125	55	126
rect	54	126	55	127
rect	54	127	55	128
rect	54	128	55	129
rect	54	129	55	130
rect	54	130	55	131
rect	54	131	55	132
rect	54	132	55	133
rect	54	133	55	134
rect	54	134	55	135
rect	54	135	55	136
rect	54	136	55	137
rect	54	137	55	138
rect	54	138	55	139
rect	54	139	55	140
rect	54	140	55	141
rect	54	141	55	142
rect	54	142	55	143
rect	54	143	55	144
rect	54	144	55	145
rect	54	145	55	146
rect	54	146	55	147
rect	54	147	55	148
rect	54	148	55	149
rect	54	149	55	150
rect	54	150	55	151
rect	54	151	55	152
rect	54	152	55	153
rect	54	153	55	154
rect	54	154	55	155
rect	54	155	55	156
rect	54	156	55	157
rect	54	157	55	158
rect	54	158	55	159
rect	54	159	55	160
rect	54	160	55	161
rect	54	161	55	162
rect	54	162	55	163
rect	54	163	55	164
rect	54	164	55	165
rect	54	165	55	166
rect	54	166	55	167
rect	54	167	55	168
rect	54	168	55	169
rect	54	169	55	170
rect	54	170	55	171
rect	54	171	55	172
rect	54	172	55	173
rect	54	173	55	174
rect	54	174	55	175
rect	54	175	55	176
rect	54	176	55	177
rect	54	177	55	178
rect	54	178	55	179
rect	54	179	55	180
rect	54	180	55	181
rect	54	181	55	182
rect	54	182	55	183
rect	54	183	55	184
rect	54	184	55	185
rect	54	185	55	186
rect	54	186	55	187
rect	54	187	55	188
rect	54	188	55	189
rect	54	189	55	190
rect	54	190	55	191
rect	54	191	55	192
rect	54	192	55	193
rect	54	193	55	194
rect	54	194	55	195
rect	54	195	55	196
rect	54	196	55	197
rect	54	197	55	198
rect	54	198	55	199
rect	54	199	55	200
rect	54	200	55	201
rect	54	201	55	202
rect	54	202	55	203
rect	54	203	55	204
rect	54	204	55	205
rect	54	205	55	206
rect	54	206	55	207
rect	54	207	55	208
rect	54	208	55	209
rect	54	209	55	210
rect	54	210	55	211
rect	54	211	55	212
rect	54	212	55	213
rect	54	213	55	214
rect	54	214	55	215
rect	54	215	55	216
rect	54	216	55	217
rect	54	217	55	218
rect	54	218	55	219
rect	54	219	55	220
rect	54	220	55	221
rect	54	221	55	222
rect	54	222	55	223
rect	54	223	55	224
rect	54	224	55	225
rect	54	225	55	226
rect	54	226	55	227
rect	54	227	55	228
rect	54	228	55	229
rect	54	229	55	230
rect	54	230	55	231
rect	54	231	55	232
rect	54	232	55	233
rect	54	233	55	234
rect	54	234	55	235
rect	54	235	55	236
rect	54	236	55	237
rect	54	237	55	238
rect	54	238	55	239
rect	54	239	55	240
rect	54	240	55	241
rect	54	241	55	242
rect	54	242	55	243
rect	55	0	56	1
rect	55	1	56	2
rect	55	2	56	3
rect	55	3	56	4
rect	55	4	56	5
rect	55	5	56	6
rect	55	6	56	7
rect	55	7	56	8
rect	55	8	56	9
rect	55	9	56	10
rect	55	10	56	11
rect	55	11	56	12
rect	55	12	56	13
rect	55	13	56	14
rect	55	14	56	15
rect	55	15	56	16
rect	55	16	56	17
rect	55	17	56	18
rect	55	18	56	19
rect	55	19	56	20
rect	55	20	56	21
rect	55	21	56	22
rect	55	22	56	23
rect	55	23	56	24
rect	55	24	56	25
rect	55	25	56	26
rect	55	26	56	27
rect	55	27	56	28
rect	55	28	56	29
rect	55	29	56	30
rect	55	30	56	31
rect	55	31	56	32
rect	55	32	56	33
rect	55	33	56	34
rect	55	34	56	35
rect	55	35	56	36
rect	55	36	56	37
rect	55	37	56	38
rect	55	38	56	39
rect	55	39	56	40
rect	55	40	56	41
rect	55	41	56	42
rect	55	42	56	43
rect	55	43	56	44
rect	55	44	56	45
rect	55	45	56	46
rect	55	46	56	47
rect	55	47	56	48
rect	55	48	56	49
rect	55	49	56	50
rect	55	50	56	51
rect	55	51	56	52
rect	55	52	56	53
rect	55	53	56	54
rect	55	54	56	55
rect	55	55	56	56
rect	55	56	56	57
rect	55	57	56	58
rect	55	58	56	59
rect	55	59	56	60
rect	55	60	56	61
rect	55	61	56	62
rect	55	62	56	63
rect	55	63	56	64
rect	55	64	56	65
rect	55	65	56	66
rect	55	66	56	67
rect	55	67	56	68
rect	55	68	56	69
rect	55	69	56	70
rect	55	70	56	71
rect	55	71	56	72
rect	55	72	56	73
rect	55	73	56	74
rect	55	74	56	75
rect	55	75	56	76
rect	55	76	56	77
rect	55	77	56	78
rect	55	78	56	79
rect	55	79	56	80
rect	55	80	56	81
rect	55	81	56	82
rect	55	82	56	83
rect	55	83	56	84
rect	55	84	56	85
rect	55	85	56	86
rect	55	86	56	87
rect	55	87	56	88
rect	55	88	56	89
rect	55	89	56	90
rect	55	90	56	91
rect	55	91	56	92
rect	55	92	56	93
rect	55	93	56	94
rect	55	94	56	95
rect	55	95	56	96
rect	55	96	56	97
rect	55	97	56	98
rect	55	98	56	99
rect	55	99	56	100
rect	55	100	56	101
rect	55	101	56	102
rect	55	102	56	103
rect	55	103	56	104
rect	55	104	56	105
rect	55	105	56	106
rect	55	106	56	107
rect	55	107	56	108
rect	55	108	56	109
rect	55	109	56	110
rect	55	110	56	111
rect	55	111	56	112
rect	55	112	56	113
rect	55	113	56	114
rect	55	114	56	115
rect	55	115	56	116
rect	55	116	56	117
rect	55	117	56	118
rect	55	118	56	119
rect	55	119	56	120
rect	55	120	56	121
rect	55	121	56	122
rect	55	122	56	123
rect	55	123	56	124
rect	55	124	56	125
rect	55	125	56	126
rect	55	126	56	127
rect	55	127	56	128
rect	55	128	56	129
rect	55	129	56	130
rect	55	130	56	131
rect	55	131	56	132
rect	55	132	56	133
rect	55	133	56	134
rect	55	134	56	135
rect	55	135	56	136
rect	55	136	56	137
rect	55	137	56	138
rect	55	138	56	139
rect	55	139	56	140
rect	55	140	56	141
rect	55	141	56	142
rect	55	142	56	143
rect	55	143	56	144
rect	55	144	56	145
rect	55	145	56	146
rect	55	146	56	147
rect	55	147	56	148
rect	55	148	56	149
rect	55	149	56	150
rect	55	150	56	151
rect	55	151	56	152
rect	55	152	56	153
rect	55	153	56	154
rect	55	154	56	155
rect	55	155	56	156
rect	55	156	56	157
rect	55	157	56	158
rect	55	158	56	159
rect	55	159	56	160
rect	55	160	56	161
rect	55	161	56	162
rect	55	162	56	163
rect	55	163	56	164
rect	55	164	56	165
rect	55	165	56	166
rect	55	166	56	167
rect	55	167	56	168
rect	55	168	56	169
rect	55	169	56	170
rect	55	170	56	171
rect	55	171	56	172
rect	55	172	56	173
rect	55	173	56	174
rect	55	174	56	175
rect	55	175	56	176
rect	55	176	56	177
rect	55	177	56	178
rect	55	178	56	179
rect	55	179	56	180
rect	55	180	56	181
rect	55	181	56	182
rect	55	182	56	183
rect	55	183	56	184
rect	55	184	56	185
rect	55	185	56	186
rect	55	186	56	187
rect	55	187	56	188
rect	55	188	56	189
rect	55	189	56	190
rect	55	190	56	191
rect	55	191	56	192
rect	55	192	56	193
rect	55	193	56	194
rect	55	194	56	195
rect	55	195	56	196
rect	55	196	56	197
rect	55	197	56	198
rect	55	198	56	199
rect	55	199	56	200
rect	55	200	56	201
rect	55	201	56	202
rect	55	202	56	203
rect	55	203	56	204
rect	55	204	56	205
rect	55	205	56	206
rect	55	206	56	207
rect	55	207	56	208
rect	55	208	56	209
rect	55	209	56	210
rect	55	210	56	211
rect	55	211	56	212
rect	55	212	56	213
rect	55	213	56	214
rect	55	214	56	215
rect	55	215	56	216
rect	55	216	56	217
rect	55	217	56	218
rect	55	218	56	219
rect	55	219	56	220
rect	55	220	56	221
rect	55	221	56	222
rect	55	222	56	223
rect	55	223	56	224
rect	55	224	56	225
rect	55	225	56	226
rect	55	226	56	227
rect	55	227	56	228
rect	55	228	56	229
rect	55	229	56	230
rect	55	230	56	231
rect	55	231	56	232
rect	55	232	56	233
rect	55	233	56	234
rect	55	234	56	235
rect	55	235	56	236
rect	55	236	56	237
rect	55	237	56	238
rect	55	238	56	239
rect	55	239	56	240
rect	55	240	56	241
rect	55	241	56	242
rect	55	242	56	243
rect	56	0	57	1
rect	56	1	57	2
rect	56	2	57	3
rect	56	3	57	4
rect	56	4	57	5
rect	56	5	57	6
rect	56	6	57	7
rect	56	7	57	8
rect	56	8	57	9
rect	56	9	57	10
rect	56	10	57	11
rect	56	11	57	12
rect	56	12	57	13
rect	56	13	57	14
rect	56	14	57	15
rect	56	15	57	16
rect	56	16	57	17
rect	56	17	57	18
rect	56	18	57	19
rect	56	19	57	20
rect	56	20	57	21
rect	56	21	57	22
rect	56	22	57	23
rect	56	23	57	24
rect	56	24	57	25
rect	56	25	57	26
rect	56	26	57	27
rect	56	27	57	28
rect	56	28	57	29
rect	56	29	57	30
rect	56	30	57	31
rect	56	31	57	32
rect	56	32	57	33
rect	56	33	57	34
rect	56	34	57	35
rect	56	35	57	36
rect	56	36	57	37
rect	56	37	57	38
rect	56	38	57	39
rect	56	39	57	40
rect	56	40	57	41
rect	56	41	57	42
rect	56	42	57	43
rect	56	43	57	44
rect	56	44	57	45
rect	56	45	57	46
rect	56	46	57	47
rect	56	47	57	48
rect	56	48	57	49
rect	56	49	57	50
rect	56	50	57	51
rect	56	51	57	52
rect	56	52	57	53
rect	56	53	57	54
rect	56	54	57	55
rect	56	55	57	56
rect	56	56	57	57
rect	56	57	57	58
rect	56	58	57	59
rect	56	59	57	60
rect	56	60	57	61
rect	56	61	57	62
rect	56	62	57	63
rect	56	63	57	64
rect	56	64	57	65
rect	56	65	57	66
rect	56	66	57	67
rect	56	67	57	68
rect	56	68	57	69
rect	56	69	57	70
rect	56	70	57	71
rect	56	71	57	72
rect	56	72	57	73
rect	56	73	57	74
rect	56	74	57	75
rect	56	75	57	76
rect	56	76	57	77
rect	56	77	57	78
rect	56	78	57	79
rect	56	79	57	80
rect	56	80	57	81
rect	56	81	57	82
rect	56	82	57	83
rect	56	83	57	84
rect	56	84	57	85
rect	56	85	57	86
rect	56	86	57	87
rect	56	87	57	88
rect	56	88	57	89
rect	56	89	57	90
rect	56	90	57	91
rect	56	91	57	92
rect	56	92	57	93
rect	56	93	57	94
rect	56	94	57	95
rect	56	95	57	96
rect	56	96	57	97
rect	56	97	57	98
rect	56	98	57	99
rect	56	99	57	100
rect	56	100	57	101
rect	56	101	57	102
rect	56	102	57	103
rect	56	103	57	104
rect	56	104	57	105
rect	56	105	57	106
rect	56	106	57	107
rect	56	107	57	108
rect	56	108	57	109
rect	56	109	57	110
rect	56	110	57	111
rect	56	111	57	112
rect	56	112	57	113
rect	56	113	57	114
rect	56	114	57	115
rect	56	115	57	116
rect	56	116	57	117
rect	56	117	57	118
rect	56	118	57	119
rect	56	119	57	120
rect	56	120	57	121
rect	56	121	57	122
rect	56	122	57	123
rect	56	123	57	124
rect	56	124	57	125
rect	56	125	57	126
rect	56	126	57	127
rect	56	127	57	128
rect	56	128	57	129
rect	56	129	57	130
rect	56	130	57	131
rect	56	131	57	132
rect	56	132	57	133
rect	56	133	57	134
rect	56	134	57	135
rect	56	135	57	136
rect	56	136	57	137
rect	56	137	57	138
rect	56	138	57	139
rect	56	139	57	140
rect	56	140	57	141
rect	56	141	57	142
rect	56	142	57	143
rect	56	143	57	144
rect	56	144	57	145
rect	56	145	57	146
rect	56	146	57	147
rect	56	147	57	148
rect	56	148	57	149
rect	56	149	57	150
rect	56	150	57	151
rect	56	151	57	152
rect	56	152	57	153
rect	56	153	57	154
rect	56	154	57	155
rect	56	155	57	156
rect	56	156	57	157
rect	56	157	57	158
rect	56	158	57	159
rect	56	159	57	160
rect	56	160	57	161
rect	56	161	57	162
rect	56	162	57	163
rect	56	163	57	164
rect	56	164	57	165
rect	56	165	57	166
rect	56	166	57	167
rect	56	167	57	168
rect	56	168	57	169
rect	56	169	57	170
rect	56	170	57	171
rect	56	171	57	172
rect	56	172	57	173
rect	56	173	57	174
rect	56	174	57	175
rect	56	175	57	176
rect	56	176	57	177
rect	56	177	57	178
rect	56	178	57	179
rect	56	179	57	180
rect	56	180	57	181
rect	56	181	57	182
rect	56	182	57	183
rect	56	183	57	184
rect	56	184	57	185
rect	56	185	57	186
rect	56	186	57	187
rect	56	187	57	188
rect	56	188	57	189
rect	56	189	57	190
rect	56	190	57	191
rect	56	191	57	192
rect	56	192	57	193
rect	56	193	57	194
rect	56	194	57	195
rect	56	195	57	196
rect	56	196	57	197
rect	56	197	57	198
rect	56	198	57	199
rect	56	199	57	200
rect	56	200	57	201
rect	56	201	57	202
rect	56	202	57	203
rect	56	203	57	204
rect	56	204	57	205
rect	56	205	57	206
rect	56	206	57	207
rect	56	207	57	208
rect	56	208	57	209
rect	56	209	57	210
rect	56	210	57	211
rect	56	211	57	212
rect	56	212	57	213
rect	56	213	57	214
rect	56	214	57	215
rect	56	215	57	216
rect	56	216	57	217
rect	56	217	57	218
rect	56	218	57	219
rect	56	219	57	220
rect	56	220	57	221
rect	56	221	57	222
rect	56	222	57	223
rect	56	223	57	224
rect	56	224	57	225
rect	56	225	57	226
rect	56	226	57	227
rect	56	227	57	228
rect	56	228	57	229
rect	56	229	57	230
rect	56	230	57	231
rect	56	231	57	232
rect	56	232	57	233
rect	56	233	57	234
rect	56	234	57	235
rect	56	235	57	236
rect	56	236	57	237
rect	56	237	57	238
rect	56	238	57	239
rect	56	239	57	240
rect	56	240	57	241
rect	56	241	57	242
rect	56	242	57	243
rect	57	0	58	1
rect	57	1	58	2
rect	57	2	58	3
rect	57	3	58	4
rect	57	4	58	5
rect	57	5	58	6
rect	57	6	58	7
rect	57	7	58	8
rect	57	8	58	9
rect	57	9	58	10
rect	57	10	58	11
rect	57	11	58	12
rect	57	12	58	13
rect	57	13	58	14
rect	57	14	58	15
rect	57	15	58	16
rect	57	16	58	17
rect	57	17	58	18
rect	57	18	58	19
rect	57	19	58	20
rect	57	20	58	21
rect	57	21	58	22
rect	57	22	58	23
rect	57	23	58	24
rect	57	24	58	25
rect	57	25	58	26
rect	57	26	58	27
rect	57	27	58	28
rect	57	28	58	29
rect	57	29	58	30
rect	57	30	58	31
rect	57	31	58	32
rect	57	32	58	33
rect	57	33	58	34
rect	57	34	58	35
rect	57	35	58	36
rect	57	36	58	37
rect	57	37	58	38
rect	57	38	58	39
rect	57	39	58	40
rect	57	40	58	41
rect	57	41	58	42
rect	57	42	58	43
rect	57	43	58	44
rect	57	44	58	45
rect	57	45	58	46
rect	57	46	58	47
rect	57	47	58	48
rect	57	48	58	49
rect	57	49	58	50
rect	57	50	58	51
rect	57	51	58	52
rect	57	52	58	53
rect	57	53	58	54
rect	57	54	58	55
rect	57	55	58	56
rect	57	56	58	57
rect	57	57	58	58
rect	57	58	58	59
rect	57	59	58	60
rect	57	60	58	61
rect	57	61	58	62
rect	57	62	58	63
rect	57	63	58	64
rect	57	64	58	65
rect	57	65	58	66
rect	57	66	58	67
rect	57	67	58	68
rect	57	68	58	69
rect	57	69	58	70
rect	57	70	58	71
rect	57	71	58	72
rect	57	72	58	73
rect	57	73	58	74
rect	57	74	58	75
rect	57	75	58	76
rect	57	76	58	77
rect	57	77	58	78
rect	57	78	58	79
rect	57	79	58	80
rect	57	80	58	81
rect	57	81	58	82
rect	57	82	58	83
rect	57	83	58	84
rect	57	84	58	85
rect	57	85	58	86
rect	57	86	58	87
rect	57	87	58	88
rect	57	88	58	89
rect	57	89	58	90
rect	57	90	58	91
rect	57	91	58	92
rect	57	92	58	93
rect	57	93	58	94
rect	57	94	58	95
rect	57	95	58	96
rect	57	96	58	97
rect	57	97	58	98
rect	57	98	58	99
rect	57	99	58	100
rect	57	100	58	101
rect	57	101	58	102
rect	57	102	58	103
rect	57	103	58	104
rect	57	104	58	105
rect	57	105	58	106
rect	57	106	58	107
rect	57	107	58	108
rect	57	108	58	109
rect	57	109	58	110
rect	57	110	58	111
rect	57	111	58	112
rect	57	112	58	113
rect	57	113	58	114
rect	57	114	58	115
rect	57	115	58	116
rect	57	116	58	117
rect	57	117	58	118
rect	57	118	58	119
rect	57	119	58	120
rect	57	120	58	121
rect	57	121	58	122
rect	57	122	58	123
rect	57	123	58	124
rect	57	124	58	125
rect	57	125	58	126
rect	57	126	58	127
rect	57	127	58	128
rect	57	128	58	129
rect	57	129	58	130
rect	57	130	58	131
rect	57	131	58	132
rect	57	132	58	133
rect	57	133	58	134
rect	57	134	58	135
rect	57	135	58	136
rect	57	136	58	137
rect	57	137	58	138
rect	57	138	58	139
rect	57	139	58	140
rect	57	140	58	141
rect	57	141	58	142
rect	57	142	58	143
rect	57	143	58	144
rect	57	144	58	145
rect	57	145	58	146
rect	57	146	58	147
rect	57	147	58	148
rect	57	148	58	149
rect	57	149	58	150
rect	57	150	58	151
rect	57	151	58	152
rect	57	152	58	153
rect	57	153	58	154
rect	57	154	58	155
rect	57	155	58	156
rect	57	156	58	157
rect	57	157	58	158
rect	57	158	58	159
rect	57	159	58	160
rect	57	160	58	161
rect	57	161	58	162
rect	57	162	58	163
rect	57	163	58	164
rect	57	164	58	165
rect	57	165	58	166
rect	57	166	58	167
rect	57	167	58	168
rect	57	168	58	169
rect	57	169	58	170
rect	57	170	58	171
rect	57	171	58	172
rect	57	172	58	173
rect	57	173	58	174
rect	57	174	58	175
rect	57	175	58	176
rect	57	176	58	177
rect	57	177	58	178
rect	57	178	58	179
rect	57	179	58	180
rect	57	180	58	181
rect	57	181	58	182
rect	57	182	58	183
rect	57	183	58	184
rect	57	184	58	185
rect	57	185	58	186
rect	57	186	58	187
rect	57	187	58	188
rect	57	188	58	189
rect	57	189	58	190
rect	57	190	58	191
rect	57	191	58	192
rect	57	192	58	193
rect	57	193	58	194
rect	57	194	58	195
rect	57	195	58	196
rect	57	196	58	197
rect	57	197	58	198
rect	57	198	58	199
rect	57	199	58	200
rect	57	200	58	201
rect	57	201	58	202
rect	57	202	58	203
rect	57	203	58	204
rect	57	204	58	205
rect	57	205	58	206
rect	57	206	58	207
rect	57	207	58	208
rect	57	208	58	209
rect	57	209	58	210
rect	57	210	58	211
rect	57	211	58	212
rect	57	212	58	213
rect	57	213	58	214
rect	57	214	58	215
rect	57	215	58	216
rect	57	216	58	217
rect	57	217	58	218
rect	57	218	58	219
rect	57	219	58	220
rect	57	220	58	221
rect	57	221	58	222
rect	57	222	58	223
rect	57	223	58	224
rect	57	224	58	225
rect	57	225	58	226
rect	57	226	58	227
rect	57	227	58	228
rect	57	228	58	229
rect	57	229	58	230
rect	57	230	58	231
rect	57	231	58	232
rect	57	232	58	233
rect	57	233	58	234
rect	57	234	58	235
rect	57	235	58	236
rect	57	236	58	237
rect	57	237	58	238
rect	57	238	58	239
rect	57	239	58	240
rect	57	240	58	241
rect	57	241	58	242
rect	57	242	58	243
rect	75	0	76	1
rect	75	1	76	2
rect	75	2	76	3
rect	75	3	76	4
rect	75	4	76	5
rect	75	5	76	6
rect	75	6	76	7
rect	75	7	76	8
rect	75	8	76	9
rect	75	9	76	10
rect	75	10	76	11
rect	75	11	76	12
rect	75	12	76	13
rect	75	13	76	14
rect	75	14	76	15
rect	75	15	76	16
rect	75	16	76	17
rect	75	17	76	18
rect	75	18	76	19
rect	75	19	76	20
rect	75	20	76	21
rect	75	21	76	22
rect	75	22	76	23
rect	75	23	76	24
rect	75	24	76	25
rect	75	25	76	26
rect	75	26	76	27
rect	75	27	76	28
rect	75	28	76	29
rect	75	29	76	30
rect	75	30	76	31
rect	75	31	76	32
rect	75	32	76	33
rect	75	33	76	34
rect	75	34	76	35
rect	75	35	76	36
rect	75	36	76	37
rect	75	37	76	38
rect	75	38	76	39
rect	75	39	76	40
rect	75	40	76	41
rect	75	41	76	42
rect	75	42	76	43
rect	75	43	76	44
rect	75	44	76	45
rect	75	45	76	46
rect	75	46	76	47
rect	75	47	76	48
rect	75	48	76	49
rect	75	49	76	50
rect	75	50	76	51
rect	75	51	76	52
rect	75	52	76	53
rect	75	53	76	54
rect	75	54	76	55
rect	75	55	76	56
rect	75	56	76	57
rect	75	57	76	58
rect	75	58	76	59
rect	75	59	76	60
rect	75	60	76	61
rect	75	61	76	62
rect	75	62	76	63
rect	75	63	76	64
rect	75	64	76	65
rect	75	65	76	66
rect	75	66	76	67
rect	75	67	76	68
rect	75	68	76	69
rect	75	69	76	70
rect	75	70	76	71
rect	75	71	76	72
rect	75	72	76	73
rect	75	73	76	74
rect	75	74	76	75
rect	75	75	76	76
rect	75	76	76	77
rect	75	77	76	78
rect	75	78	76	79
rect	75	79	76	80
rect	75	80	76	81
rect	75	81	76	82
rect	75	82	76	83
rect	75	83	76	84
rect	75	84	76	85
rect	75	85	76	86
rect	75	86	76	87
rect	75	87	76	88
rect	75	88	76	89
rect	75	89	76	90
rect	75	90	76	91
rect	75	91	76	92
rect	75	92	76	93
rect	75	93	76	94
rect	75	94	76	95
rect	75	95	76	96
rect	75	96	76	97
rect	75	97	76	98
rect	75	98	76	99
rect	75	99	76	100
rect	75	100	76	101
rect	75	101	76	102
rect	75	102	76	103
rect	75	103	76	104
rect	75	104	76	105
rect	75	105	76	106
rect	75	106	76	107
rect	75	107	76	108
rect	75	108	76	109
rect	75	109	76	110
rect	75	110	76	111
rect	75	111	76	112
rect	75	112	76	113
rect	75	113	76	114
rect	75	114	76	115
rect	75	115	76	116
rect	75	116	76	117
rect	75	117	76	118
rect	75	118	76	119
rect	75	119	76	120
rect	75	120	76	121
rect	75	121	76	122
rect	75	122	76	123
rect	75	123	76	124
rect	75	124	76	125
rect	75	125	76	126
rect	75	126	76	127
rect	75	127	76	128
rect	75	128	76	129
rect	75	129	76	130
rect	75	130	76	131
rect	75	131	76	132
rect	75	132	76	133
rect	75	133	76	134
rect	75	134	76	135
rect	75	135	76	136
rect	75	136	76	137
rect	75	137	76	138
rect	75	138	76	139
rect	75	139	76	140
rect	75	140	76	141
rect	75	141	76	142
rect	75	142	76	143
rect	75	143	76	144
rect	75	144	76	145
rect	75	145	76	146
rect	75	146	76	147
rect	75	147	76	148
rect	75	148	76	149
rect	75	149	76	150
rect	75	150	76	151
rect	75	151	76	152
rect	75	152	76	153
rect	75	153	76	154
rect	75	154	76	155
rect	75	155	76	156
rect	75	156	76	157
rect	75	157	76	158
rect	75	158	76	159
rect	75	159	76	160
rect	75	160	76	161
rect	75	161	76	162
rect	75	162	76	163
rect	75	163	76	164
rect	75	164	76	165
rect	75	165	76	166
rect	75	166	76	167
rect	75	167	76	168
rect	75	168	76	169
rect	75	169	76	170
rect	75	170	76	171
rect	75	171	76	172
rect	75	172	76	173
rect	75	173	76	174
rect	75	174	76	175
rect	75	175	76	176
rect	75	176	76	177
rect	75	177	76	178
rect	75	178	76	179
rect	75	179	76	180
rect	75	180	76	181
rect	75	181	76	182
rect	75	182	76	183
rect	75	183	76	184
rect	75	184	76	185
rect	75	185	76	186
rect	75	186	76	187
rect	75	187	76	188
rect	75	188	76	189
rect	75	189	76	190
rect	75	190	76	191
rect	75	191	76	192
rect	75	192	76	193
rect	75	193	76	194
rect	75	194	76	195
rect	75	195	76	196
rect	75	196	76	197
rect	75	197	76	198
rect	75	198	76	199
rect	75	199	76	200
rect	75	200	76	201
rect	75	201	76	202
rect	75	202	76	203
rect	75	203	76	204
rect	75	204	76	205
rect	75	205	76	206
rect	75	206	76	207
rect	75	207	76	208
rect	75	208	76	209
rect	75	209	76	210
rect	75	210	76	211
rect	75	211	76	212
rect	75	212	76	213
rect	75	213	76	214
rect	75	214	76	215
rect	75	215	76	216
rect	75	216	76	217
rect	75	217	76	218
rect	75	218	76	219
rect	75	219	76	220
rect	75	220	76	221
rect	75	221	76	222
rect	75	222	76	223
rect	75	223	76	224
rect	75	224	76	225
rect	75	225	76	226
rect	75	226	76	227
rect	75	227	76	228
rect	75	228	76	229
rect	75	229	76	230
rect	75	230	76	231
rect	75	231	76	232
rect	75	232	76	233
rect	75	233	76	234
rect	75	234	76	235
rect	75	235	76	236
rect	75	236	76	237
rect	75	237	76	238
rect	75	238	76	239
rect	75	239	76	240
rect	75	240	76	241
rect	75	241	76	242
rect	75	242	76	243
rect	75	243	76	244
rect	75	244	76	245
rect	75	245	76	246
rect	75	246	76	247
rect	75	247	76	248
rect	75	248	76	249
rect	75	249	76	250
rect	75	250	76	251
rect	75	251	76	252
rect	75	252	76	253
rect	75	253	76	254
rect	75	254	76	255
rect	75	255	76	256
rect	75	256	76	257
rect	75	257	76	258
rect	75	258	76	259
rect	75	259	76	260
rect	75	260	76	261
rect	75	261	76	262
rect	75	262	76	263
rect	75	263	76	264
rect	75	264	76	265
rect	75	265	76	266
rect	75	266	76	267
rect	75	267	76	268
rect	75	268	76	269
rect	75	269	76	270
rect	75	270	76	271
rect	75	271	76	272
rect	75	272	76	273
rect	75	273	76	274
rect	75	274	76	275
rect	75	275	76	276
rect	75	276	76	277
rect	75	277	76	278
rect	75	278	76	279
rect	75	279	76	280
rect	75	280	76	281
rect	75	281	76	282
rect	75	282	76	283
rect	75	283	76	284
rect	75	284	76	285
rect	75	285	76	286
rect	75	286	76	287
rect	75	287	76	288
rect	75	288	76	289
rect	75	289	76	290
rect	75	290	76	291
rect	76	0	77	1
rect	76	1	77	2
rect	76	2	77	3
rect	76	3	77	4
rect	76	4	77	5
rect	76	5	77	6
rect	76	6	77	7
rect	76	7	77	8
rect	76	8	77	9
rect	76	9	77	10
rect	76	10	77	11
rect	76	11	77	12
rect	76	12	77	13
rect	76	13	77	14
rect	76	14	77	15
rect	76	15	77	16
rect	76	16	77	17
rect	76	17	77	18
rect	76	18	77	19
rect	76	19	77	20
rect	76	20	77	21
rect	76	21	77	22
rect	76	22	77	23
rect	76	23	77	24
rect	76	24	77	25
rect	76	25	77	26
rect	76	26	77	27
rect	76	27	77	28
rect	76	28	77	29
rect	76	29	77	30
rect	76	30	77	31
rect	76	31	77	32
rect	76	32	77	33
rect	76	33	77	34
rect	76	34	77	35
rect	76	35	77	36
rect	76	36	77	37
rect	76	37	77	38
rect	76	38	77	39
rect	76	39	77	40
rect	76	40	77	41
rect	76	41	77	42
rect	76	42	77	43
rect	76	43	77	44
rect	76	44	77	45
rect	76	45	77	46
rect	76	46	77	47
rect	76	47	77	48
rect	76	48	77	49
rect	76	49	77	50
rect	76	50	77	51
rect	76	51	77	52
rect	76	52	77	53
rect	76	53	77	54
rect	76	54	77	55
rect	76	55	77	56
rect	76	56	77	57
rect	76	57	77	58
rect	76	58	77	59
rect	76	59	77	60
rect	76	60	77	61
rect	76	61	77	62
rect	76	62	77	63
rect	76	63	77	64
rect	76	64	77	65
rect	76	65	77	66
rect	76	66	77	67
rect	76	67	77	68
rect	76	68	77	69
rect	76	69	77	70
rect	76	70	77	71
rect	76	71	77	72
rect	76	72	77	73
rect	76	73	77	74
rect	76	74	77	75
rect	76	75	77	76
rect	76	76	77	77
rect	76	77	77	78
rect	76	78	77	79
rect	76	79	77	80
rect	76	80	77	81
rect	76	81	77	82
rect	76	82	77	83
rect	76	83	77	84
rect	76	84	77	85
rect	76	85	77	86
rect	76	86	77	87
rect	76	87	77	88
rect	76	88	77	89
rect	76	89	77	90
rect	76	90	77	91
rect	76	91	77	92
rect	76	92	77	93
rect	76	93	77	94
rect	76	94	77	95
rect	76	95	77	96
rect	76	96	77	97
rect	76	97	77	98
rect	76	98	77	99
rect	76	99	77	100
rect	76	100	77	101
rect	76	101	77	102
rect	76	102	77	103
rect	76	103	77	104
rect	76	104	77	105
rect	76	105	77	106
rect	76	106	77	107
rect	76	107	77	108
rect	76	108	77	109
rect	76	109	77	110
rect	76	110	77	111
rect	76	111	77	112
rect	76	112	77	113
rect	76	113	77	114
rect	76	114	77	115
rect	76	115	77	116
rect	76	116	77	117
rect	76	117	77	118
rect	76	118	77	119
rect	76	119	77	120
rect	76	120	77	121
rect	76	121	77	122
rect	76	122	77	123
rect	76	123	77	124
rect	76	124	77	125
rect	76	125	77	126
rect	76	126	77	127
rect	76	127	77	128
rect	76	128	77	129
rect	76	129	77	130
rect	76	130	77	131
rect	76	131	77	132
rect	76	132	77	133
rect	76	133	77	134
rect	76	134	77	135
rect	76	135	77	136
rect	76	136	77	137
rect	76	137	77	138
rect	76	138	77	139
rect	76	139	77	140
rect	76	140	77	141
rect	76	141	77	142
rect	76	142	77	143
rect	76	143	77	144
rect	76	144	77	145
rect	76	145	77	146
rect	76	146	77	147
rect	76	147	77	148
rect	76	148	77	149
rect	76	149	77	150
rect	76	150	77	151
rect	76	151	77	152
rect	76	152	77	153
rect	76	153	77	154
rect	76	154	77	155
rect	76	155	77	156
rect	76	156	77	157
rect	76	157	77	158
rect	76	158	77	159
rect	76	159	77	160
rect	76	160	77	161
rect	76	161	77	162
rect	76	162	77	163
rect	76	163	77	164
rect	76	164	77	165
rect	76	165	77	166
rect	76	166	77	167
rect	76	167	77	168
rect	76	168	77	169
rect	76	169	77	170
rect	76	170	77	171
rect	76	171	77	172
rect	76	172	77	173
rect	76	173	77	174
rect	76	174	77	175
rect	76	175	77	176
rect	76	176	77	177
rect	76	177	77	178
rect	76	178	77	179
rect	76	179	77	180
rect	76	180	77	181
rect	76	181	77	182
rect	76	182	77	183
rect	76	183	77	184
rect	76	184	77	185
rect	76	185	77	186
rect	76	186	77	187
rect	76	187	77	188
rect	76	188	77	189
rect	76	189	77	190
rect	76	190	77	191
rect	76	191	77	192
rect	76	192	77	193
rect	76	193	77	194
rect	76	194	77	195
rect	76	195	77	196
rect	76	196	77	197
rect	76	197	77	198
rect	76	198	77	199
rect	76	199	77	200
rect	76	200	77	201
rect	76	201	77	202
rect	76	202	77	203
rect	76	203	77	204
rect	76	204	77	205
rect	76	205	77	206
rect	76	206	77	207
rect	76	207	77	208
rect	76	208	77	209
rect	76	209	77	210
rect	76	210	77	211
rect	76	211	77	212
rect	76	212	77	213
rect	76	213	77	214
rect	76	214	77	215
rect	76	215	77	216
rect	76	216	77	217
rect	76	217	77	218
rect	76	218	77	219
rect	76	219	77	220
rect	76	220	77	221
rect	76	221	77	222
rect	76	222	77	223
rect	76	223	77	224
rect	76	224	77	225
rect	76	225	77	226
rect	76	226	77	227
rect	76	227	77	228
rect	76	228	77	229
rect	76	229	77	230
rect	76	230	77	231
rect	76	231	77	232
rect	76	232	77	233
rect	76	233	77	234
rect	76	234	77	235
rect	76	235	77	236
rect	76	236	77	237
rect	76	237	77	238
rect	76	238	77	239
rect	76	239	77	240
rect	76	240	77	241
rect	76	241	77	242
rect	76	242	77	243
rect	76	243	77	244
rect	76	244	77	245
rect	76	245	77	246
rect	76	246	77	247
rect	76	247	77	248
rect	76	248	77	249
rect	76	249	77	250
rect	76	250	77	251
rect	76	251	77	252
rect	76	252	77	253
rect	76	253	77	254
rect	76	254	77	255
rect	76	255	77	256
rect	76	256	77	257
rect	76	257	77	258
rect	76	258	77	259
rect	76	259	77	260
rect	76	260	77	261
rect	76	261	77	262
rect	76	262	77	263
rect	76	263	77	264
rect	76	264	77	265
rect	76	265	77	266
rect	76	266	77	267
rect	76	267	77	268
rect	76	268	77	269
rect	76	269	77	270
rect	76	270	77	271
rect	76	271	77	272
rect	76	272	77	273
rect	76	273	77	274
rect	76	274	77	275
rect	76	275	77	276
rect	76	276	77	277
rect	76	277	77	278
rect	76	278	77	279
rect	76	279	77	280
rect	76	280	77	281
rect	76	281	77	282
rect	76	282	77	283
rect	76	283	77	284
rect	76	284	77	285
rect	76	285	77	286
rect	76	286	77	287
rect	76	287	77	288
rect	76	288	77	289
rect	76	289	77	290
rect	76	290	77	291
rect	77	0	78	1
rect	77	1	78	2
rect	77	2	78	3
rect	77	3	78	4
rect	77	4	78	5
rect	77	5	78	6
rect	77	6	78	7
rect	77	7	78	8
rect	77	8	78	9
rect	77	9	78	10
rect	77	10	78	11
rect	77	11	78	12
rect	77	12	78	13
rect	77	13	78	14
rect	77	14	78	15
rect	77	15	78	16
rect	77	16	78	17
rect	77	17	78	18
rect	77	18	78	19
rect	77	19	78	20
rect	77	20	78	21
rect	77	21	78	22
rect	77	22	78	23
rect	77	23	78	24
rect	77	24	78	25
rect	77	25	78	26
rect	77	26	78	27
rect	77	27	78	28
rect	77	28	78	29
rect	77	29	78	30
rect	77	30	78	31
rect	77	31	78	32
rect	77	32	78	33
rect	77	33	78	34
rect	77	34	78	35
rect	77	35	78	36
rect	77	36	78	37
rect	77	37	78	38
rect	77	38	78	39
rect	77	39	78	40
rect	77	40	78	41
rect	77	41	78	42
rect	77	42	78	43
rect	77	43	78	44
rect	77	44	78	45
rect	77	45	78	46
rect	77	46	78	47
rect	77	47	78	48
rect	77	48	78	49
rect	77	49	78	50
rect	77	50	78	51
rect	77	51	78	52
rect	77	52	78	53
rect	77	53	78	54
rect	77	54	78	55
rect	77	55	78	56
rect	77	56	78	57
rect	77	57	78	58
rect	77	58	78	59
rect	77	59	78	60
rect	77	60	78	61
rect	77	61	78	62
rect	77	62	78	63
rect	77	63	78	64
rect	77	64	78	65
rect	77	65	78	66
rect	77	66	78	67
rect	77	67	78	68
rect	77	68	78	69
rect	77	69	78	70
rect	77	70	78	71
rect	77	71	78	72
rect	77	72	78	73
rect	77	73	78	74
rect	77	74	78	75
rect	77	75	78	76
rect	77	76	78	77
rect	77	77	78	78
rect	77	78	78	79
rect	77	79	78	80
rect	77	80	78	81
rect	77	81	78	82
rect	77	82	78	83
rect	77	83	78	84
rect	77	84	78	85
rect	77	85	78	86
rect	77	86	78	87
rect	77	87	78	88
rect	77	88	78	89
rect	77	89	78	90
rect	77	90	78	91
rect	77	91	78	92
rect	77	92	78	93
rect	77	93	78	94
rect	77	94	78	95
rect	77	95	78	96
rect	77	96	78	97
rect	77	97	78	98
rect	77	98	78	99
rect	77	99	78	100
rect	77	100	78	101
rect	77	101	78	102
rect	77	102	78	103
rect	77	103	78	104
rect	77	104	78	105
rect	77	105	78	106
rect	77	106	78	107
rect	77	107	78	108
rect	77	108	78	109
rect	77	109	78	110
rect	77	110	78	111
rect	77	111	78	112
rect	77	112	78	113
rect	77	113	78	114
rect	77	114	78	115
rect	77	115	78	116
rect	77	116	78	117
rect	77	117	78	118
rect	77	118	78	119
rect	77	119	78	120
rect	77	120	78	121
rect	77	121	78	122
rect	77	122	78	123
rect	77	123	78	124
rect	77	124	78	125
rect	77	125	78	126
rect	77	126	78	127
rect	77	127	78	128
rect	77	128	78	129
rect	77	129	78	130
rect	77	130	78	131
rect	77	131	78	132
rect	77	132	78	133
rect	77	133	78	134
rect	77	134	78	135
rect	77	135	78	136
rect	77	136	78	137
rect	77	137	78	138
rect	77	138	78	139
rect	77	139	78	140
rect	77	140	78	141
rect	77	141	78	142
rect	77	142	78	143
rect	77	143	78	144
rect	77	144	78	145
rect	77	145	78	146
rect	77	146	78	147
rect	77	147	78	148
rect	77	148	78	149
rect	77	149	78	150
rect	77	150	78	151
rect	77	151	78	152
rect	77	152	78	153
rect	77	153	78	154
rect	77	154	78	155
rect	77	155	78	156
rect	77	156	78	157
rect	77	157	78	158
rect	77	158	78	159
rect	77	159	78	160
rect	77	160	78	161
rect	77	161	78	162
rect	77	162	78	163
rect	77	163	78	164
rect	77	164	78	165
rect	77	165	78	166
rect	77	166	78	167
rect	77	167	78	168
rect	77	168	78	169
rect	77	169	78	170
rect	77	170	78	171
rect	77	171	78	172
rect	77	172	78	173
rect	77	173	78	174
rect	77	174	78	175
rect	77	175	78	176
rect	77	176	78	177
rect	77	177	78	178
rect	77	178	78	179
rect	77	179	78	180
rect	77	180	78	181
rect	77	181	78	182
rect	77	182	78	183
rect	77	183	78	184
rect	77	184	78	185
rect	77	185	78	186
rect	77	186	78	187
rect	77	187	78	188
rect	77	188	78	189
rect	77	189	78	190
rect	77	190	78	191
rect	77	191	78	192
rect	77	192	78	193
rect	77	193	78	194
rect	77	194	78	195
rect	77	195	78	196
rect	77	196	78	197
rect	77	197	78	198
rect	77	198	78	199
rect	77	199	78	200
rect	77	200	78	201
rect	77	201	78	202
rect	77	202	78	203
rect	77	203	78	204
rect	77	204	78	205
rect	77	205	78	206
rect	77	206	78	207
rect	77	207	78	208
rect	77	208	78	209
rect	77	209	78	210
rect	77	210	78	211
rect	77	211	78	212
rect	77	212	78	213
rect	77	213	78	214
rect	77	214	78	215
rect	77	215	78	216
rect	77	216	78	217
rect	77	217	78	218
rect	77	218	78	219
rect	77	219	78	220
rect	77	220	78	221
rect	77	221	78	222
rect	77	222	78	223
rect	77	223	78	224
rect	77	224	78	225
rect	77	225	78	226
rect	77	226	78	227
rect	77	227	78	228
rect	77	228	78	229
rect	77	229	78	230
rect	77	230	78	231
rect	77	231	78	232
rect	77	232	78	233
rect	77	233	78	234
rect	77	234	78	235
rect	77	235	78	236
rect	77	236	78	237
rect	77	237	78	238
rect	77	238	78	239
rect	77	239	78	240
rect	77	240	78	241
rect	77	241	78	242
rect	77	242	78	243
rect	77	243	78	244
rect	77	244	78	245
rect	77	245	78	246
rect	77	246	78	247
rect	77	247	78	248
rect	77	248	78	249
rect	77	249	78	250
rect	77	250	78	251
rect	77	251	78	252
rect	77	252	78	253
rect	77	253	78	254
rect	77	254	78	255
rect	77	255	78	256
rect	77	256	78	257
rect	77	257	78	258
rect	77	258	78	259
rect	77	259	78	260
rect	77	260	78	261
rect	77	261	78	262
rect	77	262	78	263
rect	77	263	78	264
rect	77	264	78	265
rect	77	265	78	266
rect	77	266	78	267
rect	77	267	78	268
rect	77	268	78	269
rect	77	269	78	270
rect	77	270	78	271
rect	77	271	78	272
rect	77	272	78	273
rect	77	273	78	274
rect	77	274	78	275
rect	77	275	78	276
rect	77	276	78	277
rect	77	277	78	278
rect	77	278	78	279
rect	77	279	78	280
rect	77	280	78	281
rect	77	281	78	282
rect	77	282	78	283
rect	77	283	78	284
rect	77	284	78	285
rect	77	285	78	286
rect	77	286	78	287
rect	77	287	78	288
rect	77	288	78	289
rect	77	289	78	290
rect	77	290	78	291
rect	78	0	79	1
rect	78	1	79	2
rect	78	2	79	3
rect	78	3	79	4
rect	78	4	79	5
rect	78	5	79	6
rect	78	6	79	7
rect	78	7	79	8
rect	78	8	79	9
rect	78	9	79	10
rect	78	10	79	11
rect	78	11	79	12
rect	78	12	79	13
rect	78	13	79	14
rect	78	14	79	15
rect	78	15	79	16
rect	78	16	79	17
rect	78	17	79	18
rect	78	18	79	19
rect	78	19	79	20
rect	78	20	79	21
rect	78	21	79	22
rect	78	22	79	23
rect	78	23	79	24
rect	78	24	79	25
rect	78	25	79	26
rect	78	26	79	27
rect	78	27	79	28
rect	78	28	79	29
rect	78	29	79	30
rect	78	30	79	31
rect	78	31	79	32
rect	78	32	79	33
rect	78	33	79	34
rect	78	34	79	35
rect	78	35	79	36
rect	78	36	79	37
rect	78	37	79	38
rect	78	38	79	39
rect	78	39	79	40
rect	78	40	79	41
rect	78	41	79	42
rect	78	42	79	43
rect	78	43	79	44
rect	78	44	79	45
rect	78	45	79	46
rect	78	46	79	47
rect	78	47	79	48
rect	78	48	79	49
rect	78	49	79	50
rect	78	50	79	51
rect	78	51	79	52
rect	78	52	79	53
rect	78	53	79	54
rect	78	54	79	55
rect	78	55	79	56
rect	78	56	79	57
rect	78	57	79	58
rect	78	58	79	59
rect	78	59	79	60
rect	78	60	79	61
rect	78	61	79	62
rect	78	62	79	63
rect	78	63	79	64
rect	78	64	79	65
rect	78	65	79	66
rect	78	66	79	67
rect	78	67	79	68
rect	78	68	79	69
rect	78	69	79	70
rect	78	70	79	71
rect	78	71	79	72
rect	78	72	79	73
rect	78	73	79	74
rect	78	74	79	75
rect	78	75	79	76
rect	78	76	79	77
rect	78	77	79	78
rect	78	78	79	79
rect	78	79	79	80
rect	78	80	79	81
rect	78	81	79	82
rect	78	82	79	83
rect	78	83	79	84
rect	78	84	79	85
rect	78	85	79	86
rect	78	86	79	87
rect	78	87	79	88
rect	78	88	79	89
rect	78	89	79	90
rect	78	90	79	91
rect	78	91	79	92
rect	78	92	79	93
rect	78	93	79	94
rect	78	94	79	95
rect	78	95	79	96
rect	78	96	79	97
rect	78	97	79	98
rect	78	98	79	99
rect	78	99	79	100
rect	78	100	79	101
rect	78	101	79	102
rect	78	102	79	103
rect	78	103	79	104
rect	78	104	79	105
rect	78	105	79	106
rect	78	106	79	107
rect	78	107	79	108
rect	78	108	79	109
rect	78	109	79	110
rect	78	110	79	111
rect	78	111	79	112
rect	78	112	79	113
rect	78	113	79	114
rect	78	114	79	115
rect	78	115	79	116
rect	78	116	79	117
rect	78	117	79	118
rect	78	118	79	119
rect	78	119	79	120
rect	78	120	79	121
rect	78	121	79	122
rect	78	122	79	123
rect	78	123	79	124
rect	78	124	79	125
rect	78	125	79	126
rect	78	126	79	127
rect	78	127	79	128
rect	78	128	79	129
rect	78	129	79	130
rect	78	130	79	131
rect	78	131	79	132
rect	78	132	79	133
rect	78	133	79	134
rect	78	134	79	135
rect	78	135	79	136
rect	78	136	79	137
rect	78	137	79	138
rect	78	138	79	139
rect	78	139	79	140
rect	78	140	79	141
rect	78	141	79	142
rect	78	142	79	143
rect	78	143	79	144
rect	78	144	79	145
rect	78	145	79	146
rect	78	146	79	147
rect	78	147	79	148
rect	78	148	79	149
rect	78	149	79	150
rect	78	150	79	151
rect	78	151	79	152
rect	78	152	79	153
rect	78	153	79	154
rect	78	154	79	155
rect	78	155	79	156
rect	78	156	79	157
rect	78	157	79	158
rect	78	158	79	159
rect	78	159	79	160
rect	78	160	79	161
rect	78	161	79	162
rect	78	162	79	163
rect	78	163	79	164
rect	78	164	79	165
rect	78	165	79	166
rect	78	166	79	167
rect	78	167	79	168
rect	78	168	79	169
rect	78	169	79	170
rect	78	170	79	171
rect	78	171	79	172
rect	78	172	79	173
rect	78	173	79	174
rect	78	174	79	175
rect	78	175	79	176
rect	78	176	79	177
rect	78	177	79	178
rect	78	178	79	179
rect	78	179	79	180
rect	78	180	79	181
rect	78	181	79	182
rect	78	182	79	183
rect	78	183	79	184
rect	78	184	79	185
rect	78	185	79	186
rect	78	186	79	187
rect	78	187	79	188
rect	78	188	79	189
rect	78	189	79	190
rect	78	190	79	191
rect	78	191	79	192
rect	78	192	79	193
rect	78	193	79	194
rect	78	194	79	195
rect	78	195	79	196
rect	78	196	79	197
rect	78	197	79	198
rect	78	198	79	199
rect	78	199	79	200
rect	78	200	79	201
rect	78	201	79	202
rect	78	202	79	203
rect	78	203	79	204
rect	78	204	79	205
rect	78	205	79	206
rect	78	206	79	207
rect	78	207	79	208
rect	78	208	79	209
rect	78	209	79	210
rect	78	210	79	211
rect	78	211	79	212
rect	78	212	79	213
rect	78	213	79	214
rect	78	214	79	215
rect	78	215	79	216
rect	78	216	79	217
rect	78	217	79	218
rect	78	218	79	219
rect	78	219	79	220
rect	78	220	79	221
rect	78	221	79	222
rect	78	222	79	223
rect	78	223	79	224
rect	78	224	79	225
rect	78	225	79	226
rect	78	226	79	227
rect	78	227	79	228
rect	78	228	79	229
rect	78	229	79	230
rect	78	230	79	231
rect	78	231	79	232
rect	78	232	79	233
rect	78	233	79	234
rect	78	234	79	235
rect	78	235	79	236
rect	78	236	79	237
rect	78	237	79	238
rect	78	238	79	239
rect	78	239	79	240
rect	78	240	79	241
rect	78	241	79	242
rect	78	242	79	243
rect	78	243	79	244
rect	78	244	79	245
rect	78	245	79	246
rect	78	246	79	247
rect	78	247	79	248
rect	78	248	79	249
rect	78	249	79	250
rect	78	250	79	251
rect	78	251	79	252
rect	78	252	79	253
rect	78	253	79	254
rect	78	254	79	255
rect	78	255	79	256
rect	78	256	79	257
rect	78	257	79	258
rect	78	258	79	259
rect	78	259	79	260
rect	78	260	79	261
rect	78	261	79	262
rect	78	262	79	263
rect	78	263	79	264
rect	78	264	79	265
rect	78	265	79	266
rect	78	266	79	267
rect	78	267	79	268
rect	78	268	79	269
rect	78	269	79	270
rect	78	270	79	271
rect	78	271	79	272
rect	78	272	79	273
rect	78	273	79	274
rect	78	274	79	275
rect	78	275	79	276
rect	78	276	79	277
rect	78	277	79	278
rect	78	278	79	279
rect	78	279	79	280
rect	78	280	79	281
rect	78	281	79	282
rect	78	282	79	283
rect	78	283	79	284
rect	78	284	79	285
rect	78	285	79	286
rect	78	286	79	287
rect	78	287	79	288
rect	78	288	79	289
rect	78	289	79	290
rect	78	290	79	291
rect	79	0	80	1
rect	79	1	80	2
rect	79	2	80	3
rect	79	3	80	4
rect	79	4	80	5
rect	79	5	80	6
rect	79	6	80	7
rect	79	7	80	8
rect	79	8	80	9
rect	79	9	80	10
rect	79	10	80	11
rect	79	11	80	12
rect	79	12	80	13
rect	79	13	80	14
rect	79	14	80	15
rect	79	15	80	16
rect	79	16	80	17
rect	79	17	80	18
rect	79	18	80	19
rect	79	19	80	20
rect	79	20	80	21
rect	79	21	80	22
rect	79	22	80	23
rect	79	23	80	24
rect	79	24	80	25
rect	79	25	80	26
rect	79	26	80	27
rect	79	27	80	28
rect	79	28	80	29
rect	79	29	80	30
rect	79	30	80	31
rect	79	31	80	32
rect	79	32	80	33
rect	79	33	80	34
rect	79	34	80	35
rect	79	35	80	36
rect	79	36	80	37
rect	79	37	80	38
rect	79	38	80	39
rect	79	39	80	40
rect	79	40	80	41
rect	79	41	80	42
rect	79	42	80	43
rect	79	43	80	44
rect	79	44	80	45
rect	79	45	80	46
rect	79	46	80	47
rect	79	47	80	48
rect	79	48	80	49
rect	79	49	80	50
rect	79	50	80	51
rect	79	51	80	52
rect	79	52	80	53
rect	79	53	80	54
rect	79	54	80	55
rect	79	55	80	56
rect	79	56	80	57
rect	79	57	80	58
rect	79	58	80	59
rect	79	59	80	60
rect	79	60	80	61
rect	79	61	80	62
rect	79	62	80	63
rect	79	63	80	64
rect	79	64	80	65
rect	79	65	80	66
rect	79	66	80	67
rect	79	67	80	68
rect	79	68	80	69
rect	79	69	80	70
rect	79	70	80	71
rect	79	71	80	72
rect	79	72	80	73
rect	79	73	80	74
rect	79	74	80	75
rect	79	75	80	76
rect	79	76	80	77
rect	79	77	80	78
rect	79	78	80	79
rect	79	79	80	80
rect	79	80	80	81
rect	79	81	80	82
rect	79	82	80	83
rect	79	83	80	84
rect	79	84	80	85
rect	79	85	80	86
rect	79	86	80	87
rect	79	87	80	88
rect	79	88	80	89
rect	79	89	80	90
rect	79	90	80	91
rect	79	91	80	92
rect	79	92	80	93
rect	79	93	80	94
rect	79	94	80	95
rect	79	95	80	96
rect	79	96	80	97
rect	79	97	80	98
rect	79	98	80	99
rect	79	99	80	100
rect	79	100	80	101
rect	79	101	80	102
rect	79	102	80	103
rect	79	103	80	104
rect	79	104	80	105
rect	79	105	80	106
rect	79	106	80	107
rect	79	107	80	108
rect	79	108	80	109
rect	79	109	80	110
rect	79	110	80	111
rect	79	111	80	112
rect	79	112	80	113
rect	79	113	80	114
rect	79	114	80	115
rect	79	115	80	116
rect	79	116	80	117
rect	79	117	80	118
rect	79	118	80	119
rect	79	119	80	120
rect	79	120	80	121
rect	79	121	80	122
rect	79	122	80	123
rect	79	123	80	124
rect	79	124	80	125
rect	79	125	80	126
rect	79	126	80	127
rect	79	127	80	128
rect	79	128	80	129
rect	79	129	80	130
rect	79	130	80	131
rect	79	131	80	132
rect	79	132	80	133
rect	79	133	80	134
rect	79	134	80	135
rect	79	135	80	136
rect	79	136	80	137
rect	79	137	80	138
rect	79	138	80	139
rect	79	139	80	140
rect	79	140	80	141
rect	79	141	80	142
rect	79	142	80	143
rect	79	143	80	144
rect	79	144	80	145
rect	79	145	80	146
rect	79	146	80	147
rect	79	147	80	148
rect	79	148	80	149
rect	79	149	80	150
rect	79	150	80	151
rect	79	151	80	152
rect	79	152	80	153
rect	79	153	80	154
rect	79	154	80	155
rect	79	155	80	156
rect	79	156	80	157
rect	79	157	80	158
rect	79	158	80	159
rect	79	159	80	160
rect	79	160	80	161
rect	79	161	80	162
rect	79	162	80	163
rect	79	163	80	164
rect	79	164	80	165
rect	79	165	80	166
rect	79	166	80	167
rect	79	167	80	168
rect	79	168	80	169
rect	79	169	80	170
rect	79	170	80	171
rect	79	171	80	172
rect	79	172	80	173
rect	79	173	80	174
rect	79	174	80	175
rect	79	175	80	176
rect	79	176	80	177
rect	79	177	80	178
rect	79	178	80	179
rect	79	179	80	180
rect	79	180	80	181
rect	79	181	80	182
rect	79	182	80	183
rect	79	183	80	184
rect	79	184	80	185
rect	79	185	80	186
rect	79	186	80	187
rect	79	187	80	188
rect	79	188	80	189
rect	79	189	80	190
rect	79	190	80	191
rect	79	191	80	192
rect	79	192	80	193
rect	79	193	80	194
rect	79	194	80	195
rect	79	195	80	196
rect	79	196	80	197
rect	79	197	80	198
rect	79	198	80	199
rect	79	199	80	200
rect	79	200	80	201
rect	79	201	80	202
rect	79	202	80	203
rect	79	203	80	204
rect	79	204	80	205
rect	79	205	80	206
rect	79	206	80	207
rect	79	207	80	208
rect	79	208	80	209
rect	79	209	80	210
rect	79	210	80	211
rect	79	211	80	212
rect	79	212	80	213
rect	79	213	80	214
rect	79	214	80	215
rect	79	215	80	216
rect	79	216	80	217
rect	79	217	80	218
rect	79	218	80	219
rect	79	219	80	220
rect	79	220	80	221
rect	79	221	80	222
rect	79	222	80	223
rect	79	223	80	224
rect	79	224	80	225
rect	79	225	80	226
rect	79	226	80	227
rect	79	227	80	228
rect	79	228	80	229
rect	79	229	80	230
rect	79	230	80	231
rect	79	231	80	232
rect	79	232	80	233
rect	79	233	80	234
rect	79	234	80	235
rect	79	235	80	236
rect	79	236	80	237
rect	79	237	80	238
rect	79	238	80	239
rect	79	239	80	240
rect	79	240	80	241
rect	79	241	80	242
rect	79	242	80	243
rect	79	243	80	244
rect	79	244	80	245
rect	79	245	80	246
rect	79	246	80	247
rect	79	247	80	248
rect	79	248	80	249
rect	79	249	80	250
rect	79	250	80	251
rect	79	251	80	252
rect	79	252	80	253
rect	79	253	80	254
rect	79	254	80	255
rect	79	255	80	256
rect	79	256	80	257
rect	79	257	80	258
rect	79	258	80	259
rect	79	259	80	260
rect	79	260	80	261
rect	79	261	80	262
rect	79	262	80	263
rect	79	263	80	264
rect	79	264	80	265
rect	79	265	80	266
rect	79	266	80	267
rect	79	267	80	268
rect	79	268	80	269
rect	79	269	80	270
rect	79	270	80	271
rect	79	271	80	272
rect	79	272	80	273
rect	79	273	80	274
rect	79	274	80	275
rect	79	275	80	276
rect	79	276	80	277
rect	79	277	80	278
rect	79	278	80	279
rect	79	279	80	280
rect	79	280	80	281
rect	79	281	80	282
rect	79	282	80	283
rect	79	283	80	284
rect	79	284	80	285
rect	79	285	80	286
rect	79	286	80	287
rect	79	287	80	288
rect	79	288	80	289
rect	79	289	80	290
rect	79	290	80	291
rect	80	0	81	1
rect	80	1	81	2
rect	80	2	81	3
rect	80	3	81	4
rect	80	4	81	5
rect	80	5	81	6
rect	80	6	81	7
rect	80	7	81	8
rect	80	8	81	9
rect	80	9	81	10
rect	80	10	81	11
rect	80	11	81	12
rect	80	12	81	13
rect	80	13	81	14
rect	80	14	81	15
rect	80	15	81	16
rect	80	16	81	17
rect	80	17	81	18
rect	80	18	81	19
rect	80	19	81	20
rect	80	20	81	21
rect	80	21	81	22
rect	80	22	81	23
rect	80	23	81	24
rect	80	24	81	25
rect	80	25	81	26
rect	80	26	81	27
rect	80	27	81	28
rect	80	28	81	29
rect	80	29	81	30
rect	80	30	81	31
rect	80	31	81	32
rect	80	32	81	33
rect	80	33	81	34
rect	80	34	81	35
rect	80	35	81	36
rect	80	36	81	37
rect	80	37	81	38
rect	80	38	81	39
rect	80	39	81	40
rect	80	40	81	41
rect	80	41	81	42
rect	80	42	81	43
rect	80	43	81	44
rect	80	44	81	45
rect	80	45	81	46
rect	80	46	81	47
rect	80	47	81	48
rect	80	48	81	49
rect	80	49	81	50
rect	80	50	81	51
rect	80	51	81	52
rect	80	52	81	53
rect	80	53	81	54
rect	80	54	81	55
rect	80	55	81	56
rect	80	56	81	57
rect	80	57	81	58
rect	80	58	81	59
rect	80	59	81	60
rect	80	60	81	61
rect	80	61	81	62
rect	80	62	81	63
rect	80	63	81	64
rect	80	64	81	65
rect	80	65	81	66
rect	80	66	81	67
rect	80	67	81	68
rect	80	68	81	69
rect	80	69	81	70
rect	80	70	81	71
rect	80	71	81	72
rect	80	72	81	73
rect	80	73	81	74
rect	80	74	81	75
rect	80	75	81	76
rect	80	76	81	77
rect	80	77	81	78
rect	80	78	81	79
rect	80	79	81	80
rect	80	80	81	81
rect	80	81	81	82
rect	80	82	81	83
rect	80	83	81	84
rect	80	84	81	85
rect	80	85	81	86
rect	80	86	81	87
rect	80	87	81	88
rect	80	88	81	89
rect	80	89	81	90
rect	80	90	81	91
rect	80	91	81	92
rect	80	92	81	93
rect	80	93	81	94
rect	80	94	81	95
rect	80	95	81	96
rect	80	96	81	97
rect	80	97	81	98
rect	80	98	81	99
rect	80	99	81	100
rect	80	100	81	101
rect	80	101	81	102
rect	80	102	81	103
rect	80	103	81	104
rect	80	104	81	105
rect	80	105	81	106
rect	80	106	81	107
rect	80	107	81	108
rect	80	108	81	109
rect	80	109	81	110
rect	80	110	81	111
rect	80	111	81	112
rect	80	112	81	113
rect	80	113	81	114
rect	80	114	81	115
rect	80	115	81	116
rect	80	116	81	117
rect	80	117	81	118
rect	80	118	81	119
rect	80	119	81	120
rect	80	120	81	121
rect	80	121	81	122
rect	80	122	81	123
rect	80	123	81	124
rect	80	124	81	125
rect	80	125	81	126
rect	80	126	81	127
rect	80	127	81	128
rect	80	128	81	129
rect	80	129	81	130
rect	80	130	81	131
rect	80	131	81	132
rect	80	132	81	133
rect	80	133	81	134
rect	80	134	81	135
rect	80	135	81	136
rect	80	136	81	137
rect	80	137	81	138
rect	80	138	81	139
rect	80	139	81	140
rect	80	140	81	141
rect	80	141	81	142
rect	80	142	81	143
rect	80	143	81	144
rect	80	144	81	145
rect	80	145	81	146
rect	80	146	81	147
rect	80	147	81	148
rect	80	148	81	149
rect	80	149	81	150
rect	80	150	81	151
rect	80	151	81	152
rect	80	152	81	153
rect	80	153	81	154
rect	80	154	81	155
rect	80	155	81	156
rect	80	156	81	157
rect	80	157	81	158
rect	80	158	81	159
rect	80	159	81	160
rect	80	160	81	161
rect	80	161	81	162
rect	80	162	81	163
rect	80	163	81	164
rect	80	164	81	165
rect	80	165	81	166
rect	80	166	81	167
rect	80	167	81	168
rect	80	168	81	169
rect	80	169	81	170
rect	80	170	81	171
rect	80	171	81	172
rect	80	172	81	173
rect	80	173	81	174
rect	80	174	81	175
rect	80	175	81	176
rect	80	176	81	177
rect	80	177	81	178
rect	80	178	81	179
rect	80	179	81	180
rect	80	180	81	181
rect	80	181	81	182
rect	80	182	81	183
rect	80	183	81	184
rect	80	184	81	185
rect	80	185	81	186
rect	80	186	81	187
rect	80	187	81	188
rect	80	188	81	189
rect	80	189	81	190
rect	80	190	81	191
rect	80	191	81	192
rect	80	192	81	193
rect	80	193	81	194
rect	80	194	81	195
rect	80	195	81	196
rect	80	196	81	197
rect	80	197	81	198
rect	80	198	81	199
rect	80	199	81	200
rect	80	200	81	201
rect	80	201	81	202
rect	80	202	81	203
rect	80	203	81	204
rect	80	204	81	205
rect	80	205	81	206
rect	80	206	81	207
rect	80	207	81	208
rect	80	208	81	209
rect	80	209	81	210
rect	80	210	81	211
rect	80	211	81	212
rect	80	212	81	213
rect	80	213	81	214
rect	80	214	81	215
rect	80	215	81	216
rect	80	216	81	217
rect	80	217	81	218
rect	80	218	81	219
rect	80	219	81	220
rect	80	220	81	221
rect	80	221	81	222
rect	80	222	81	223
rect	80	223	81	224
rect	80	224	81	225
rect	80	225	81	226
rect	80	226	81	227
rect	80	227	81	228
rect	80	228	81	229
rect	80	229	81	230
rect	80	230	81	231
rect	80	231	81	232
rect	80	232	81	233
rect	80	233	81	234
rect	80	234	81	235
rect	80	235	81	236
rect	80	236	81	237
rect	80	237	81	238
rect	80	238	81	239
rect	80	239	81	240
rect	80	240	81	241
rect	80	241	81	242
rect	80	242	81	243
rect	80	243	81	244
rect	80	244	81	245
rect	80	245	81	246
rect	80	246	81	247
rect	80	247	81	248
rect	80	248	81	249
rect	80	249	81	250
rect	80	250	81	251
rect	80	251	81	252
rect	80	252	81	253
rect	80	253	81	254
rect	80	254	81	255
rect	80	255	81	256
rect	80	256	81	257
rect	80	257	81	258
rect	80	258	81	259
rect	80	259	81	260
rect	80	260	81	261
rect	80	261	81	262
rect	80	262	81	263
rect	80	263	81	264
rect	80	264	81	265
rect	80	265	81	266
rect	80	266	81	267
rect	80	267	81	268
rect	80	268	81	269
rect	80	269	81	270
rect	80	270	81	271
rect	80	271	81	272
rect	80	272	81	273
rect	80	273	81	274
rect	80	274	81	275
rect	80	275	81	276
rect	80	276	81	277
rect	80	277	81	278
rect	80	278	81	279
rect	80	279	81	280
rect	80	280	81	281
rect	80	281	81	282
rect	80	282	81	283
rect	80	283	81	284
rect	80	284	81	285
rect	80	285	81	286
rect	80	286	81	287
rect	80	287	81	288
rect	80	288	81	289
rect	80	289	81	290
rect	80	290	81	291
rect	100	0	101	1
rect	100	1	101	2
rect	100	2	101	3
rect	100	3	101	4
rect	100	4	101	5
rect	100	5	101	6
rect	100	6	101	7
rect	100	7	101	8
rect	100	8	101	9
rect	100	9	101	10
rect	100	10	101	11
rect	100	11	101	12
rect	100	12	101	13
rect	100	13	101	14
rect	100	14	101	15
rect	100	15	101	16
rect	100	16	101	17
rect	100	17	101	18
rect	100	18	101	19
rect	100	19	101	20
rect	100	20	101	21
rect	100	21	101	22
rect	100	22	101	23
rect	100	23	101	24
rect	100	24	101	25
rect	100	25	101	26
rect	100	26	101	27
rect	100	27	101	28
rect	100	28	101	29
rect	100	29	101	30
rect	100	30	101	31
rect	100	31	101	32
rect	100	32	101	33
rect	100	33	101	34
rect	100	34	101	35
rect	100	35	101	36
rect	100	36	101	37
rect	100	37	101	38
rect	100	38	101	39
rect	100	39	101	40
rect	100	40	101	41
rect	100	41	101	42
rect	100	42	101	43
rect	100	43	101	44
rect	100	44	101	45
rect	100	45	101	46
rect	100	46	101	47
rect	100	47	101	48
rect	100	48	101	49
rect	100	49	101	50
rect	100	50	101	51
rect	100	51	101	52
rect	100	52	101	53
rect	100	53	101	54
rect	100	54	101	55
rect	100	55	101	56
rect	100	56	101	57
rect	100	57	101	58
rect	100	58	101	59
rect	100	59	101	60
rect	100	60	101	61
rect	100	61	101	62
rect	100	62	101	63
rect	100	63	101	64
rect	100	64	101	65
rect	100	65	101	66
rect	100	66	101	67
rect	100	67	101	68
rect	100	68	101	69
rect	100	69	101	70
rect	100	70	101	71
rect	100	71	101	72
rect	100	72	101	73
rect	100	73	101	74
rect	100	74	101	75
rect	100	75	101	76
rect	100	76	101	77
rect	100	77	101	78
rect	100	78	101	79
rect	100	79	101	80
rect	100	80	101	81
rect	100	81	101	82
rect	100	82	101	83
rect	100	83	101	84
rect	100	84	101	85
rect	100	85	101	86
rect	100	86	101	87
rect	100	87	101	88
rect	100	88	101	89
rect	100	89	101	90
rect	100	90	101	91
rect	100	91	101	92
rect	100	92	101	93
rect	100	93	101	94
rect	100	94	101	95
rect	100	95	101	96
rect	100	96	101	97
rect	100	97	101	98
rect	100	98	101	99
rect	100	99	101	100
rect	100	100	101	101
rect	100	101	101	102
rect	100	102	101	103
rect	100	103	101	104
rect	100	104	101	105
rect	100	105	101	106
rect	100	106	101	107
rect	100	107	101	108
rect	100	108	101	109
rect	100	109	101	110
rect	100	110	101	111
rect	100	111	101	112
rect	100	112	101	113
rect	100	113	101	114
rect	100	114	101	115
rect	100	115	101	116
rect	100	116	101	117
rect	100	117	101	118
rect	100	118	101	119
rect	100	119	101	120
rect	100	120	101	121
rect	100	121	101	122
rect	100	122	101	123
rect	100	123	101	124
rect	100	124	101	125
rect	100	125	101	126
rect	100	126	101	127
rect	100	127	101	128
rect	100	128	101	129
rect	100	129	101	130
rect	100	130	101	131
rect	100	131	101	132
rect	100	132	101	133
rect	100	133	101	134
rect	100	134	101	135
rect	100	135	101	136
rect	100	136	101	137
rect	100	137	101	138
rect	100	138	101	139
rect	100	139	101	140
rect	100	140	101	141
rect	100	141	101	142
rect	100	142	101	143
rect	100	143	101	144
rect	100	144	101	145
rect	100	145	101	146
rect	100	146	101	147
rect	100	147	101	148
rect	100	148	101	149
rect	100	149	101	150
rect	100	150	101	151
rect	100	151	101	152
rect	100	152	101	153
rect	100	153	101	154
rect	100	154	101	155
rect	100	155	101	156
rect	100	156	101	157
rect	100	157	101	158
rect	100	158	101	159
rect	100	159	101	160
rect	100	160	101	161
rect	100	161	101	162
rect	100	162	101	163
rect	100	163	101	164
rect	100	164	101	165
rect	100	165	101	166
rect	100	166	101	167
rect	100	167	101	168
rect	100	168	101	169
rect	100	169	101	170
rect	100	170	101	171
rect	100	171	101	172
rect	100	172	101	173
rect	100	173	101	174
rect	100	174	101	175
rect	100	175	101	176
rect	100	176	101	177
rect	100	177	101	178
rect	100	178	101	179
rect	100	179	101	180
rect	100	180	101	181
rect	100	181	101	182
rect	100	182	101	183
rect	100	183	101	184
rect	100	184	101	185
rect	100	185	101	186
rect	100	186	101	187
rect	100	187	101	188
rect	100	188	101	189
rect	100	189	101	190
rect	100	190	101	191
rect	100	191	101	192
rect	100	192	101	193
rect	100	193	101	194
rect	100	194	101	195
rect	100	195	101	196
rect	100	196	101	197
rect	100	197	101	198
rect	100	198	101	199
rect	100	199	101	200
rect	100	200	101	201
rect	100	201	101	202
rect	100	202	101	203
rect	100	203	101	204
rect	100	204	101	205
rect	100	205	101	206
rect	100	206	101	207
rect	100	207	101	208
rect	100	208	101	209
rect	100	209	101	210
rect	100	210	101	211
rect	100	211	101	212
rect	100	212	101	213
rect	100	213	101	214
rect	100	214	101	215
rect	100	215	101	216
rect	100	216	101	217
rect	100	217	101	218
rect	100	218	101	219
rect	100	219	101	220
rect	100	220	101	221
rect	100	221	101	222
rect	100	222	101	223
rect	100	223	101	224
rect	100	224	101	225
rect	100	225	101	226
rect	100	226	101	227
rect	100	227	101	228
rect	100	228	101	229
rect	100	229	101	230
rect	100	230	101	231
rect	100	231	101	232
rect	100	232	101	233
rect	100	233	101	234
rect	100	234	101	235
rect	100	235	101	236
rect	100	236	101	237
rect	100	237	101	238
rect	100	238	101	239
rect	100	239	101	240
rect	100	240	101	241
rect	100	241	101	242
rect	100	242	101	243
rect	100	243	101	244
rect	100	244	101	245
rect	100	245	101	246
rect	100	246	101	247
rect	100	247	101	248
rect	100	248	101	249
rect	100	249	101	250
rect	100	250	101	251
rect	100	251	101	252
rect	100	252	101	253
rect	100	253	101	254
rect	100	254	101	255
rect	100	255	101	256
rect	100	256	101	257
rect	100	257	101	258
rect	100	258	101	259
rect	100	259	101	260
rect	100	260	101	261
rect	100	261	101	262
rect	100	262	101	263
rect	100	263	101	264
rect	100	264	101	265
rect	100	265	101	266
rect	100	266	101	267
rect	100	267	101	268
rect	100	268	101	269
rect	100	269	101	270
rect	100	270	101	271
rect	100	271	101	272
rect	100	272	101	273
rect	100	273	101	274
rect	100	274	101	275
rect	100	275	101	276
rect	100	276	101	277
rect	100	277	101	278
rect	100	278	101	279
rect	100	279	101	280
rect	100	280	101	281
rect	100	281	101	282
rect	100	282	101	283
rect	100	283	101	284
rect	100	284	101	285
rect	100	285	101	286
rect	100	286	101	287
rect	100	287	101	288
rect	100	288	101	289
rect	100	289	101	290
rect	100	290	101	291
rect	100	291	101	292
rect	100	292	101	293
rect	100	293	101	294
rect	100	294	101	295
rect	100	295	101	296
rect	100	296	101	297
rect	100	297	101	298
rect	100	298	101	299
rect	100	299	101	300
rect	100	300	101	301
rect	100	301	101	302
rect	100	302	101	303
rect	100	303	101	304
rect	100	304	101	305
rect	100	305	101	306
rect	100	306	101	307
rect	100	307	101	308
rect	100	308	101	309
rect	100	309	101	310
rect	100	310	101	311
rect	100	311	101	312
rect	101	0	102	1
rect	101	1	102	2
rect	101	2	102	3
rect	101	3	102	4
rect	101	4	102	5
rect	101	5	102	6
rect	101	6	102	7
rect	101	7	102	8
rect	101	8	102	9
rect	101	9	102	10
rect	101	10	102	11
rect	101	11	102	12
rect	101	12	102	13
rect	101	13	102	14
rect	101	14	102	15
rect	101	15	102	16
rect	101	16	102	17
rect	101	17	102	18
rect	101	18	102	19
rect	101	19	102	20
rect	101	20	102	21
rect	101	21	102	22
rect	101	22	102	23
rect	101	23	102	24
rect	101	24	102	25
rect	101	25	102	26
rect	101	26	102	27
rect	101	27	102	28
rect	101	28	102	29
rect	101	29	102	30
rect	101	30	102	31
rect	101	31	102	32
rect	101	32	102	33
rect	101	33	102	34
rect	101	34	102	35
rect	101	35	102	36
rect	101	36	102	37
rect	101	37	102	38
rect	101	38	102	39
rect	101	39	102	40
rect	101	40	102	41
rect	101	41	102	42
rect	101	42	102	43
rect	101	43	102	44
rect	101	44	102	45
rect	101	45	102	46
rect	101	46	102	47
rect	101	47	102	48
rect	101	48	102	49
rect	101	49	102	50
rect	101	50	102	51
rect	101	51	102	52
rect	101	52	102	53
rect	101	53	102	54
rect	101	54	102	55
rect	101	55	102	56
rect	101	56	102	57
rect	101	57	102	58
rect	101	58	102	59
rect	101	59	102	60
rect	101	60	102	61
rect	101	61	102	62
rect	101	62	102	63
rect	101	63	102	64
rect	101	64	102	65
rect	101	65	102	66
rect	101	66	102	67
rect	101	67	102	68
rect	101	68	102	69
rect	101	69	102	70
rect	101	70	102	71
rect	101	71	102	72
rect	101	72	102	73
rect	101	73	102	74
rect	101	74	102	75
rect	101	75	102	76
rect	101	76	102	77
rect	101	77	102	78
rect	101	78	102	79
rect	101	79	102	80
rect	101	80	102	81
rect	101	81	102	82
rect	101	82	102	83
rect	101	83	102	84
rect	101	84	102	85
rect	101	85	102	86
rect	101	86	102	87
rect	101	87	102	88
rect	101	88	102	89
rect	101	89	102	90
rect	101	90	102	91
rect	101	91	102	92
rect	101	92	102	93
rect	101	93	102	94
rect	101	94	102	95
rect	101	95	102	96
rect	101	96	102	97
rect	101	97	102	98
rect	101	98	102	99
rect	101	99	102	100
rect	101	100	102	101
rect	101	101	102	102
rect	101	102	102	103
rect	101	103	102	104
rect	101	104	102	105
rect	101	105	102	106
rect	101	106	102	107
rect	101	107	102	108
rect	101	108	102	109
rect	101	109	102	110
rect	101	110	102	111
rect	101	111	102	112
rect	101	112	102	113
rect	101	113	102	114
rect	101	114	102	115
rect	101	115	102	116
rect	101	116	102	117
rect	101	117	102	118
rect	101	118	102	119
rect	101	119	102	120
rect	101	120	102	121
rect	101	121	102	122
rect	101	122	102	123
rect	101	123	102	124
rect	101	124	102	125
rect	101	125	102	126
rect	101	126	102	127
rect	101	127	102	128
rect	101	128	102	129
rect	101	129	102	130
rect	101	130	102	131
rect	101	131	102	132
rect	101	132	102	133
rect	101	133	102	134
rect	101	134	102	135
rect	101	135	102	136
rect	101	136	102	137
rect	101	137	102	138
rect	101	138	102	139
rect	101	139	102	140
rect	101	140	102	141
rect	101	141	102	142
rect	101	142	102	143
rect	101	143	102	144
rect	101	144	102	145
rect	101	145	102	146
rect	101	146	102	147
rect	101	147	102	148
rect	101	148	102	149
rect	101	149	102	150
rect	101	150	102	151
rect	101	151	102	152
rect	101	152	102	153
rect	101	153	102	154
rect	101	154	102	155
rect	101	155	102	156
rect	101	156	102	157
rect	101	157	102	158
rect	101	158	102	159
rect	101	159	102	160
rect	101	160	102	161
rect	101	161	102	162
rect	101	162	102	163
rect	101	163	102	164
rect	101	164	102	165
rect	101	165	102	166
rect	101	166	102	167
rect	101	167	102	168
rect	101	168	102	169
rect	101	169	102	170
rect	101	170	102	171
rect	101	171	102	172
rect	101	172	102	173
rect	101	173	102	174
rect	101	174	102	175
rect	101	175	102	176
rect	101	176	102	177
rect	101	177	102	178
rect	101	178	102	179
rect	101	179	102	180
rect	101	180	102	181
rect	101	181	102	182
rect	101	182	102	183
rect	101	183	102	184
rect	101	184	102	185
rect	101	185	102	186
rect	101	186	102	187
rect	101	187	102	188
rect	101	188	102	189
rect	101	189	102	190
rect	101	190	102	191
rect	101	191	102	192
rect	101	192	102	193
rect	101	193	102	194
rect	101	194	102	195
rect	101	195	102	196
rect	101	196	102	197
rect	101	197	102	198
rect	101	198	102	199
rect	101	199	102	200
rect	101	200	102	201
rect	101	201	102	202
rect	101	202	102	203
rect	101	203	102	204
rect	101	204	102	205
rect	101	205	102	206
rect	101	206	102	207
rect	101	207	102	208
rect	101	208	102	209
rect	101	209	102	210
rect	101	210	102	211
rect	101	211	102	212
rect	101	212	102	213
rect	101	213	102	214
rect	101	214	102	215
rect	101	215	102	216
rect	101	216	102	217
rect	101	217	102	218
rect	101	218	102	219
rect	101	219	102	220
rect	101	220	102	221
rect	101	221	102	222
rect	101	222	102	223
rect	101	223	102	224
rect	101	224	102	225
rect	101	225	102	226
rect	101	226	102	227
rect	101	227	102	228
rect	101	228	102	229
rect	101	229	102	230
rect	101	230	102	231
rect	101	231	102	232
rect	101	232	102	233
rect	101	233	102	234
rect	101	234	102	235
rect	101	235	102	236
rect	101	236	102	237
rect	101	237	102	238
rect	101	238	102	239
rect	101	239	102	240
rect	101	240	102	241
rect	101	241	102	242
rect	101	242	102	243
rect	101	243	102	244
rect	101	244	102	245
rect	101	245	102	246
rect	101	246	102	247
rect	101	247	102	248
rect	101	248	102	249
rect	101	249	102	250
rect	101	250	102	251
rect	101	251	102	252
rect	101	252	102	253
rect	101	253	102	254
rect	101	254	102	255
rect	101	255	102	256
rect	101	256	102	257
rect	101	257	102	258
rect	101	258	102	259
rect	101	259	102	260
rect	101	260	102	261
rect	101	261	102	262
rect	101	262	102	263
rect	101	263	102	264
rect	101	264	102	265
rect	101	265	102	266
rect	101	266	102	267
rect	101	267	102	268
rect	101	268	102	269
rect	101	269	102	270
rect	101	270	102	271
rect	101	271	102	272
rect	101	272	102	273
rect	101	273	102	274
rect	101	274	102	275
rect	101	275	102	276
rect	101	276	102	277
rect	101	277	102	278
rect	101	278	102	279
rect	101	279	102	280
rect	101	280	102	281
rect	101	281	102	282
rect	101	282	102	283
rect	101	283	102	284
rect	101	284	102	285
rect	101	285	102	286
rect	101	286	102	287
rect	101	287	102	288
rect	101	288	102	289
rect	101	289	102	290
rect	101	290	102	291
rect	101	291	102	292
rect	101	292	102	293
rect	101	293	102	294
rect	101	294	102	295
rect	101	295	102	296
rect	101	296	102	297
rect	101	297	102	298
rect	101	298	102	299
rect	101	299	102	300
rect	101	300	102	301
rect	101	301	102	302
rect	101	302	102	303
rect	101	303	102	304
rect	101	304	102	305
rect	101	305	102	306
rect	101	306	102	307
rect	101	307	102	308
rect	101	308	102	309
rect	101	309	102	310
rect	101	310	102	311
rect	101	311	102	312
rect	102	0	103	1
rect	102	1	103	2
rect	102	2	103	3
rect	102	3	103	4
rect	102	4	103	5
rect	102	5	103	6
rect	102	6	103	7
rect	102	7	103	8
rect	102	8	103	9
rect	102	9	103	10
rect	102	10	103	11
rect	102	11	103	12
rect	102	12	103	13
rect	102	13	103	14
rect	102	14	103	15
rect	102	15	103	16
rect	102	16	103	17
rect	102	17	103	18
rect	102	18	103	19
rect	102	19	103	20
rect	102	20	103	21
rect	102	21	103	22
rect	102	22	103	23
rect	102	23	103	24
rect	102	24	103	25
rect	102	25	103	26
rect	102	26	103	27
rect	102	27	103	28
rect	102	28	103	29
rect	102	29	103	30
rect	102	30	103	31
rect	102	31	103	32
rect	102	32	103	33
rect	102	33	103	34
rect	102	34	103	35
rect	102	35	103	36
rect	102	36	103	37
rect	102	37	103	38
rect	102	38	103	39
rect	102	39	103	40
rect	102	40	103	41
rect	102	41	103	42
rect	102	42	103	43
rect	102	43	103	44
rect	102	44	103	45
rect	102	45	103	46
rect	102	46	103	47
rect	102	47	103	48
rect	102	48	103	49
rect	102	49	103	50
rect	102	50	103	51
rect	102	51	103	52
rect	102	52	103	53
rect	102	53	103	54
rect	102	54	103	55
rect	102	55	103	56
rect	102	56	103	57
rect	102	57	103	58
rect	102	58	103	59
rect	102	59	103	60
rect	102	60	103	61
rect	102	61	103	62
rect	102	62	103	63
rect	102	63	103	64
rect	102	64	103	65
rect	102	65	103	66
rect	102	66	103	67
rect	102	67	103	68
rect	102	68	103	69
rect	102	69	103	70
rect	102	70	103	71
rect	102	71	103	72
rect	102	72	103	73
rect	102	73	103	74
rect	102	74	103	75
rect	102	75	103	76
rect	102	76	103	77
rect	102	77	103	78
rect	102	78	103	79
rect	102	79	103	80
rect	102	80	103	81
rect	102	81	103	82
rect	102	82	103	83
rect	102	83	103	84
rect	102	84	103	85
rect	102	85	103	86
rect	102	86	103	87
rect	102	87	103	88
rect	102	88	103	89
rect	102	89	103	90
rect	102	90	103	91
rect	102	91	103	92
rect	102	92	103	93
rect	102	93	103	94
rect	102	94	103	95
rect	102	95	103	96
rect	102	96	103	97
rect	102	97	103	98
rect	102	98	103	99
rect	102	99	103	100
rect	102	100	103	101
rect	102	101	103	102
rect	102	102	103	103
rect	102	103	103	104
rect	102	104	103	105
rect	102	105	103	106
rect	102	106	103	107
rect	102	107	103	108
rect	102	108	103	109
rect	102	109	103	110
rect	102	110	103	111
rect	102	111	103	112
rect	102	112	103	113
rect	102	113	103	114
rect	102	114	103	115
rect	102	115	103	116
rect	102	116	103	117
rect	102	117	103	118
rect	102	118	103	119
rect	102	119	103	120
rect	102	120	103	121
rect	102	121	103	122
rect	102	122	103	123
rect	102	123	103	124
rect	102	124	103	125
rect	102	125	103	126
rect	102	126	103	127
rect	102	127	103	128
rect	102	128	103	129
rect	102	129	103	130
rect	102	130	103	131
rect	102	131	103	132
rect	102	132	103	133
rect	102	133	103	134
rect	102	134	103	135
rect	102	135	103	136
rect	102	136	103	137
rect	102	137	103	138
rect	102	138	103	139
rect	102	139	103	140
rect	102	140	103	141
rect	102	141	103	142
rect	102	142	103	143
rect	102	143	103	144
rect	102	144	103	145
rect	102	145	103	146
rect	102	146	103	147
rect	102	147	103	148
rect	102	148	103	149
rect	102	149	103	150
rect	102	150	103	151
rect	102	151	103	152
rect	102	152	103	153
rect	102	153	103	154
rect	102	154	103	155
rect	102	155	103	156
rect	102	156	103	157
rect	102	157	103	158
rect	102	158	103	159
rect	102	159	103	160
rect	102	160	103	161
rect	102	161	103	162
rect	102	162	103	163
rect	102	163	103	164
rect	102	164	103	165
rect	102	165	103	166
rect	102	166	103	167
rect	102	167	103	168
rect	102	168	103	169
rect	102	169	103	170
rect	102	170	103	171
rect	102	171	103	172
rect	102	172	103	173
rect	102	173	103	174
rect	102	174	103	175
rect	102	175	103	176
rect	102	176	103	177
rect	102	177	103	178
rect	102	178	103	179
rect	102	179	103	180
rect	102	180	103	181
rect	102	181	103	182
rect	102	182	103	183
rect	102	183	103	184
rect	102	184	103	185
rect	102	185	103	186
rect	102	186	103	187
rect	102	187	103	188
rect	102	188	103	189
rect	102	189	103	190
rect	102	190	103	191
rect	102	191	103	192
rect	102	192	103	193
rect	102	193	103	194
rect	102	194	103	195
rect	102	195	103	196
rect	102	196	103	197
rect	102	197	103	198
rect	102	198	103	199
rect	102	199	103	200
rect	102	200	103	201
rect	102	201	103	202
rect	102	202	103	203
rect	102	203	103	204
rect	102	204	103	205
rect	102	205	103	206
rect	102	206	103	207
rect	102	207	103	208
rect	102	208	103	209
rect	102	209	103	210
rect	102	210	103	211
rect	102	211	103	212
rect	102	212	103	213
rect	102	213	103	214
rect	102	214	103	215
rect	102	215	103	216
rect	102	216	103	217
rect	102	217	103	218
rect	102	218	103	219
rect	102	219	103	220
rect	102	220	103	221
rect	102	221	103	222
rect	102	222	103	223
rect	102	223	103	224
rect	102	224	103	225
rect	102	225	103	226
rect	102	226	103	227
rect	102	227	103	228
rect	102	228	103	229
rect	102	229	103	230
rect	102	230	103	231
rect	102	231	103	232
rect	102	232	103	233
rect	102	233	103	234
rect	102	234	103	235
rect	102	235	103	236
rect	102	236	103	237
rect	102	237	103	238
rect	102	238	103	239
rect	102	239	103	240
rect	102	240	103	241
rect	102	241	103	242
rect	102	242	103	243
rect	102	243	103	244
rect	102	244	103	245
rect	102	245	103	246
rect	102	246	103	247
rect	102	247	103	248
rect	102	248	103	249
rect	102	249	103	250
rect	102	250	103	251
rect	102	251	103	252
rect	102	252	103	253
rect	102	253	103	254
rect	102	254	103	255
rect	102	255	103	256
rect	102	256	103	257
rect	102	257	103	258
rect	102	258	103	259
rect	102	259	103	260
rect	102	260	103	261
rect	102	261	103	262
rect	102	262	103	263
rect	102	263	103	264
rect	102	264	103	265
rect	102	265	103	266
rect	102	266	103	267
rect	102	267	103	268
rect	102	268	103	269
rect	102	269	103	270
rect	102	270	103	271
rect	102	271	103	272
rect	102	272	103	273
rect	102	273	103	274
rect	102	274	103	275
rect	102	275	103	276
rect	102	276	103	277
rect	102	277	103	278
rect	102	278	103	279
rect	102	279	103	280
rect	102	280	103	281
rect	102	281	103	282
rect	102	282	103	283
rect	102	283	103	284
rect	102	284	103	285
rect	102	285	103	286
rect	102	286	103	287
rect	102	287	103	288
rect	102	288	103	289
rect	102	289	103	290
rect	102	290	103	291
rect	102	291	103	292
rect	102	292	103	293
rect	102	293	103	294
rect	102	294	103	295
rect	102	295	103	296
rect	102	296	103	297
rect	102	297	103	298
rect	102	298	103	299
rect	102	299	103	300
rect	102	300	103	301
rect	102	301	103	302
rect	102	302	103	303
rect	102	303	103	304
rect	102	304	103	305
rect	102	305	103	306
rect	102	306	103	307
rect	102	307	103	308
rect	102	308	103	309
rect	102	309	103	310
rect	102	310	103	311
rect	102	311	103	312
rect	103	0	104	1
rect	103	1	104	2
rect	103	2	104	3
rect	103	3	104	4
rect	103	4	104	5
rect	103	5	104	6
rect	103	6	104	7
rect	103	7	104	8
rect	103	8	104	9
rect	103	9	104	10
rect	103	10	104	11
rect	103	11	104	12
rect	103	12	104	13
rect	103	13	104	14
rect	103	14	104	15
rect	103	15	104	16
rect	103	16	104	17
rect	103	17	104	18
rect	103	18	104	19
rect	103	19	104	20
rect	103	20	104	21
rect	103	21	104	22
rect	103	22	104	23
rect	103	23	104	24
rect	103	24	104	25
rect	103	25	104	26
rect	103	26	104	27
rect	103	27	104	28
rect	103	28	104	29
rect	103	29	104	30
rect	103	30	104	31
rect	103	31	104	32
rect	103	32	104	33
rect	103	33	104	34
rect	103	34	104	35
rect	103	35	104	36
rect	103	36	104	37
rect	103	37	104	38
rect	103	38	104	39
rect	103	39	104	40
rect	103	40	104	41
rect	103	41	104	42
rect	103	42	104	43
rect	103	43	104	44
rect	103	44	104	45
rect	103	45	104	46
rect	103	46	104	47
rect	103	47	104	48
rect	103	48	104	49
rect	103	49	104	50
rect	103	50	104	51
rect	103	51	104	52
rect	103	52	104	53
rect	103	53	104	54
rect	103	54	104	55
rect	103	55	104	56
rect	103	56	104	57
rect	103	57	104	58
rect	103	58	104	59
rect	103	59	104	60
rect	103	60	104	61
rect	103	61	104	62
rect	103	62	104	63
rect	103	63	104	64
rect	103	64	104	65
rect	103	65	104	66
rect	103	66	104	67
rect	103	67	104	68
rect	103	68	104	69
rect	103	69	104	70
rect	103	70	104	71
rect	103	71	104	72
rect	103	72	104	73
rect	103	73	104	74
rect	103	74	104	75
rect	103	75	104	76
rect	103	76	104	77
rect	103	77	104	78
rect	103	78	104	79
rect	103	79	104	80
rect	103	80	104	81
rect	103	81	104	82
rect	103	82	104	83
rect	103	83	104	84
rect	103	84	104	85
rect	103	85	104	86
rect	103	86	104	87
rect	103	87	104	88
rect	103	88	104	89
rect	103	89	104	90
rect	103	90	104	91
rect	103	91	104	92
rect	103	92	104	93
rect	103	93	104	94
rect	103	94	104	95
rect	103	95	104	96
rect	103	96	104	97
rect	103	97	104	98
rect	103	98	104	99
rect	103	99	104	100
rect	103	100	104	101
rect	103	101	104	102
rect	103	102	104	103
rect	103	103	104	104
rect	103	104	104	105
rect	103	105	104	106
rect	103	106	104	107
rect	103	107	104	108
rect	103	108	104	109
rect	103	109	104	110
rect	103	110	104	111
rect	103	111	104	112
rect	103	112	104	113
rect	103	113	104	114
rect	103	114	104	115
rect	103	115	104	116
rect	103	116	104	117
rect	103	117	104	118
rect	103	118	104	119
rect	103	119	104	120
rect	103	120	104	121
rect	103	121	104	122
rect	103	122	104	123
rect	103	123	104	124
rect	103	124	104	125
rect	103	125	104	126
rect	103	126	104	127
rect	103	127	104	128
rect	103	128	104	129
rect	103	129	104	130
rect	103	130	104	131
rect	103	131	104	132
rect	103	132	104	133
rect	103	133	104	134
rect	103	134	104	135
rect	103	135	104	136
rect	103	136	104	137
rect	103	137	104	138
rect	103	138	104	139
rect	103	139	104	140
rect	103	140	104	141
rect	103	141	104	142
rect	103	142	104	143
rect	103	143	104	144
rect	103	144	104	145
rect	103	145	104	146
rect	103	146	104	147
rect	103	147	104	148
rect	103	148	104	149
rect	103	149	104	150
rect	103	150	104	151
rect	103	151	104	152
rect	103	152	104	153
rect	103	153	104	154
rect	103	154	104	155
rect	103	155	104	156
rect	103	156	104	157
rect	103	157	104	158
rect	103	158	104	159
rect	103	159	104	160
rect	103	160	104	161
rect	103	161	104	162
rect	103	162	104	163
rect	103	163	104	164
rect	103	164	104	165
rect	103	165	104	166
rect	103	166	104	167
rect	103	167	104	168
rect	103	168	104	169
rect	103	169	104	170
rect	103	170	104	171
rect	103	171	104	172
rect	103	172	104	173
rect	103	173	104	174
rect	103	174	104	175
rect	103	175	104	176
rect	103	176	104	177
rect	103	177	104	178
rect	103	178	104	179
rect	103	179	104	180
rect	103	180	104	181
rect	103	181	104	182
rect	103	182	104	183
rect	103	183	104	184
rect	103	184	104	185
rect	103	185	104	186
rect	103	186	104	187
rect	103	187	104	188
rect	103	188	104	189
rect	103	189	104	190
rect	103	190	104	191
rect	103	191	104	192
rect	103	192	104	193
rect	103	193	104	194
rect	103	194	104	195
rect	103	195	104	196
rect	103	196	104	197
rect	103	197	104	198
rect	103	198	104	199
rect	103	199	104	200
rect	103	200	104	201
rect	103	201	104	202
rect	103	202	104	203
rect	103	203	104	204
rect	103	204	104	205
rect	103	205	104	206
rect	103	206	104	207
rect	103	207	104	208
rect	103	208	104	209
rect	103	209	104	210
rect	103	210	104	211
rect	103	211	104	212
rect	103	212	104	213
rect	103	213	104	214
rect	103	214	104	215
rect	103	215	104	216
rect	103	216	104	217
rect	103	217	104	218
rect	103	218	104	219
rect	103	219	104	220
rect	103	220	104	221
rect	103	221	104	222
rect	103	222	104	223
rect	103	223	104	224
rect	103	224	104	225
rect	103	225	104	226
rect	103	226	104	227
rect	103	227	104	228
rect	103	228	104	229
rect	103	229	104	230
rect	103	230	104	231
rect	103	231	104	232
rect	103	232	104	233
rect	103	233	104	234
rect	103	234	104	235
rect	103	235	104	236
rect	103	236	104	237
rect	103	237	104	238
rect	103	238	104	239
rect	103	239	104	240
rect	103	240	104	241
rect	103	241	104	242
rect	103	242	104	243
rect	103	243	104	244
rect	103	244	104	245
rect	103	245	104	246
rect	103	246	104	247
rect	103	247	104	248
rect	103	248	104	249
rect	103	249	104	250
rect	103	250	104	251
rect	103	251	104	252
rect	103	252	104	253
rect	103	253	104	254
rect	103	254	104	255
rect	103	255	104	256
rect	103	256	104	257
rect	103	257	104	258
rect	103	258	104	259
rect	103	259	104	260
rect	103	260	104	261
rect	103	261	104	262
rect	103	262	104	263
rect	103	263	104	264
rect	103	264	104	265
rect	103	265	104	266
rect	103	266	104	267
rect	103	267	104	268
rect	103	268	104	269
rect	103	269	104	270
rect	103	270	104	271
rect	103	271	104	272
rect	103	272	104	273
rect	103	273	104	274
rect	103	274	104	275
rect	103	275	104	276
rect	103	276	104	277
rect	103	277	104	278
rect	103	278	104	279
rect	103	279	104	280
rect	103	280	104	281
rect	103	281	104	282
rect	103	282	104	283
rect	103	283	104	284
rect	103	284	104	285
rect	103	285	104	286
rect	103	286	104	287
rect	103	287	104	288
rect	103	288	104	289
rect	103	289	104	290
rect	103	290	104	291
rect	103	291	104	292
rect	103	292	104	293
rect	103	293	104	294
rect	103	294	104	295
rect	103	295	104	296
rect	103	296	104	297
rect	103	297	104	298
rect	103	298	104	299
rect	103	299	104	300
rect	103	300	104	301
rect	103	301	104	302
rect	103	302	104	303
rect	103	303	104	304
rect	103	304	104	305
rect	103	305	104	306
rect	103	306	104	307
rect	103	307	104	308
rect	103	308	104	309
rect	103	309	104	310
rect	103	310	104	311
rect	103	311	104	312
rect	104	0	105	1
rect	104	1	105	2
rect	104	2	105	3
rect	104	3	105	4
rect	104	4	105	5
rect	104	5	105	6
rect	104	6	105	7
rect	104	7	105	8
rect	104	8	105	9
rect	104	9	105	10
rect	104	10	105	11
rect	104	11	105	12
rect	104	12	105	13
rect	104	13	105	14
rect	104	14	105	15
rect	104	15	105	16
rect	104	16	105	17
rect	104	17	105	18
rect	104	18	105	19
rect	104	19	105	20
rect	104	20	105	21
rect	104	21	105	22
rect	104	22	105	23
rect	104	23	105	24
rect	104	24	105	25
rect	104	25	105	26
rect	104	26	105	27
rect	104	27	105	28
rect	104	28	105	29
rect	104	29	105	30
rect	104	30	105	31
rect	104	31	105	32
rect	104	32	105	33
rect	104	33	105	34
rect	104	34	105	35
rect	104	35	105	36
rect	104	36	105	37
rect	104	37	105	38
rect	104	38	105	39
rect	104	39	105	40
rect	104	40	105	41
rect	104	41	105	42
rect	104	42	105	43
rect	104	43	105	44
rect	104	44	105	45
rect	104	45	105	46
rect	104	46	105	47
rect	104	47	105	48
rect	104	48	105	49
rect	104	49	105	50
rect	104	50	105	51
rect	104	51	105	52
rect	104	52	105	53
rect	104	53	105	54
rect	104	54	105	55
rect	104	55	105	56
rect	104	56	105	57
rect	104	57	105	58
rect	104	58	105	59
rect	104	59	105	60
rect	104	60	105	61
rect	104	61	105	62
rect	104	62	105	63
rect	104	63	105	64
rect	104	64	105	65
rect	104	65	105	66
rect	104	66	105	67
rect	104	67	105	68
rect	104	68	105	69
rect	104	69	105	70
rect	104	70	105	71
rect	104	71	105	72
rect	104	72	105	73
rect	104	73	105	74
rect	104	74	105	75
rect	104	75	105	76
rect	104	76	105	77
rect	104	77	105	78
rect	104	78	105	79
rect	104	79	105	80
rect	104	80	105	81
rect	104	81	105	82
rect	104	82	105	83
rect	104	83	105	84
rect	104	84	105	85
rect	104	85	105	86
rect	104	86	105	87
rect	104	87	105	88
rect	104	88	105	89
rect	104	89	105	90
rect	104	90	105	91
rect	104	91	105	92
rect	104	92	105	93
rect	104	93	105	94
rect	104	94	105	95
rect	104	95	105	96
rect	104	96	105	97
rect	104	97	105	98
rect	104	98	105	99
rect	104	99	105	100
rect	104	100	105	101
rect	104	101	105	102
rect	104	102	105	103
rect	104	103	105	104
rect	104	104	105	105
rect	104	105	105	106
rect	104	106	105	107
rect	104	107	105	108
rect	104	108	105	109
rect	104	109	105	110
rect	104	110	105	111
rect	104	111	105	112
rect	104	112	105	113
rect	104	113	105	114
rect	104	114	105	115
rect	104	115	105	116
rect	104	116	105	117
rect	104	117	105	118
rect	104	118	105	119
rect	104	119	105	120
rect	104	120	105	121
rect	104	121	105	122
rect	104	122	105	123
rect	104	123	105	124
rect	104	124	105	125
rect	104	125	105	126
rect	104	126	105	127
rect	104	127	105	128
rect	104	128	105	129
rect	104	129	105	130
rect	104	130	105	131
rect	104	131	105	132
rect	104	132	105	133
rect	104	133	105	134
rect	104	134	105	135
rect	104	135	105	136
rect	104	136	105	137
rect	104	137	105	138
rect	104	138	105	139
rect	104	139	105	140
rect	104	140	105	141
rect	104	141	105	142
rect	104	142	105	143
rect	104	143	105	144
rect	104	144	105	145
rect	104	145	105	146
rect	104	146	105	147
rect	104	147	105	148
rect	104	148	105	149
rect	104	149	105	150
rect	104	150	105	151
rect	104	151	105	152
rect	104	152	105	153
rect	104	153	105	154
rect	104	154	105	155
rect	104	155	105	156
rect	104	156	105	157
rect	104	157	105	158
rect	104	158	105	159
rect	104	159	105	160
rect	104	160	105	161
rect	104	161	105	162
rect	104	162	105	163
rect	104	163	105	164
rect	104	164	105	165
rect	104	165	105	166
rect	104	166	105	167
rect	104	167	105	168
rect	104	168	105	169
rect	104	169	105	170
rect	104	170	105	171
rect	104	171	105	172
rect	104	172	105	173
rect	104	173	105	174
rect	104	174	105	175
rect	104	175	105	176
rect	104	176	105	177
rect	104	177	105	178
rect	104	178	105	179
rect	104	179	105	180
rect	104	180	105	181
rect	104	181	105	182
rect	104	182	105	183
rect	104	183	105	184
rect	104	184	105	185
rect	104	185	105	186
rect	104	186	105	187
rect	104	187	105	188
rect	104	188	105	189
rect	104	189	105	190
rect	104	190	105	191
rect	104	191	105	192
rect	104	192	105	193
rect	104	193	105	194
rect	104	194	105	195
rect	104	195	105	196
rect	104	196	105	197
rect	104	197	105	198
rect	104	198	105	199
rect	104	199	105	200
rect	104	200	105	201
rect	104	201	105	202
rect	104	202	105	203
rect	104	203	105	204
rect	104	204	105	205
rect	104	205	105	206
rect	104	206	105	207
rect	104	207	105	208
rect	104	208	105	209
rect	104	209	105	210
rect	104	210	105	211
rect	104	211	105	212
rect	104	212	105	213
rect	104	213	105	214
rect	104	214	105	215
rect	104	215	105	216
rect	104	216	105	217
rect	104	217	105	218
rect	104	218	105	219
rect	104	219	105	220
rect	104	220	105	221
rect	104	221	105	222
rect	104	222	105	223
rect	104	223	105	224
rect	104	224	105	225
rect	104	225	105	226
rect	104	226	105	227
rect	104	227	105	228
rect	104	228	105	229
rect	104	229	105	230
rect	104	230	105	231
rect	104	231	105	232
rect	104	232	105	233
rect	104	233	105	234
rect	104	234	105	235
rect	104	235	105	236
rect	104	236	105	237
rect	104	237	105	238
rect	104	238	105	239
rect	104	239	105	240
rect	104	240	105	241
rect	104	241	105	242
rect	104	242	105	243
rect	104	243	105	244
rect	104	244	105	245
rect	104	245	105	246
rect	104	246	105	247
rect	104	247	105	248
rect	104	248	105	249
rect	104	249	105	250
rect	104	250	105	251
rect	104	251	105	252
rect	104	252	105	253
rect	104	253	105	254
rect	104	254	105	255
rect	104	255	105	256
rect	104	256	105	257
rect	104	257	105	258
rect	104	258	105	259
rect	104	259	105	260
rect	104	260	105	261
rect	104	261	105	262
rect	104	262	105	263
rect	104	263	105	264
rect	104	264	105	265
rect	104	265	105	266
rect	104	266	105	267
rect	104	267	105	268
rect	104	268	105	269
rect	104	269	105	270
rect	104	270	105	271
rect	104	271	105	272
rect	104	272	105	273
rect	104	273	105	274
rect	104	274	105	275
rect	104	275	105	276
rect	104	276	105	277
rect	104	277	105	278
rect	104	278	105	279
rect	104	279	105	280
rect	104	280	105	281
rect	104	281	105	282
rect	104	282	105	283
rect	104	283	105	284
rect	104	284	105	285
rect	104	285	105	286
rect	104	286	105	287
rect	104	287	105	288
rect	104	288	105	289
rect	104	289	105	290
rect	104	290	105	291
rect	104	291	105	292
rect	104	292	105	293
rect	104	293	105	294
rect	104	294	105	295
rect	104	295	105	296
rect	104	296	105	297
rect	104	297	105	298
rect	104	298	105	299
rect	104	299	105	300
rect	104	300	105	301
rect	104	301	105	302
rect	104	302	105	303
rect	104	303	105	304
rect	104	304	105	305
rect	104	305	105	306
rect	104	306	105	307
rect	104	307	105	308
rect	104	308	105	309
rect	104	309	105	310
rect	104	310	105	311
rect	104	311	105	312
rect	105	0	106	1
rect	105	1	106	2
rect	105	2	106	3
rect	105	3	106	4
rect	105	4	106	5
rect	105	5	106	6
rect	105	6	106	7
rect	105	7	106	8
rect	105	8	106	9
rect	105	9	106	10
rect	105	10	106	11
rect	105	11	106	12
rect	105	12	106	13
rect	105	13	106	14
rect	105	14	106	15
rect	105	15	106	16
rect	105	16	106	17
rect	105	17	106	18
rect	105	18	106	19
rect	105	19	106	20
rect	105	20	106	21
rect	105	21	106	22
rect	105	22	106	23
rect	105	23	106	24
rect	105	24	106	25
rect	105	25	106	26
rect	105	26	106	27
rect	105	27	106	28
rect	105	28	106	29
rect	105	29	106	30
rect	105	30	106	31
rect	105	31	106	32
rect	105	32	106	33
rect	105	33	106	34
rect	105	34	106	35
rect	105	35	106	36
rect	105	36	106	37
rect	105	37	106	38
rect	105	38	106	39
rect	105	39	106	40
rect	105	40	106	41
rect	105	41	106	42
rect	105	42	106	43
rect	105	43	106	44
rect	105	44	106	45
rect	105	45	106	46
rect	105	46	106	47
rect	105	47	106	48
rect	105	48	106	49
rect	105	49	106	50
rect	105	50	106	51
rect	105	51	106	52
rect	105	52	106	53
rect	105	53	106	54
rect	105	54	106	55
rect	105	55	106	56
rect	105	56	106	57
rect	105	57	106	58
rect	105	58	106	59
rect	105	59	106	60
rect	105	60	106	61
rect	105	61	106	62
rect	105	62	106	63
rect	105	63	106	64
rect	105	64	106	65
rect	105	65	106	66
rect	105	66	106	67
rect	105	67	106	68
rect	105	68	106	69
rect	105	69	106	70
rect	105	70	106	71
rect	105	71	106	72
rect	105	72	106	73
rect	105	73	106	74
rect	105	74	106	75
rect	105	75	106	76
rect	105	76	106	77
rect	105	77	106	78
rect	105	78	106	79
rect	105	79	106	80
rect	105	80	106	81
rect	105	81	106	82
rect	105	82	106	83
rect	105	83	106	84
rect	105	84	106	85
rect	105	85	106	86
rect	105	86	106	87
rect	105	87	106	88
rect	105	88	106	89
rect	105	89	106	90
rect	105	90	106	91
rect	105	91	106	92
rect	105	92	106	93
rect	105	93	106	94
rect	105	94	106	95
rect	105	95	106	96
rect	105	96	106	97
rect	105	97	106	98
rect	105	98	106	99
rect	105	99	106	100
rect	105	100	106	101
rect	105	101	106	102
rect	105	102	106	103
rect	105	103	106	104
rect	105	104	106	105
rect	105	105	106	106
rect	105	106	106	107
rect	105	107	106	108
rect	105	108	106	109
rect	105	109	106	110
rect	105	110	106	111
rect	105	111	106	112
rect	105	112	106	113
rect	105	113	106	114
rect	105	114	106	115
rect	105	115	106	116
rect	105	116	106	117
rect	105	117	106	118
rect	105	118	106	119
rect	105	119	106	120
rect	105	120	106	121
rect	105	121	106	122
rect	105	122	106	123
rect	105	123	106	124
rect	105	124	106	125
rect	105	125	106	126
rect	105	126	106	127
rect	105	127	106	128
rect	105	128	106	129
rect	105	129	106	130
rect	105	130	106	131
rect	105	131	106	132
rect	105	132	106	133
rect	105	133	106	134
rect	105	134	106	135
rect	105	135	106	136
rect	105	136	106	137
rect	105	137	106	138
rect	105	138	106	139
rect	105	139	106	140
rect	105	140	106	141
rect	105	141	106	142
rect	105	142	106	143
rect	105	143	106	144
rect	105	144	106	145
rect	105	145	106	146
rect	105	146	106	147
rect	105	147	106	148
rect	105	148	106	149
rect	105	149	106	150
rect	105	150	106	151
rect	105	151	106	152
rect	105	152	106	153
rect	105	153	106	154
rect	105	154	106	155
rect	105	155	106	156
rect	105	156	106	157
rect	105	157	106	158
rect	105	158	106	159
rect	105	159	106	160
rect	105	160	106	161
rect	105	161	106	162
rect	105	162	106	163
rect	105	163	106	164
rect	105	164	106	165
rect	105	165	106	166
rect	105	166	106	167
rect	105	167	106	168
rect	105	168	106	169
rect	105	169	106	170
rect	105	170	106	171
rect	105	171	106	172
rect	105	172	106	173
rect	105	173	106	174
rect	105	174	106	175
rect	105	175	106	176
rect	105	176	106	177
rect	105	177	106	178
rect	105	178	106	179
rect	105	179	106	180
rect	105	180	106	181
rect	105	181	106	182
rect	105	182	106	183
rect	105	183	106	184
rect	105	184	106	185
rect	105	185	106	186
rect	105	186	106	187
rect	105	187	106	188
rect	105	188	106	189
rect	105	189	106	190
rect	105	190	106	191
rect	105	191	106	192
rect	105	192	106	193
rect	105	193	106	194
rect	105	194	106	195
rect	105	195	106	196
rect	105	196	106	197
rect	105	197	106	198
rect	105	198	106	199
rect	105	199	106	200
rect	105	200	106	201
rect	105	201	106	202
rect	105	202	106	203
rect	105	203	106	204
rect	105	204	106	205
rect	105	205	106	206
rect	105	206	106	207
rect	105	207	106	208
rect	105	208	106	209
rect	105	209	106	210
rect	105	210	106	211
rect	105	211	106	212
rect	105	212	106	213
rect	105	213	106	214
rect	105	214	106	215
rect	105	215	106	216
rect	105	216	106	217
rect	105	217	106	218
rect	105	218	106	219
rect	105	219	106	220
rect	105	220	106	221
rect	105	221	106	222
rect	105	222	106	223
rect	105	223	106	224
rect	105	224	106	225
rect	105	225	106	226
rect	105	226	106	227
rect	105	227	106	228
rect	105	228	106	229
rect	105	229	106	230
rect	105	230	106	231
rect	105	231	106	232
rect	105	232	106	233
rect	105	233	106	234
rect	105	234	106	235
rect	105	235	106	236
rect	105	236	106	237
rect	105	237	106	238
rect	105	238	106	239
rect	105	239	106	240
rect	105	240	106	241
rect	105	241	106	242
rect	105	242	106	243
rect	105	243	106	244
rect	105	244	106	245
rect	105	245	106	246
rect	105	246	106	247
rect	105	247	106	248
rect	105	248	106	249
rect	105	249	106	250
rect	105	250	106	251
rect	105	251	106	252
rect	105	252	106	253
rect	105	253	106	254
rect	105	254	106	255
rect	105	255	106	256
rect	105	256	106	257
rect	105	257	106	258
rect	105	258	106	259
rect	105	259	106	260
rect	105	260	106	261
rect	105	261	106	262
rect	105	262	106	263
rect	105	263	106	264
rect	105	264	106	265
rect	105	265	106	266
rect	105	266	106	267
rect	105	267	106	268
rect	105	268	106	269
rect	105	269	106	270
rect	105	270	106	271
rect	105	271	106	272
rect	105	272	106	273
rect	105	273	106	274
rect	105	274	106	275
rect	105	275	106	276
rect	105	276	106	277
rect	105	277	106	278
rect	105	278	106	279
rect	105	279	106	280
rect	105	280	106	281
rect	105	281	106	282
rect	105	282	106	283
rect	105	283	106	284
rect	105	284	106	285
rect	105	285	106	286
rect	105	286	106	287
rect	105	287	106	288
rect	105	288	106	289
rect	105	289	106	290
rect	105	290	106	291
rect	105	291	106	292
rect	105	292	106	293
rect	105	293	106	294
rect	105	294	106	295
rect	105	295	106	296
rect	105	296	106	297
rect	105	297	106	298
rect	105	298	106	299
rect	105	299	106	300
rect	105	300	106	301
rect	105	301	106	302
rect	105	302	106	303
rect	105	303	106	304
rect	105	304	106	305
rect	105	305	106	306
rect	105	306	106	307
rect	105	307	106	308
rect	105	308	106	309
rect	105	309	106	310
rect	105	310	106	311
rect	105	311	106	312
rect	139	0	140	1
rect	139	1	140	2
rect	139	2	140	3
rect	139	3	140	4
rect	139	4	140	5
rect	139	5	140	6
rect	139	6	140	7
rect	139	7	140	8
rect	139	8	140	9
rect	139	9	140	10
rect	139	10	140	11
rect	139	11	140	12
rect	139	12	140	13
rect	139	13	140	14
rect	139	14	140	15
rect	139	15	140	16
rect	139	16	140	17
rect	139	17	140	18
rect	139	18	140	19
rect	139	19	140	20
rect	139	20	140	21
rect	139	21	140	22
rect	139	22	140	23
rect	139	23	140	24
rect	139	24	140	25
rect	139	25	140	26
rect	139	26	140	27
rect	139	27	140	28
rect	139	28	140	29
rect	139	29	140	30
rect	139	30	140	31
rect	139	31	140	32
rect	139	32	140	33
rect	139	33	140	34
rect	139	34	140	35
rect	139	35	140	36
rect	139	36	140	37
rect	139	37	140	38
rect	139	38	140	39
rect	139	39	140	40
rect	139	40	140	41
rect	139	41	140	42
rect	139	42	140	43
rect	139	43	140	44
rect	139	44	140	45
rect	139	45	140	46
rect	139	46	140	47
rect	139	47	140	48
rect	139	48	140	49
rect	139	49	140	50
rect	139	50	140	51
rect	139	51	140	52
rect	139	52	140	53
rect	139	53	140	54
rect	139	54	140	55
rect	139	55	140	56
rect	139	56	140	57
rect	139	57	140	58
rect	139	58	140	59
rect	139	59	140	60
rect	139	60	140	61
rect	139	61	140	62
rect	139	62	140	63
rect	139	63	140	64
rect	139	64	140	65
rect	139	65	140	66
rect	139	66	140	67
rect	139	67	140	68
rect	139	68	140	69
rect	139	69	140	70
rect	139	70	140	71
rect	139	71	140	72
rect	139	72	140	73
rect	139	73	140	74
rect	139	74	140	75
rect	139	75	140	76
rect	139	76	140	77
rect	139	77	140	78
rect	139	78	140	79
rect	139	79	140	80
rect	139	80	140	81
rect	139	81	140	82
rect	139	82	140	83
rect	139	83	140	84
rect	139	84	140	85
rect	139	85	140	86
rect	139	86	140	87
rect	139	87	140	88
rect	139	88	140	89
rect	139	89	140	90
rect	139	90	140	91
rect	139	91	140	92
rect	139	92	140	93
rect	139	93	140	94
rect	139	94	140	95
rect	139	95	140	96
rect	139	96	140	97
rect	139	97	140	98
rect	139	98	140	99
rect	139	99	140	100
rect	139	100	140	101
rect	139	101	140	102
rect	139	102	140	103
rect	139	103	140	104
rect	139	104	140	105
rect	139	105	140	106
rect	139	106	140	107
rect	139	107	140	108
rect	139	108	140	109
rect	139	109	140	110
rect	139	110	140	111
rect	139	111	140	112
rect	139	112	140	113
rect	139	113	140	114
rect	139	114	140	115
rect	139	115	140	116
rect	139	116	140	117
rect	139	117	140	118
rect	139	118	140	119
rect	139	119	140	120
rect	139	120	140	121
rect	139	121	140	122
rect	139	122	140	123
rect	139	123	140	124
rect	139	124	140	125
rect	139	125	140	126
rect	139	126	140	127
rect	139	127	140	128
rect	139	128	140	129
rect	139	129	140	130
rect	139	130	140	131
rect	139	131	140	132
rect	139	132	140	133
rect	139	133	140	134
rect	139	134	140	135
rect	139	135	140	136
rect	139	136	140	137
rect	139	137	140	138
rect	139	138	140	139
rect	139	139	140	140
rect	139	140	140	141
rect	139	141	140	142
rect	139	142	140	143
rect	139	143	140	144
rect	139	144	140	145
rect	139	145	140	146
rect	139	146	140	147
rect	139	147	140	148
rect	139	148	140	149
rect	139	149	140	150
rect	139	150	140	151
rect	139	151	140	152
rect	139	152	140	153
rect	139	153	140	154
rect	139	154	140	155
rect	139	155	140	156
rect	139	156	140	157
rect	139	157	140	158
rect	139	158	140	159
rect	139	159	140	160
rect	139	160	140	161
rect	139	161	140	162
rect	139	162	140	163
rect	139	163	140	164
rect	139	164	140	165
rect	139	165	140	166
rect	139	166	140	167
rect	139	167	140	168
rect	139	168	140	169
rect	139	169	140	170
rect	139	170	140	171
rect	139	171	140	172
rect	139	172	140	173
rect	139	173	140	174
rect	139	174	140	175
rect	139	175	140	176
rect	139	176	140	177
rect	139	177	140	178
rect	139	178	140	179
rect	139	179	140	180
rect	139	180	140	181
rect	139	181	140	182
rect	139	182	140	183
rect	139	183	140	184
rect	139	184	140	185
rect	139	185	140	186
rect	139	186	140	187
rect	139	187	140	188
rect	139	188	140	189
rect	139	189	140	190
rect	139	190	140	191
rect	139	191	140	192
rect	139	192	140	193
rect	139	193	140	194
rect	139	194	140	195
rect	139	195	140	196
rect	139	196	140	197
rect	139	197	140	198
rect	139	198	140	199
rect	139	199	140	200
rect	139	200	140	201
rect	139	201	140	202
rect	139	202	140	203
rect	139	203	140	204
rect	139	204	140	205
rect	139	205	140	206
rect	139	206	140	207
rect	139	207	140	208
rect	139	208	140	209
rect	139	209	140	210
rect	139	210	140	211
rect	139	211	140	212
rect	139	212	140	213
rect	139	213	140	214
rect	139	214	140	215
rect	139	215	140	216
rect	139	216	140	217
rect	139	217	140	218
rect	139	218	140	219
rect	139	219	140	220
rect	139	220	140	221
rect	139	221	140	222
rect	139	222	140	223
rect	139	223	140	224
rect	139	224	140	225
rect	139	225	140	226
rect	139	226	140	227
rect	139	227	140	228
rect	139	228	140	229
rect	139	229	140	230
rect	139	230	140	231
rect	139	231	140	232
rect	139	232	140	233
rect	139	233	140	234
rect	139	234	140	235
rect	139	235	140	236
rect	139	236	140	237
rect	139	237	140	238
rect	139	238	140	239
rect	139	239	140	240
rect	139	240	140	241
rect	139	241	140	242
rect	139	242	140	243
rect	139	243	140	244
rect	139	244	140	245
rect	139	245	140	246
rect	139	246	140	247
rect	139	247	140	248
rect	139	248	140	249
rect	139	249	140	250
rect	139	250	140	251
rect	139	251	140	252
rect	139	252	140	253
rect	139	253	140	254
rect	139	254	140	255
rect	139	255	140	256
rect	139	256	140	257
rect	139	257	140	258
rect	139	258	140	259
rect	139	259	140	260
rect	139	260	140	261
rect	139	261	140	262
rect	139	262	140	263
rect	139	263	140	264
rect	139	264	140	265
rect	139	265	140	266
rect	139	266	140	267
rect	139	267	140	268
rect	139	268	140	269
rect	139	269	140	270
rect	139	270	140	271
rect	139	271	140	272
rect	139	272	140	273
rect	139	273	140	274
rect	139	274	140	275
rect	139	275	140	276
rect	139	276	140	277
rect	139	277	140	278
rect	139	278	140	279
rect	139	279	140	280
rect	139	280	140	281
rect	139	281	140	282
rect	139	282	140	283
rect	139	283	140	284
rect	139	284	140	285
rect	139	285	140	286
rect	139	286	140	287
rect	139	287	140	288
rect	139	288	140	289
rect	139	289	140	290
rect	139	290	140	291
rect	139	291	140	292
rect	139	292	140	293
rect	139	293	140	294
rect	139	294	140	295
rect	139	295	140	296
rect	139	296	140	297
rect	139	297	140	298
rect	139	298	140	299
rect	139	299	140	300
rect	139	300	140	301
rect	139	301	140	302
rect	139	302	140	303
rect	139	303	140	304
rect	139	304	140	305
rect	139	305	140	306
rect	139	306	140	307
rect	139	307	140	308
rect	139	308	140	309
rect	139	309	140	310
rect	139	310	140	311
rect	139	311	140	312
rect	139	312	140	313
rect	139	313	140	314
rect	139	314	140	315
rect	139	315	140	316
rect	139	316	140	317
rect	139	317	140	318
rect	139	318	140	319
rect	139	319	140	320
rect	139	320	140	321
rect	139	321	140	322
rect	139	322	140	323
rect	139	323	140	324
rect	140	0	141	1
rect	140	1	141	2
rect	140	2	141	3
rect	140	3	141	4
rect	140	4	141	5
rect	140	5	141	6
rect	140	6	141	7
rect	140	7	141	8
rect	140	8	141	9
rect	140	9	141	10
rect	140	10	141	11
rect	140	11	141	12
rect	140	12	141	13
rect	140	13	141	14
rect	140	14	141	15
rect	140	15	141	16
rect	140	16	141	17
rect	140	17	141	18
rect	140	18	141	19
rect	140	19	141	20
rect	140	20	141	21
rect	140	21	141	22
rect	140	22	141	23
rect	140	23	141	24
rect	140	24	141	25
rect	140	25	141	26
rect	140	26	141	27
rect	140	27	141	28
rect	140	28	141	29
rect	140	29	141	30
rect	140	30	141	31
rect	140	31	141	32
rect	140	32	141	33
rect	140	33	141	34
rect	140	34	141	35
rect	140	35	141	36
rect	140	36	141	37
rect	140	37	141	38
rect	140	38	141	39
rect	140	39	141	40
rect	140	40	141	41
rect	140	41	141	42
rect	140	42	141	43
rect	140	43	141	44
rect	140	44	141	45
rect	140	45	141	46
rect	140	46	141	47
rect	140	47	141	48
rect	140	48	141	49
rect	140	49	141	50
rect	140	50	141	51
rect	140	51	141	52
rect	140	52	141	53
rect	140	53	141	54
rect	140	54	141	55
rect	140	55	141	56
rect	140	56	141	57
rect	140	57	141	58
rect	140	58	141	59
rect	140	59	141	60
rect	140	60	141	61
rect	140	61	141	62
rect	140	62	141	63
rect	140	63	141	64
rect	140	64	141	65
rect	140	65	141	66
rect	140	66	141	67
rect	140	67	141	68
rect	140	68	141	69
rect	140	69	141	70
rect	140	70	141	71
rect	140	71	141	72
rect	140	72	141	73
rect	140	73	141	74
rect	140	74	141	75
rect	140	75	141	76
rect	140	76	141	77
rect	140	77	141	78
rect	140	78	141	79
rect	140	79	141	80
rect	140	80	141	81
rect	140	81	141	82
rect	140	82	141	83
rect	140	83	141	84
rect	140	84	141	85
rect	140	85	141	86
rect	140	86	141	87
rect	140	87	141	88
rect	140	88	141	89
rect	140	89	141	90
rect	140	90	141	91
rect	140	91	141	92
rect	140	92	141	93
rect	140	93	141	94
rect	140	94	141	95
rect	140	95	141	96
rect	140	96	141	97
rect	140	97	141	98
rect	140	98	141	99
rect	140	99	141	100
rect	140	100	141	101
rect	140	101	141	102
rect	140	102	141	103
rect	140	103	141	104
rect	140	104	141	105
rect	140	105	141	106
rect	140	106	141	107
rect	140	107	141	108
rect	140	108	141	109
rect	140	109	141	110
rect	140	110	141	111
rect	140	111	141	112
rect	140	112	141	113
rect	140	113	141	114
rect	140	114	141	115
rect	140	115	141	116
rect	140	116	141	117
rect	140	117	141	118
rect	140	118	141	119
rect	140	119	141	120
rect	140	120	141	121
rect	140	121	141	122
rect	140	122	141	123
rect	140	123	141	124
rect	140	124	141	125
rect	140	125	141	126
rect	140	126	141	127
rect	140	127	141	128
rect	140	128	141	129
rect	140	129	141	130
rect	140	130	141	131
rect	140	131	141	132
rect	140	132	141	133
rect	140	133	141	134
rect	140	134	141	135
rect	140	135	141	136
rect	140	136	141	137
rect	140	137	141	138
rect	140	138	141	139
rect	140	139	141	140
rect	140	140	141	141
rect	140	141	141	142
rect	140	142	141	143
rect	140	143	141	144
rect	140	144	141	145
rect	140	145	141	146
rect	140	146	141	147
rect	140	147	141	148
rect	140	148	141	149
rect	140	149	141	150
rect	140	150	141	151
rect	140	151	141	152
rect	140	152	141	153
rect	140	153	141	154
rect	140	154	141	155
rect	140	155	141	156
rect	140	156	141	157
rect	140	157	141	158
rect	140	158	141	159
rect	140	159	141	160
rect	140	160	141	161
rect	140	161	141	162
rect	140	162	141	163
rect	140	163	141	164
rect	140	164	141	165
rect	140	165	141	166
rect	140	166	141	167
rect	140	167	141	168
rect	140	168	141	169
rect	140	169	141	170
rect	140	170	141	171
rect	140	171	141	172
rect	140	172	141	173
rect	140	173	141	174
rect	140	174	141	175
rect	140	175	141	176
rect	140	176	141	177
rect	140	177	141	178
rect	140	178	141	179
rect	140	179	141	180
rect	140	180	141	181
rect	140	181	141	182
rect	140	182	141	183
rect	140	183	141	184
rect	140	184	141	185
rect	140	185	141	186
rect	140	186	141	187
rect	140	187	141	188
rect	140	188	141	189
rect	140	189	141	190
rect	140	190	141	191
rect	140	191	141	192
rect	140	192	141	193
rect	140	193	141	194
rect	140	194	141	195
rect	140	195	141	196
rect	140	196	141	197
rect	140	197	141	198
rect	140	198	141	199
rect	140	199	141	200
rect	140	200	141	201
rect	140	201	141	202
rect	140	202	141	203
rect	140	203	141	204
rect	140	204	141	205
rect	140	205	141	206
rect	140	206	141	207
rect	140	207	141	208
rect	140	208	141	209
rect	140	209	141	210
rect	140	210	141	211
rect	140	211	141	212
rect	140	212	141	213
rect	140	213	141	214
rect	140	214	141	215
rect	140	215	141	216
rect	140	216	141	217
rect	140	217	141	218
rect	140	218	141	219
rect	140	219	141	220
rect	140	220	141	221
rect	140	221	141	222
rect	140	222	141	223
rect	140	223	141	224
rect	140	224	141	225
rect	140	225	141	226
rect	140	226	141	227
rect	140	227	141	228
rect	140	228	141	229
rect	140	229	141	230
rect	140	230	141	231
rect	140	231	141	232
rect	140	232	141	233
rect	140	233	141	234
rect	140	234	141	235
rect	140	235	141	236
rect	140	236	141	237
rect	140	237	141	238
rect	140	238	141	239
rect	140	239	141	240
rect	140	240	141	241
rect	140	241	141	242
rect	140	242	141	243
rect	140	243	141	244
rect	140	244	141	245
rect	140	245	141	246
rect	140	246	141	247
rect	140	247	141	248
rect	140	248	141	249
rect	140	249	141	250
rect	140	250	141	251
rect	140	251	141	252
rect	140	252	141	253
rect	140	253	141	254
rect	140	254	141	255
rect	140	255	141	256
rect	140	256	141	257
rect	140	257	141	258
rect	140	258	141	259
rect	140	259	141	260
rect	140	260	141	261
rect	140	261	141	262
rect	140	262	141	263
rect	140	263	141	264
rect	140	264	141	265
rect	140	265	141	266
rect	140	266	141	267
rect	140	267	141	268
rect	140	268	141	269
rect	140	269	141	270
rect	140	270	141	271
rect	140	271	141	272
rect	140	272	141	273
rect	140	273	141	274
rect	140	274	141	275
rect	140	275	141	276
rect	140	276	141	277
rect	140	277	141	278
rect	140	278	141	279
rect	140	279	141	280
rect	140	280	141	281
rect	140	281	141	282
rect	140	282	141	283
rect	140	283	141	284
rect	140	284	141	285
rect	140	285	141	286
rect	140	286	141	287
rect	140	287	141	288
rect	140	288	141	289
rect	140	289	141	290
rect	140	290	141	291
rect	140	291	141	292
rect	140	292	141	293
rect	140	293	141	294
rect	140	294	141	295
rect	140	295	141	296
rect	140	296	141	297
rect	140	297	141	298
rect	140	298	141	299
rect	140	299	141	300
rect	140	300	141	301
rect	140	301	141	302
rect	140	302	141	303
rect	140	303	141	304
rect	140	304	141	305
rect	140	305	141	306
rect	140	306	141	307
rect	140	307	141	308
rect	140	308	141	309
rect	140	309	141	310
rect	140	310	141	311
rect	140	311	141	312
rect	140	312	141	313
rect	140	313	141	314
rect	140	314	141	315
rect	140	315	141	316
rect	140	316	141	317
rect	140	317	141	318
rect	140	318	141	319
rect	140	319	141	320
rect	140	320	141	321
rect	140	321	141	322
rect	140	322	141	323
rect	140	323	141	324
rect	141	0	142	1
rect	141	1	142	2
rect	141	2	142	3
rect	141	3	142	4
rect	141	4	142	5
rect	141	5	142	6
rect	141	6	142	7
rect	141	7	142	8
rect	141	8	142	9
rect	141	9	142	10
rect	141	10	142	11
rect	141	11	142	12
rect	141	12	142	13
rect	141	13	142	14
rect	141	14	142	15
rect	141	15	142	16
rect	141	16	142	17
rect	141	17	142	18
rect	141	18	142	19
rect	141	19	142	20
rect	141	20	142	21
rect	141	21	142	22
rect	141	22	142	23
rect	141	23	142	24
rect	141	24	142	25
rect	141	25	142	26
rect	141	26	142	27
rect	141	27	142	28
rect	141	28	142	29
rect	141	29	142	30
rect	141	30	142	31
rect	141	31	142	32
rect	141	32	142	33
rect	141	33	142	34
rect	141	34	142	35
rect	141	35	142	36
rect	141	36	142	37
rect	141	37	142	38
rect	141	38	142	39
rect	141	39	142	40
rect	141	40	142	41
rect	141	41	142	42
rect	141	42	142	43
rect	141	43	142	44
rect	141	44	142	45
rect	141	45	142	46
rect	141	46	142	47
rect	141	47	142	48
rect	141	48	142	49
rect	141	49	142	50
rect	141	50	142	51
rect	141	51	142	52
rect	141	52	142	53
rect	141	53	142	54
rect	141	54	142	55
rect	141	55	142	56
rect	141	56	142	57
rect	141	57	142	58
rect	141	58	142	59
rect	141	59	142	60
rect	141	60	142	61
rect	141	61	142	62
rect	141	62	142	63
rect	141	63	142	64
rect	141	64	142	65
rect	141	65	142	66
rect	141	66	142	67
rect	141	67	142	68
rect	141	68	142	69
rect	141	69	142	70
rect	141	70	142	71
rect	141	71	142	72
rect	141	72	142	73
rect	141	73	142	74
rect	141	74	142	75
rect	141	75	142	76
rect	141	76	142	77
rect	141	77	142	78
rect	141	78	142	79
rect	141	79	142	80
rect	141	80	142	81
rect	141	81	142	82
rect	141	82	142	83
rect	141	83	142	84
rect	141	84	142	85
rect	141	85	142	86
rect	141	86	142	87
rect	141	87	142	88
rect	141	88	142	89
rect	141	89	142	90
rect	141	90	142	91
rect	141	91	142	92
rect	141	92	142	93
rect	141	93	142	94
rect	141	94	142	95
rect	141	95	142	96
rect	141	96	142	97
rect	141	97	142	98
rect	141	98	142	99
rect	141	99	142	100
rect	141	100	142	101
rect	141	101	142	102
rect	141	102	142	103
rect	141	103	142	104
rect	141	104	142	105
rect	141	105	142	106
rect	141	106	142	107
rect	141	107	142	108
rect	141	108	142	109
rect	141	109	142	110
rect	141	110	142	111
rect	141	111	142	112
rect	141	112	142	113
rect	141	113	142	114
rect	141	114	142	115
rect	141	115	142	116
rect	141	116	142	117
rect	141	117	142	118
rect	141	118	142	119
rect	141	119	142	120
rect	141	120	142	121
rect	141	121	142	122
rect	141	122	142	123
rect	141	123	142	124
rect	141	124	142	125
rect	141	125	142	126
rect	141	126	142	127
rect	141	127	142	128
rect	141	128	142	129
rect	141	129	142	130
rect	141	130	142	131
rect	141	131	142	132
rect	141	132	142	133
rect	141	133	142	134
rect	141	134	142	135
rect	141	135	142	136
rect	141	136	142	137
rect	141	137	142	138
rect	141	138	142	139
rect	141	139	142	140
rect	141	140	142	141
rect	141	141	142	142
rect	141	142	142	143
rect	141	143	142	144
rect	141	144	142	145
rect	141	145	142	146
rect	141	146	142	147
rect	141	147	142	148
rect	141	148	142	149
rect	141	149	142	150
rect	141	150	142	151
rect	141	151	142	152
rect	141	152	142	153
rect	141	153	142	154
rect	141	154	142	155
rect	141	155	142	156
rect	141	156	142	157
rect	141	157	142	158
rect	141	158	142	159
rect	141	159	142	160
rect	141	160	142	161
rect	141	161	142	162
rect	141	162	142	163
rect	141	163	142	164
rect	141	164	142	165
rect	141	165	142	166
rect	141	166	142	167
rect	141	167	142	168
rect	141	168	142	169
rect	141	169	142	170
rect	141	170	142	171
rect	141	171	142	172
rect	141	172	142	173
rect	141	173	142	174
rect	141	174	142	175
rect	141	175	142	176
rect	141	176	142	177
rect	141	177	142	178
rect	141	178	142	179
rect	141	179	142	180
rect	141	180	142	181
rect	141	181	142	182
rect	141	182	142	183
rect	141	183	142	184
rect	141	184	142	185
rect	141	185	142	186
rect	141	186	142	187
rect	141	187	142	188
rect	141	188	142	189
rect	141	189	142	190
rect	141	190	142	191
rect	141	191	142	192
rect	141	192	142	193
rect	141	193	142	194
rect	141	194	142	195
rect	141	195	142	196
rect	141	196	142	197
rect	141	197	142	198
rect	141	198	142	199
rect	141	199	142	200
rect	141	200	142	201
rect	141	201	142	202
rect	141	202	142	203
rect	141	203	142	204
rect	141	204	142	205
rect	141	205	142	206
rect	141	206	142	207
rect	141	207	142	208
rect	141	208	142	209
rect	141	209	142	210
rect	141	210	142	211
rect	141	211	142	212
rect	141	212	142	213
rect	141	213	142	214
rect	141	214	142	215
rect	141	215	142	216
rect	141	216	142	217
rect	141	217	142	218
rect	141	218	142	219
rect	141	219	142	220
rect	141	220	142	221
rect	141	221	142	222
rect	141	222	142	223
rect	141	223	142	224
rect	141	224	142	225
rect	141	225	142	226
rect	141	226	142	227
rect	141	227	142	228
rect	141	228	142	229
rect	141	229	142	230
rect	141	230	142	231
rect	141	231	142	232
rect	141	232	142	233
rect	141	233	142	234
rect	141	234	142	235
rect	141	235	142	236
rect	141	236	142	237
rect	141	237	142	238
rect	141	238	142	239
rect	141	239	142	240
rect	141	240	142	241
rect	141	241	142	242
rect	141	242	142	243
rect	141	243	142	244
rect	141	244	142	245
rect	141	245	142	246
rect	141	246	142	247
rect	141	247	142	248
rect	141	248	142	249
rect	141	249	142	250
rect	141	250	142	251
rect	141	251	142	252
rect	141	252	142	253
rect	141	253	142	254
rect	141	254	142	255
rect	141	255	142	256
rect	141	256	142	257
rect	141	257	142	258
rect	141	258	142	259
rect	141	259	142	260
rect	141	260	142	261
rect	141	261	142	262
rect	141	262	142	263
rect	141	263	142	264
rect	141	264	142	265
rect	141	265	142	266
rect	141	266	142	267
rect	141	267	142	268
rect	141	268	142	269
rect	141	269	142	270
rect	141	270	142	271
rect	141	271	142	272
rect	141	272	142	273
rect	141	273	142	274
rect	141	274	142	275
rect	141	275	142	276
rect	141	276	142	277
rect	141	277	142	278
rect	141	278	142	279
rect	141	279	142	280
rect	141	280	142	281
rect	141	281	142	282
rect	141	282	142	283
rect	141	283	142	284
rect	141	284	142	285
rect	141	285	142	286
rect	141	286	142	287
rect	141	287	142	288
rect	141	288	142	289
rect	141	289	142	290
rect	141	290	142	291
rect	141	291	142	292
rect	141	292	142	293
rect	141	293	142	294
rect	141	294	142	295
rect	141	295	142	296
rect	141	296	142	297
rect	141	297	142	298
rect	141	298	142	299
rect	141	299	142	300
rect	141	300	142	301
rect	141	301	142	302
rect	141	302	142	303
rect	141	303	142	304
rect	141	304	142	305
rect	141	305	142	306
rect	141	306	142	307
rect	141	307	142	308
rect	141	308	142	309
rect	141	309	142	310
rect	141	310	142	311
rect	141	311	142	312
rect	141	312	142	313
rect	141	313	142	314
rect	141	314	142	315
rect	141	315	142	316
rect	141	316	142	317
rect	141	317	142	318
rect	141	318	142	319
rect	141	319	142	320
rect	141	320	142	321
rect	141	321	142	322
rect	141	322	142	323
rect	141	323	142	324
rect	142	0	143	1
rect	142	1	143	2
rect	142	2	143	3
rect	142	3	143	4
rect	142	4	143	5
rect	142	5	143	6
rect	142	6	143	7
rect	142	7	143	8
rect	142	8	143	9
rect	142	9	143	10
rect	142	10	143	11
rect	142	11	143	12
rect	142	12	143	13
rect	142	13	143	14
rect	142	14	143	15
rect	142	15	143	16
rect	142	16	143	17
rect	142	17	143	18
rect	142	18	143	19
rect	142	19	143	20
rect	142	20	143	21
rect	142	21	143	22
rect	142	22	143	23
rect	142	23	143	24
rect	142	24	143	25
rect	142	25	143	26
rect	142	26	143	27
rect	142	27	143	28
rect	142	28	143	29
rect	142	29	143	30
rect	142	30	143	31
rect	142	31	143	32
rect	142	32	143	33
rect	142	33	143	34
rect	142	34	143	35
rect	142	35	143	36
rect	142	36	143	37
rect	142	37	143	38
rect	142	38	143	39
rect	142	39	143	40
rect	142	40	143	41
rect	142	41	143	42
rect	142	42	143	43
rect	142	43	143	44
rect	142	44	143	45
rect	142	45	143	46
rect	142	46	143	47
rect	142	47	143	48
rect	142	48	143	49
rect	142	49	143	50
rect	142	50	143	51
rect	142	51	143	52
rect	142	52	143	53
rect	142	53	143	54
rect	142	54	143	55
rect	142	55	143	56
rect	142	56	143	57
rect	142	57	143	58
rect	142	58	143	59
rect	142	59	143	60
rect	142	60	143	61
rect	142	61	143	62
rect	142	62	143	63
rect	142	63	143	64
rect	142	64	143	65
rect	142	65	143	66
rect	142	66	143	67
rect	142	67	143	68
rect	142	68	143	69
rect	142	69	143	70
rect	142	70	143	71
rect	142	71	143	72
rect	142	72	143	73
rect	142	73	143	74
rect	142	74	143	75
rect	142	75	143	76
rect	142	76	143	77
rect	142	77	143	78
rect	142	78	143	79
rect	142	79	143	80
rect	142	80	143	81
rect	142	81	143	82
rect	142	82	143	83
rect	142	83	143	84
rect	142	84	143	85
rect	142	85	143	86
rect	142	86	143	87
rect	142	87	143	88
rect	142	88	143	89
rect	142	89	143	90
rect	142	90	143	91
rect	142	91	143	92
rect	142	92	143	93
rect	142	93	143	94
rect	142	94	143	95
rect	142	95	143	96
rect	142	96	143	97
rect	142	97	143	98
rect	142	98	143	99
rect	142	99	143	100
rect	142	100	143	101
rect	142	101	143	102
rect	142	102	143	103
rect	142	103	143	104
rect	142	104	143	105
rect	142	105	143	106
rect	142	106	143	107
rect	142	107	143	108
rect	142	108	143	109
rect	142	109	143	110
rect	142	110	143	111
rect	142	111	143	112
rect	142	112	143	113
rect	142	113	143	114
rect	142	114	143	115
rect	142	115	143	116
rect	142	116	143	117
rect	142	117	143	118
rect	142	118	143	119
rect	142	119	143	120
rect	142	120	143	121
rect	142	121	143	122
rect	142	122	143	123
rect	142	123	143	124
rect	142	124	143	125
rect	142	125	143	126
rect	142	126	143	127
rect	142	127	143	128
rect	142	128	143	129
rect	142	129	143	130
rect	142	130	143	131
rect	142	131	143	132
rect	142	132	143	133
rect	142	133	143	134
rect	142	134	143	135
rect	142	135	143	136
rect	142	136	143	137
rect	142	137	143	138
rect	142	138	143	139
rect	142	139	143	140
rect	142	140	143	141
rect	142	141	143	142
rect	142	142	143	143
rect	142	143	143	144
rect	142	144	143	145
rect	142	145	143	146
rect	142	146	143	147
rect	142	147	143	148
rect	142	148	143	149
rect	142	149	143	150
rect	142	150	143	151
rect	142	151	143	152
rect	142	152	143	153
rect	142	153	143	154
rect	142	154	143	155
rect	142	155	143	156
rect	142	156	143	157
rect	142	157	143	158
rect	142	158	143	159
rect	142	159	143	160
rect	142	160	143	161
rect	142	161	143	162
rect	142	162	143	163
rect	142	163	143	164
rect	142	164	143	165
rect	142	165	143	166
rect	142	166	143	167
rect	142	167	143	168
rect	142	168	143	169
rect	142	169	143	170
rect	142	170	143	171
rect	142	171	143	172
rect	142	172	143	173
rect	142	173	143	174
rect	142	174	143	175
rect	142	175	143	176
rect	142	176	143	177
rect	142	177	143	178
rect	142	178	143	179
rect	142	179	143	180
rect	142	180	143	181
rect	142	181	143	182
rect	142	182	143	183
rect	142	183	143	184
rect	142	184	143	185
rect	142	185	143	186
rect	142	186	143	187
rect	142	187	143	188
rect	142	188	143	189
rect	142	189	143	190
rect	142	190	143	191
rect	142	191	143	192
rect	142	192	143	193
rect	142	193	143	194
rect	142	194	143	195
rect	142	195	143	196
rect	142	196	143	197
rect	142	197	143	198
rect	142	198	143	199
rect	142	199	143	200
rect	142	200	143	201
rect	142	201	143	202
rect	142	202	143	203
rect	142	203	143	204
rect	142	204	143	205
rect	142	205	143	206
rect	142	206	143	207
rect	142	207	143	208
rect	142	208	143	209
rect	142	209	143	210
rect	142	210	143	211
rect	142	211	143	212
rect	142	212	143	213
rect	142	213	143	214
rect	142	214	143	215
rect	142	215	143	216
rect	142	216	143	217
rect	142	217	143	218
rect	142	218	143	219
rect	142	219	143	220
rect	142	220	143	221
rect	142	221	143	222
rect	142	222	143	223
rect	142	223	143	224
rect	142	224	143	225
rect	142	225	143	226
rect	142	226	143	227
rect	142	227	143	228
rect	142	228	143	229
rect	142	229	143	230
rect	142	230	143	231
rect	142	231	143	232
rect	142	232	143	233
rect	142	233	143	234
rect	142	234	143	235
rect	142	235	143	236
rect	142	236	143	237
rect	142	237	143	238
rect	142	238	143	239
rect	142	239	143	240
rect	142	240	143	241
rect	142	241	143	242
rect	142	242	143	243
rect	142	243	143	244
rect	142	244	143	245
rect	142	245	143	246
rect	142	246	143	247
rect	142	247	143	248
rect	142	248	143	249
rect	142	249	143	250
rect	142	250	143	251
rect	142	251	143	252
rect	142	252	143	253
rect	142	253	143	254
rect	142	254	143	255
rect	142	255	143	256
rect	142	256	143	257
rect	142	257	143	258
rect	142	258	143	259
rect	142	259	143	260
rect	142	260	143	261
rect	142	261	143	262
rect	142	262	143	263
rect	142	263	143	264
rect	142	264	143	265
rect	142	265	143	266
rect	142	266	143	267
rect	142	267	143	268
rect	142	268	143	269
rect	142	269	143	270
rect	142	270	143	271
rect	142	271	143	272
rect	142	272	143	273
rect	142	273	143	274
rect	142	274	143	275
rect	142	275	143	276
rect	142	276	143	277
rect	142	277	143	278
rect	142	278	143	279
rect	142	279	143	280
rect	142	280	143	281
rect	142	281	143	282
rect	142	282	143	283
rect	142	283	143	284
rect	142	284	143	285
rect	142	285	143	286
rect	142	286	143	287
rect	142	287	143	288
rect	142	288	143	289
rect	142	289	143	290
rect	142	290	143	291
rect	142	291	143	292
rect	142	292	143	293
rect	142	293	143	294
rect	142	294	143	295
rect	142	295	143	296
rect	142	296	143	297
rect	142	297	143	298
rect	142	298	143	299
rect	142	299	143	300
rect	142	300	143	301
rect	142	301	143	302
rect	142	302	143	303
rect	142	303	143	304
rect	142	304	143	305
rect	142	305	143	306
rect	142	306	143	307
rect	142	307	143	308
rect	142	308	143	309
rect	142	309	143	310
rect	142	310	143	311
rect	142	311	143	312
rect	142	312	143	313
rect	142	313	143	314
rect	142	314	143	315
rect	142	315	143	316
rect	142	316	143	317
rect	142	317	143	318
rect	142	318	143	319
rect	142	319	143	320
rect	142	320	143	321
rect	142	321	143	322
rect	142	322	143	323
rect	142	323	143	324
rect	143	0	144	1
rect	143	1	144	2
rect	143	2	144	3
rect	143	3	144	4
rect	143	4	144	5
rect	143	5	144	6
rect	143	6	144	7
rect	143	7	144	8
rect	143	8	144	9
rect	143	9	144	10
rect	143	10	144	11
rect	143	11	144	12
rect	143	12	144	13
rect	143	13	144	14
rect	143	14	144	15
rect	143	15	144	16
rect	143	16	144	17
rect	143	17	144	18
rect	143	18	144	19
rect	143	19	144	20
rect	143	20	144	21
rect	143	21	144	22
rect	143	22	144	23
rect	143	23	144	24
rect	143	24	144	25
rect	143	25	144	26
rect	143	26	144	27
rect	143	27	144	28
rect	143	28	144	29
rect	143	29	144	30
rect	143	30	144	31
rect	143	31	144	32
rect	143	32	144	33
rect	143	33	144	34
rect	143	34	144	35
rect	143	35	144	36
rect	143	36	144	37
rect	143	37	144	38
rect	143	38	144	39
rect	143	39	144	40
rect	143	40	144	41
rect	143	41	144	42
rect	143	42	144	43
rect	143	43	144	44
rect	143	44	144	45
rect	143	45	144	46
rect	143	46	144	47
rect	143	47	144	48
rect	143	48	144	49
rect	143	49	144	50
rect	143	50	144	51
rect	143	51	144	52
rect	143	52	144	53
rect	143	53	144	54
rect	143	54	144	55
rect	143	55	144	56
rect	143	56	144	57
rect	143	57	144	58
rect	143	58	144	59
rect	143	59	144	60
rect	143	60	144	61
rect	143	61	144	62
rect	143	62	144	63
rect	143	63	144	64
rect	143	64	144	65
rect	143	65	144	66
rect	143	66	144	67
rect	143	67	144	68
rect	143	68	144	69
rect	143	69	144	70
rect	143	70	144	71
rect	143	71	144	72
rect	143	72	144	73
rect	143	73	144	74
rect	143	74	144	75
rect	143	75	144	76
rect	143	76	144	77
rect	143	77	144	78
rect	143	78	144	79
rect	143	79	144	80
rect	143	80	144	81
rect	143	81	144	82
rect	143	82	144	83
rect	143	83	144	84
rect	143	84	144	85
rect	143	85	144	86
rect	143	86	144	87
rect	143	87	144	88
rect	143	88	144	89
rect	143	89	144	90
rect	143	90	144	91
rect	143	91	144	92
rect	143	92	144	93
rect	143	93	144	94
rect	143	94	144	95
rect	143	95	144	96
rect	143	96	144	97
rect	143	97	144	98
rect	143	98	144	99
rect	143	99	144	100
rect	143	100	144	101
rect	143	101	144	102
rect	143	102	144	103
rect	143	103	144	104
rect	143	104	144	105
rect	143	105	144	106
rect	143	106	144	107
rect	143	107	144	108
rect	143	108	144	109
rect	143	109	144	110
rect	143	110	144	111
rect	143	111	144	112
rect	143	112	144	113
rect	143	113	144	114
rect	143	114	144	115
rect	143	115	144	116
rect	143	116	144	117
rect	143	117	144	118
rect	143	118	144	119
rect	143	119	144	120
rect	143	120	144	121
rect	143	121	144	122
rect	143	122	144	123
rect	143	123	144	124
rect	143	124	144	125
rect	143	125	144	126
rect	143	126	144	127
rect	143	127	144	128
rect	143	128	144	129
rect	143	129	144	130
rect	143	130	144	131
rect	143	131	144	132
rect	143	132	144	133
rect	143	133	144	134
rect	143	134	144	135
rect	143	135	144	136
rect	143	136	144	137
rect	143	137	144	138
rect	143	138	144	139
rect	143	139	144	140
rect	143	140	144	141
rect	143	141	144	142
rect	143	142	144	143
rect	143	143	144	144
rect	143	144	144	145
rect	143	145	144	146
rect	143	146	144	147
rect	143	147	144	148
rect	143	148	144	149
rect	143	149	144	150
rect	143	150	144	151
rect	143	151	144	152
rect	143	152	144	153
rect	143	153	144	154
rect	143	154	144	155
rect	143	155	144	156
rect	143	156	144	157
rect	143	157	144	158
rect	143	158	144	159
rect	143	159	144	160
rect	143	160	144	161
rect	143	161	144	162
rect	143	162	144	163
rect	143	163	144	164
rect	143	164	144	165
rect	143	165	144	166
rect	143	166	144	167
rect	143	167	144	168
rect	143	168	144	169
rect	143	169	144	170
rect	143	170	144	171
rect	143	171	144	172
rect	143	172	144	173
rect	143	173	144	174
rect	143	174	144	175
rect	143	175	144	176
rect	143	176	144	177
rect	143	177	144	178
rect	143	178	144	179
rect	143	179	144	180
rect	143	180	144	181
rect	143	181	144	182
rect	143	182	144	183
rect	143	183	144	184
rect	143	184	144	185
rect	143	185	144	186
rect	143	186	144	187
rect	143	187	144	188
rect	143	188	144	189
rect	143	189	144	190
rect	143	190	144	191
rect	143	191	144	192
rect	143	192	144	193
rect	143	193	144	194
rect	143	194	144	195
rect	143	195	144	196
rect	143	196	144	197
rect	143	197	144	198
rect	143	198	144	199
rect	143	199	144	200
rect	143	200	144	201
rect	143	201	144	202
rect	143	202	144	203
rect	143	203	144	204
rect	143	204	144	205
rect	143	205	144	206
rect	143	206	144	207
rect	143	207	144	208
rect	143	208	144	209
rect	143	209	144	210
rect	143	210	144	211
rect	143	211	144	212
rect	143	212	144	213
rect	143	213	144	214
rect	143	214	144	215
rect	143	215	144	216
rect	143	216	144	217
rect	143	217	144	218
rect	143	218	144	219
rect	143	219	144	220
rect	143	220	144	221
rect	143	221	144	222
rect	143	222	144	223
rect	143	223	144	224
rect	143	224	144	225
rect	143	225	144	226
rect	143	226	144	227
rect	143	227	144	228
rect	143	228	144	229
rect	143	229	144	230
rect	143	230	144	231
rect	143	231	144	232
rect	143	232	144	233
rect	143	233	144	234
rect	143	234	144	235
rect	143	235	144	236
rect	143	236	144	237
rect	143	237	144	238
rect	143	238	144	239
rect	143	239	144	240
rect	143	240	144	241
rect	143	241	144	242
rect	143	242	144	243
rect	143	243	144	244
rect	143	244	144	245
rect	143	245	144	246
rect	143	246	144	247
rect	143	247	144	248
rect	143	248	144	249
rect	143	249	144	250
rect	143	250	144	251
rect	143	251	144	252
rect	143	252	144	253
rect	143	253	144	254
rect	143	254	144	255
rect	143	255	144	256
rect	143	256	144	257
rect	143	257	144	258
rect	143	258	144	259
rect	143	259	144	260
rect	143	260	144	261
rect	143	261	144	262
rect	143	262	144	263
rect	143	263	144	264
rect	143	264	144	265
rect	143	265	144	266
rect	143	266	144	267
rect	143	267	144	268
rect	143	268	144	269
rect	143	269	144	270
rect	143	270	144	271
rect	143	271	144	272
rect	143	272	144	273
rect	143	273	144	274
rect	143	274	144	275
rect	143	275	144	276
rect	143	276	144	277
rect	143	277	144	278
rect	143	278	144	279
rect	143	279	144	280
rect	143	280	144	281
rect	143	281	144	282
rect	143	282	144	283
rect	143	283	144	284
rect	143	284	144	285
rect	143	285	144	286
rect	143	286	144	287
rect	143	287	144	288
rect	143	288	144	289
rect	143	289	144	290
rect	143	290	144	291
rect	143	291	144	292
rect	143	292	144	293
rect	143	293	144	294
rect	143	294	144	295
rect	143	295	144	296
rect	143	296	144	297
rect	143	297	144	298
rect	143	298	144	299
rect	143	299	144	300
rect	143	300	144	301
rect	143	301	144	302
rect	143	302	144	303
rect	143	303	144	304
rect	143	304	144	305
rect	143	305	144	306
rect	143	306	144	307
rect	143	307	144	308
rect	143	308	144	309
rect	143	309	144	310
rect	143	310	144	311
rect	143	311	144	312
rect	143	312	144	313
rect	143	313	144	314
rect	143	314	144	315
rect	143	315	144	316
rect	143	316	144	317
rect	143	317	144	318
rect	143	318	144	319
rect	143	319	144	320
rect	143	320	144	321
rect	143	321	144	322
rect	143	322	144	323
rect	143	323	144	324
rect	144	0	145	1
rect	144	1	145	2
rect	144	2	145	3
rect	144	3	145	4
rect	144	4	145	5
rect	144	5	145	6
rect	144	6	145	7
rect	144	7	145	8
rect	144	8	145	9
rect	144	9	145	10
rect	144	10	145	11
rect	144	11	145	12
rect	144	12	145	13
rect	144	13	145	14
rect	144	14	145	15
rect	144	15	145	16
rect	144	16	145	17
rect	144	17	145	18
rect	144	18	145	19
rect	144	19	145	20
rect	144	20	145	21
rect	144	21	145	22
rect	144	22	145	23
rect	144	23	145	24
rect	144	24	145	25
rect	144	25	145	26
rect	144	26	145	27
rect	144	27	145	28
rect	144	28	145	29
rect	144	29	145	30
rect	144	30	145	31
rect	144	31	145	32
rect	144	32	145	33
rect	144	33	145	34
rect	144	34	145	35
rect	144	35	145	36
rect	144	36	145	37
rect	144	37	145	38
rect	144	38	145	39
rect	144	39	145	40
rect	144	40	145	41
rect	144	41	145	42
rect	144	42	145	43
rect	144	43	145	44
rect	144	44	145	45
rect	144	45	145	46
rect	144	46	145	47
rect	144	47	145	48
rect	144	48	145	49
rect	144	49	145	50
rect	144	50	145	51
rect	144	51	145	52
rect	144	52	145	53
rect	144	53	145	54
rect	144	54	145	55
rect	144	55	145	56
rect	144	56	145	57
rect	144	57	145	58
rect	144	58	145	59
rect	144	59	145	60
rect	144	60	145	61
rect	144	61	145	62
rect	144	62	145	63
rect	144	63	145	64
rect	144	64	145	65
rect	144	65	145	66
rect	144	66	145	67
rect	144	67	145	68
rect	144	68	145	69
rect	144	69	145	70
rect	144	70	145	71
rect	144	71	145	72
rect	144	72	145	73
rect	144	73	145	74
rect	144	74	145	75
rect	144	75	145	76
rect	144	76	145	77
rect	144	77	145	78
rect	144	78	145	79
rect	144	79	145	80
rect	144	80	145	81
rect	144	81	145	82
rect	144	82	145	83
rect	144	83	145	84
rect	144	84	145	85
rect	144	85	145	86
rect	144	86	145	87
rect	144	87	145	88
rect	144	88	145	89
rect	144	89	145	90
rect	144	90	145	91
rect	144	91	145	92
rect	144	92	145	93
rect	144	93	145	94
rect	144	94	145	95
rect	144	95	145	96
rect	144	96	145	97
rect	144	97	145	98
rect	144	98	145	99
rect	144	99	145	100
rect	144	100	145	101
rect	144	101	145	102
rect	144	102	145	103
rect	144	103	145	104
rect	144	104	145	105
rect	144	105	145	106
rect	144	106	145	107
rect	144	107	145	108
rect	144	108	145	109
rect	144	109	145	110
rect	144	110	145	111
rect	144	111	145	112
rect	144	112	145	113
rect	144	113	145	114
rect	144	114	145	115
rect	144	115	145	116
rect	144	116	145	117
rect	144	117	145	118
rect	144	118	145	119
rect	144	119	145	120
rect	144	120	145	121
rect	144	121	145	122
rect	144	122	145	123
rect	144	123	145	124
rect	144	124	145	125
rect	144	125	145	126
rect	144	126	145	127
rect	144	127	145	128
rect	144	128	145	129
rect	144	129	145	130
rect	144	130	145	131
rect	144	131	145	132
rect	144	132	145	133
rect	144	133	145	134
rect	144	134	145	135
rect	144	135	145	136
rect	144	136	145	137
rect	144	137	145	138
rect	144	138	145	139
rect	144	139	145	140
rect	144	140	145	141
rect	144	141	145	142
rect	144	142	145	143
rect	144	143	145	144
rect	144	144	145	145
rect	144	145	145	146
rect	144	146	145	147
rect	144	147	145	148
rect	144	148	145	149
rect	144	149	145	150
rect	144	150	145	151
rect	144	151	145	152
rect	144	152	145	153
rect	144	153	145	154
rect	144	154	145	155
rect	144	155	145	156
rect	144	156	145	157
rect	144	157	145	158
rect	144	158	145	159
rect	144	159	145	160
rect	144	160	145	161
rect	144	161	145	162
rect	144	162	145	163
rect	144	163	145	164
rect	144	164	145	165
rect	144	165	145	166
rect	144	166	145	167
rect	144	167	145	168
rect	144	168	145	169
rect	144	169	145	170
rect	144	170	145	171
rect	144	171	145	172
rect	144	172	145	173
rect	144	173	145	174
rect	144	174	145	175
rect	144	175	145	176
rect	144	176	145	177
rect	144	177	145	178
rect	144	178	145	179
rect	144	179	145	180
rect	144	180	145	181
rect	144	181	145	182
rect	144	182	145	183
rect	144	183	145	184
rect	144	184	145	185
rect	144	185	145	186
rect	144	186	145	187
rect	144	187	145	188
rect	144	188	145	189
rect	144	189	145	190
rect	144	190	145	191
rect	144	191	145	192
rect	144	192	145	193
rect	144	193	145	194
rect	144	194	145	195
rect	144	195	145	196
rect	144	196	145	197
rect	144	197	145	198
rect	144	198	145	199
rect	144	199	145	200
rect	144	200	145	201
rect	144	201	145	202
rect	144	202	145	203
rect	144	203	145	204
rect	144	204	145	205
rect	144	205	145	206
rect	144	206	145	207
rect	144	207	145	208
rect	144	208	145	209
rect	144	209	145	210
rect	144	210	145	211
rect	144	211	145	212
rect	144	212	145	213
rect	144	213	145	214
rect	144	214	145	215
rect	144	215	145	216
rect	144	216	145	217
rect	144	217	145	218
rect	144	218	145	219
rect	144	219	145	220
rect	144	220	145	221
rect	144	221	145	222
rect	144	222	145	223
rect	144	223	145	224
rect	144	224	145	225
rect	144	225	145	226
rect	144	226	145	227
rect	144	227	145	228
rect	144	228	145	229
rect	144	229	145	230
rect	144	230	145	231
rect	144	231	145	232
rect	144	232	145	233
rect	144	233	145	234
rect	144	234	145	235
rect	144	235	145	236
rect	144	236	145	237
rect	144	237	145	238
rect	144	238	145	239
rect	144	239	145	240
rect	144	240	145	241
rect	144	241	145	242
rect	144	242	145	243
rect	144	243	145	244
rect	144	244	145	245
rect	144	245	145	246
rect	144	246	145	247
rect	144	247	145	248
rect	144	248	145	249
rect	144	249	145	250
rect	144	250	145	251
rect	144	251	145	252
rect	144	252	145	253
rect	144	253	145	254
rect	144	254	145	255
rect	144	255	145	256
rect	144	256	145	257
rect	144	257	145	258
rect	144	258	145	259
rect	144	259	145	260
rect	144	260	145	261
rect	144	261	145	262
rect	144	262	145	263
rect	144	263	145	264
rect	144	264	145	265
rect	144	265	145	266
rect	144	266	145	267
rect	144	267	145	268
rect	144	268	145	269
rect	144	269	145	270
rect	144	270	145	271
rect	144	271	145	272
rect	144	272	145	273
rect	144	273	145	274
rect	144	274	145	275
rect	144	275	145	276
rect	144	276	145	277
rect	144	277	145	278
rect	144	278	145	279
rect	144	279	145	280
rect	144	280	145	281
rect	144	281	145	282
rect	144	282	145	283
rect	144	283	145	284
rect	144	284	145	285
rect	144	285	145	286
rect	144	286	145	287
rect	144	287	145	288
rect	144	288	145	289
rect	144	289	145	290
rect	144	290	145	291
rect	144	291	145	292
rect	144	292	145	293
rect	144	293	145	294
rect	144	294	145	295
rect	144	295	145	296
rect	144	296	145	297
rect	144	297	145	298
rect	144	298	145	299
rect	144	299	145	300
rect	144	300	145	301
rect	144	301	145	302
rect	144	302	145	303
rect	144	303	145	304
rect	144	304	145	305
rect	144	305	145	306
rect	144	306	145	307
rect	144	307	145	308
rect	144	308	145	309
rect	144	309	145	310
rect	144	310	145	311
rect	144	311	145	312
rect	144	312	145	313
rect	144	313	145	314
rect	144	314	145	315
rect	144	315	145	316
rect	144	316	145	317
rect	144	317	145	318
rect	144	318	145	319
rect	144	319	145	320
rect	144	320	145	321
rect	144	321	145	322
rect	144	322	145	323
rect	144	323	145	324
rect	172	0	173	1
rect	172	1	173	2
rect	172	2	173	3
rect	172	3	173	4
rect	172	4	173	5
rect	172	5	173	6
rect	172	6	173	7
rect	172	7	173	8
rect	172	8	173	9
rect	172	9	173	10
rect	172	10	173	11
rect	172	11	173	12
rect	172	12	173	13
rect	172	13	173	14
rect	172	14	173	15
rect	172	15	173	16
rect	172	16	173	17
rect	172	17	173	18
rect	172	18	173	19
rect	172	19	173	20
rect	172	20	173	21
rect	172	21	173	22
rect	172	22	173	23
rect	172	23	173	24
rect	172	24	173	25
rect	172	25	173	26
rect	172	26	173	27
rect	172	27	173	28
rect	172	28	173	29
rect	172	29	173	30
rect	172	30	173	31
rect	172	31	173	32
rect	172	32	173	33
rect	172	33	173	34
rect	172	34	173	35
rect	172	35	173	36
rect	172	36	173	37
rect	172	37	173	38
rect	172	38	173	39
rect	172	39	173	40
rect	172	40	173	41
rect	172	41	173	42
rect	172	42	173	43
rect	172	43	173	44
rect	172	44	173	45
rect	172	45	173	46
rect	172	46	173	47
rect	172	47	173	48
rect	172	48	173	49
rect	172	49	173	50
rect	172	50	173	51
rect	172	51	173	52
rect	172	52	173	53
rect	172	53	173	54
rect	172	54	173	55
rect	172	55	173	56
rect	172	56	173	57
rect	172	57	173	58
rect	172	58	173	59
rect	172	59	173	60
rect	172	60	173	61
rect	172	61	173	62
rect	172	62	173	63
rect	172	63	173	64
rect	172	64	173	65
rect	172	65	173	66
rect	172	66	173	67
rect	172	67	173	68
rect	172	68	173	69
rect	172	69	173	70
rect	172	70	173	71
rect	172	71	173	72
rect	172	72	173	73
rect	172	73	173	74
rect	172	74	173	75
rect	172	75	173	76
rect	172	76	173	77
rect	172	77	173	78
rect	172	78	173	79
rect	172	79	173	80
rect	172	80	173	81
rect	172	81	173	82
rect	172	82	173	83
rect	172	83	173	84
rect	172	84	173	85
rect	172	85	173	86
rect	172	86	173	87
rect	172	87	173	88
rect	172	88	173	89
rect	172	89	173	90
rect	172	90	173	91
rect	172	91	173	92
rect	172	92	173	93
rect	172	93	173	94
rect	172	94	173	95
rect	172	95	173	96
rect	172	96	173	97
rect	172	97	173	98
rect	172	98	173	99
rect	172	99	173	100
rect	172	100	173	101
rect	172	101	173	102
rect	172	102	173	103
rect	172	103	173	104
rect	172	104	173	105
rect	172	105	173	106
rect	172	106	173	107
rect	172	107	173	108
rect	172	108	173	109
rect	172	109	173	110
rect	172	110	173	111
rect	172	111	173	112
rect	172	112	173	113
rect	172	113	173	114
rect	172	114	173	115
rect	172	115	173	116
rect	172	116	173	117
rect	172	117	173	118
rect	172	118	173	119
rect	172	119	173	120
rect	172	120	173	121
rect	172	121	173	122
rect	172	122	173	123
rect	172	123	173	124
rect	172	124	173	125
rect	172	125	173	126
rect	172	126	173	127
rect	172	127	173	128
rect	172	128	173	129
rect	172	129	173	130
rect	172	130	173	131
rect	172	131	173	132
rect	172	132	173	133
rect	172	133	173	134
rect	172	134	173	135
rect	172	135	173	136
rect	172	136	173	137
rect	172	137	173	138
rect	172	138	173	139
rect	172	139	173	140
rect	172	140	173	141
rect	172	141	173	142
rect	172	142	173	143
rect	172	143	173	144
rect	172	144	173	145
rect	172	145	173	146
rect	172	146	173	147
rect	172	147	173	148
rect	172	148	173	149
rect	172	149	173	150
rect	172	150	173	151
rect	172	151	173	152
rect	172	152	173	153
rect	172	153	173	154
rect	172	154	173	155
rect	172	155	173	156
rect	172	156	173	157
rect	172	157	173	158
rect	172	158	173	159
rect	172	159	173	160
rect	172	160	173	161
rect	172	161	173	162
rect	172	162	173	163
rect	172	163	173	164
rect	172	164	173	165
rect	172	165	173	166
rect	172	166	173	167
rect	172	167	173	168
rect	172	168	173	169
rect	172	169	173	170
rect	172	170	173	171
rect	172	171	173	172
rect	172	172	173	173
rect	172	173	173	174
rect	172	174	173	175
rect	172	175	173	176
rect	172	176	173	177
rect	172	177	173	178
rect	172	178	173	179
rect	172	179	173	180
rect	172	180	173	181
rect	172	181	173	182
rect	172	182	173	183
rect	172	183	173	184
rect	172	184	173	185
rect	172	185	173	186
rect	172	186	173	187
rect	172	187	173	188
rect	172	188	173	189
rect	172	189	173	190
rect	172	190	173	191
rect	172	191	173	192
rect	172	192	173	193
rect	172	193	173	194
rect	172	194	173	195
rect	172	195	173	196
rect	172	196	173	197
rect	172	197	173	198
rect	172	198	173	199
rect	172	199	173	200
rect	172	200	173	201
rect	172	201	173	202
rect	172	202	173	203
rect	172	203	173	204
rect	172	204	173	205
rect	172	205	173	206
rect	172	206	173	207
rect	172	207	173	208
rect	172	208	173	209
rect	172	209	173	210
rect	172	210	173	211
rect	172	211	173	212
rect	172	212	173	213
rect	172	213	173	214
rect	172	214	173	215
rect	172	215	173	216
rect	172	216	173	217
rect	172	217	173	218
rect	172	218	173	219
rect	172	219	173	220
rect	172	220	173	221
rect	172	221	173	222
rect	172	222	173	223
rect	172	223	173	224
rect	172	224	173	225
rect	172	225	173	226
rect	172	226	173	227
rect	172	227	173	228
rect	172	228	173	229
rect	172	229	173	230
rect	172	230	173	231
rect	172	231	173	232
rect	172	232	173	233
rect	172	233	173	234
rect	172	234	173	235
rect	172	235	173	236
rect	172	236	173	237
rect	172	237	173	238
rect	172	238	173	239
rect	172	239	173	240
rect	172	240	173	241
rect	172	241	173	242
rect	172	242	173	243
rect	172	243	173	244
rect	172	244	173	245
rect	172	245	173	246
rect	172	246	173	247
rect	172	247	173	248
rect	172	248	173	249
rect	172	249	173	250
rect	172	250	173	251
rect	172	251	173	252
rect	172	252	173	253
rect	172	253	173	254
rect	172	254	173	255
rect	172	255	173	256
rect	172	256	173	257
rect	172	257	173	258
rect	172	258	173	259
rect	172	259	173	260
rect	172	260	173	261
rect	172	261	173	262
rect	172	262	173	263
rect	172	263	173	264
rect	172	264	173	265
rect	172	265	173	266
rect	172	266	173	267
rect	172	267	173	268
rect	172	268	173	269
rect	172	269	173	270
rect	172	270	173	271
rect	172	271	173	272
rect	172	272	173	273
rect	172	273	173	274
rect	172	274	173	275
rect	172	275	173	276
rect	172	276	173	277
rect	172	277	173	278
rect	172	278	173	279
rect	172	279	173	280
rect	172	280	173	281
rect	172	281	173	282
rect	172	282	173	283
rect	172	283	173	284
rect	172	284	173	285
rect	172	285	173	286
rect	172	286	173	287
rect	172	287	173	288
rect	172	288	173	289
rect	172	289	173	290
rect	172	290	173	291
rect	172	291	173	292
rect	172	292	173	293
rect	172	293	173	294
rect	172	294	173	295
rect	172	295	173	296
rect	172	296	173	297
rect	172	297	173	298
rect	172	298	173	299
rect	172	299	173	300
rect	172	300	173	301
rect	172	301	173	302
rect	172	302	173	303
rect	172	303	173	304
rect	172	304	173	305
rect	172	305	173	306
rect	172	306	173	307
rect	172	307	173	308
rect	172	308	173	309
rect	172	309	173	310
rect	172	310	173	311
rect	172	311	173	312
rect	172	312	173	313
rect	172	313	173	314
rect	172	314	173	315
rect	172	315	173	316
rect	172	316	173	317
rect	172	317	173	318
rect	172	318	173	319
rect	172	319	173	320
rect	172	320	173	321
rect	172	321	173	322
rect	172	322	173	323
rect	172	323	173	324
rect	172	324	173	325
rect	172	325	173	326
rect	172	326	173	327
rect	172	327	173	328
rect	172	328	173	329
rect	172	329	173	330
rect	173	0	174	1
rect	173	1	174	2
rect	173	2	174	3
rect	173	3	174	4
rect	173	4	174	5
rect	173	5	174	6
rect	173	6	174	7
rect	173	7	174	8
rect	173	8	174	9
rect	173	9	174	10
rect	173	10	174	11
rect	173	11	174	12
rect	173	12	174	13
rect	173	13	174	14
rect	173	14	174	15
rect	173	15	174	16
rect	173	16	174	17
rect	173	17	174	18
rect	173	18	174	19
rect	173	19	174	20
rect	173	20	174	21
rect	173	21	174	22
rect	173	22	174	23
rect	173	23	174	24
rect	173	24	174	25
rect	173	25	174	26
rect	173	26	174	27
rect	173	27	174	28
rect	173	28	174	29
rect	173	29	174	30
rect	173	30	174	31
rect	173	31	174	32
rect	173	32	174	33
rect	173	33	174	34
rect	173	34	174	35
rect	173	35	174	36
rect	173	36	174	37
rect	173	37	174	38
rect	173	38	174	39
rect	173	39	174	40
rect	173	40	174	41
rect	173	41	174	42
rect	173	42	174	43
rect	173	43	174	44
rect	173	44	174	45
rect	173	45	174	46
rect	173	46	174	47
rect	173	47	174	48
rect	173	48	174	49
rect	173	49	174	50
rect	173	50	174	51
rect	173	51	174	52
rect	173	52	174	53
rect	173	53	174	54
rect	173	54	174	55
rect	173	55	174	56
rect	173	56	174	57
rect	173	57	174	58
rect	173	58	174	59
rect	173	59	174	60
rect	173	60	174	61
rect	173	61	174	62
rect	173	62	174	63
rect	173	63	174	64
rect	173	64	174	65
rect	173	65	174	66
rect	173	66	174	67
rect	173	67	174	68
rect	173	68	174	69
rect	173	69	174	70
rect	173	70	174	71
rect	173	71	174	72
rect	173	72	174	73
rect	173	73	174	74
rect	173	74	174	75
rect	173	75	174	76
rect	173	76	174	77
rect	173	77	174	78
rect	173	78	174	79
rect	173	79	174	80
rect	173	80	174	81
rect	173	81	174	82
rect	173	82	174	83
rect	173	83	174	84
rect	173	84	174	85
rect	173	85	174	86
rect	173	86	174	87
rect	173	87	174	88
rect	173	88	174	89
rect	173	89	174	90
rect	173	90	174	91
rect	173	91	174	92
rect	173	92	174	93
rect	173	93	174	94
rect	173	94	174	95
rect	173	95	174	96
rect	173	96	174	97
rect	173	97	174	98
rect	173	98	174	99
rect	173	99	174	100
rect	173	100	174	101
rect	173	101	174	102
rect	173	102	174	103
rect	173	103	174	104
rect	173	104	174	105
rect	173	105	174	106
rect	173	106	174	107
rect	173	107	174	108
rect	173	108	174	109
rect	173	109	174	110
rect	173	110	174	111
rect	173	111	174	112
rect	173	112	174	113
rect	173	113	174	114
rect	173	114	174	115
rect	173	115	174	116
rect	173	116	174	117
rect	173	117	174	118
rect	173	118	174	119
rect	173	119	174	120
rect	173	120	174	121
rect	173	121	174	122
rect	173	122	174	123
rect	173	123	174	124
rect	173	124	174	125
rect	173	125	174	126
rect	173	126	174	127
rect	173	127	174	128
rect	173	128	174	129
rect	173	129	174	130
rect	173	130	174	131
rect	173	131	174	132
rect	173	132	174	133
rect	173	133	174	134
rect	173	134	174	135
rect	173	135	174	136
rect	173	136	174	137
rect	173	137	174	138
rect	173	138	174	139
rect	173	139	174	140
rect	173	140	174	141
rect	173	141	174	142
rect	173	142	174	143
rect	173	143	174	144
rect	173	144	174	145
rect	173	145	174	146
rect	173	146	174	147
rect	173	147	174	148
rect	173	148	174	149
rect	173	149	174	150
rect	173	150	174	151
rect	173	151	174	152
rect	173	152	174	153
rect	173	153	174	154
rect	173	154	174	155
rect	173	155	174	156
rect	173	156	174	157
rect	173	157	174	158
rect	173	158	174	159
rect	173	159	174	160
rect	173	160	174	161
rect	173	161	174	162
rect	173	162	174	163
rect	173	163	174	164
rect	173	164	174	165
rect	173	165	174	166
rect	173	166	174	167
rect	173	167	174	168
rect	173	168	174	169
rect	173	169	174	170
rect	173	170	174	171
rect	173	171	174	172
rect	173	172	174	173
rect	173	173	174	174
rect	173	174	174	175
rect	173	175	174	176
rect	173	176	174	177
rect	173	177	174	178
rect	173	178	174	179
rect	173	179	174	180
rect	173	180	174	181
rect	173	181	174	182
rect	173	182	174	183
rect	173	183	174	184
rect	173	184	174	185
rect	173	185	174	186
rect	173	186	174	187
rect	173	187	174	188
rect	173	188	174	189
rect	173	189	174	190
rect	173	190	174	191
rect	173	191	174	192
rect	173	192	174	193
rect	173	193	174	194
rect	173	194	174	195
rect	173	195	174	196
rect	173	196	174	197
rect	173	197	174	198
rect	173	198	174	199
rect	173	199	174	200
rect	173	200	174	201
rect	173	201	174	202
rect	173	202	174	203
rect	173	203	174	204
rect	173	204	174	205
rect	173	205	174	206
rect	173	206	174	207
rect	173	207	174	208
rect	173	208	174	209
rect	173	209	174	210
rect	173	210	174	211
rect	173	211	174	212
rect	173	212	174	213
rect	173	213	174	214
rect	173	214	174	215
rect	173	215	174	216
rect	173	216	174	217
rect	173	217	174	218
rect	173	218	174	219
rect	173	219	174	220
rect	173	220	174	221
rect	173	221	174	222
rect	173	222	174	223
rect	173	223	174	224
rect	173	224	174	225
rect	173	225	174	226
rect	173	226	174	227
rect	173	227	174	228
rect	173	228	174	229
rect	173	229	174	230
rect	173	230	174	231
rect	173	231	174	232
rect	173	232	174	233
rect	173	233	174	234
rect	173	234	174	235
rect	173	235	174	236
rect	173	236	174	237
rect	173	237	174	238
rect	173	238	174	239
rect	173	239	174	240
rect	173	240	174	241
rect	173	241	174	242
rect	173	242	174	243
rect	173	243	174	244
rect	173	244	174	245
rect	173	245	174	246
rect	173	246	174	247
rect	173	247	174	248
rect	173	248	174	249
rect	173	249	174	250
rect	173	250	174	251
rect	173	251	174	252
rect	173	252	174	253
rect	173	253	174	254
rect	173	254	174	255
rect	173	255	174	256
rect	173	256	174	257
rect	173	257	174	258
rect	173	258	174	259
rect	173	259	174	260
rect	173	260	174	261
rect	173	261	174	262
rect	173	262	174	263
rect	173	263	174	264
rect	173	264	174	265
rect	173	265	174	266
rect	173	266	174	267
rect	173	267	174	268
rect	173	268	174	269
rect	173	269	174	270
rect	173	270	174	271
rect	173	271	174	272
rect	173	272	174	273
rect	173	273	174	274
rect	173	274	174	275
rect	173	275	174	276
rect	173	276	174	277
rect	173	277	174	278
rect	173	278	174	279
rect	173	279	174	280
rect	173	280	174	281
rect	173	281	174	282
rect	173	282	174	283
rect	173	283	174	284
rect	173	284	174	285
rect	173	285	174	286
rect	173	286	174	287
rect	173	287	174	288
rect	173	288	174	289
rect	173	289	174	290
rect	173	290	174	291
rect	173	291	174	292
rect	173	292	174	293
rect	173	293	174	294
rect	173	294	174	295
rect	173	295	174	296
rect	173	296	174	297
rect	173	297	174	298
rect	173	298	174	299
rect	173	299	174	300
rect	173	300	174	301
rect	173	301	174	302
rect	173	302	174	303
rect	173	303	174	304
rect	173	304	174	305
rect	173	305	174	306
rect	173	306	174	307
rect	173	307	174	308
rect	173	308	174	309
rect	173	309	174	310
rect	173	310	174	311
rect	173	311	174	312
rect	173	312	174	313
rect	173	313	174	314
rect	173	314	174	315
rect	173	315	174	316
rect	173	316	174	317
rect	173	317	174	318
rect	173	318	174	319
rect	173	319	174	320
rect	173	320	174	321
rect	173	321	174	322
rect	173	322	174	323
rect	173	323	174	324
rect	173	324	174	325
rect	173	325	174	326
rect	173	326	174	327
rect	173	327	174	328
rect	173	328	174	329
rect	173	329	174	330
rect	174	0	175	1
rect	174	1	175	2
rect	174	2	175	3
rect	174	3	175	4
rect	174	4	175	5
rect	174	5	175	6
rect	174	6	175	7
rect	174	7	175	8
rect	174	8	175	9
rect	174	9	175	10
rect	174	10	175	11
rect	174	11	175	12
rect	174	12	175	13
rect	174	13	175	14
rect	174	14	175	15
rect	174	15	175	16
rect	174	16	175	17
rect	174	17	175	18
rect	174	18	175	19
rect	174	19	175	20
rect	174	20	175	21
rect	174	21	175	22
rect	174	22	175	23
rect	174	23	175	24
rect	174	24	175	25
rect	174	25	175	26
rect	174	26	175	27
rect	174	27	175	28
rect	174	28	175	29
rect	174	29	175	30
rect	174	30	175	31
rect	174	31	175	32
rect	174	32	175	33
rect	174	33	175	34
rect	174	34	175	35
rect	174	35	175	36
rect	174	36	175	37
rect	174	37	175	38
rect	174	38	175	39
rect	174	39	175	40
rect	174	40	175	41
rect	174	41	175	42
rect	174	42	175	43
rect	174	43	175	44
rect	174	44	175	45
rect	174	45	175	46
rect	174	46	175	47
rect	174	47	175	48
rect	174	48	175	49
rect	174	49	175	50
rect	174	50	175	51
rect	174	51	175	52
rect	174	52	175	53
rect	174	53	175	54
rect	174	54	175	55
rect	174	55	175	56
rect	174	56	175	57
rect	174	57	175	58
rect	174	58	175	59
rect	174	59	175	60
rect	174	60	175	61
rect	174	61	175	62
rect	174	62	175	63
rect	174	63	175	64
rect	174	64	175	65
rect	174	65	175	66
rect	174	66	175	67
rect	174	67	175	68
rect	174	68	175	69
rect	174	69	175	70
rect	174	70	175	71
rect	174	71	175	72
rect	174	72	175	73
rect	174	73	175	74
rect	174	74	175	75
rect	174	75	175	76
rect	174	76	175	77
rect	174	77	175	78
rect	174	78	175	79
rect	174	79	175	80
rect	174	80	175	81
rect	174	81	175	82
rect	174	82	175	83
rect	174	83	175	84
rect	174	84	175	85
rect	174	85	175	86
rect	174	86	175	87
rect	174	87	175	88
rect	174	88	175	89
rect	174	89	175	90
rect	174	90	175	91
rect	174	91	175	92
rect	174	92	175	93
rect	174	93	175	94
rect	174	94	175	95
rect	174	95	175	96
rect	174	96	175	97
rect	174	97	175	98
rect	174	98	175	99
rect	174	99	175	100
rect	174	100	175	101
rect	174	101	175	102
rect	174	102	175	103
rect	174	103	175	104
rect	174	104	175	105
rect	174	105	175	106
rect	174	106	175	107
rect	174	107	175	108
rect	174	108	175	109
rect	174	109	175	110
rect	174	110	175	111
rect	174	111	175	112
rect	174	112	175	113
rect	174	113	175	114
rect	174	114	175	115
rect	174	115	175	116
rect	174	116	175	117
rect	174	117	175	118
rect	174	118	175	119
rect	174	119	175	120
rect	174	120	175	121
rect	174	121	175	122
rect	174	122	175	123
rect	174	123	175	124
rect	174	124	175	125
rect	174	125	175	126
rect	174	126	175	127
rect	174	127	175	128
rect	174	128	175	129
rect	174	129	175	130
rect	174	130	175	131
rect	174	131	175	132
rect	174	132	175	133
rect	174	133	175	134
rect	174	134	175	135
rect	174	135	175	136
rect	174	136	175	137
rect	174	137	175	138
rect	174	138	175	139
rect	174	139	175	140
rect	174	140	175	141
rect	174	141	175	142
rect	174	142	175	143
rect	174	143	175	144
rect	174	144	175	145
rect	174	145	175	146
rect	174	146	175	147
rect	174	147	175	148
rect	174	148	175	149
rect	174	149	175	150
rect	174	150	175	151
rect	174	151	175	152
rect	174	152	175	153
rect	174	153	175	154
rect	174	154	175	155
rect	174	155	175	156
rect	174	156	175	157
rect	174	157	175	158
rect	174	158	175	159
rect	174	159	175	160
rect	174	160	175	161
rect	174	161	175	162
rect	174	162	175	163
rect	174	163	175	164
rect	174	164	175	165
rect	174	165	175	166
rect	174	166	175	167
rect	174	167	175	168
rect	174	168	175	169
rect	174	169	175	170
rect	174	170	175	171
rect	174	171	175	172
rect	174	172	175	173
rect	174	173	175	174
rect	174	174	175	175
rect	174	175	175	176
rect	174	176	175	177
rect	174	177	175	178
rect	174	178	175	179
rect	174	179	175	180
rect	174	180	175	181
rect	174	181	175	182
rect	174	182	175	183
rect	174	183	175	184
rect	174	184	175	185
rect	174	185	175	186
rect	174	186	175	187
rect	174	187	175	188
rect	174	188	175	189
rect	174	189	175	190
rect	174	190	175	191
rect	174	191	175	192
rect	174	192	175	193
rect	174	193	175	194
rect	174	194	175	195
rect	174	195	175	196
rect	174	196	175	197
rect	174	197	175	198
rect	174	198	175	199
rect	174	199	175	200
rect	174	200	175	201
rect	174	201	175	202
rect	174	202	175	203
rect	174	203	175	204
rect	174	204	175	205
rect	174	205	175	206
rect	174	206	175	207
rect	174	207	175	208
rect	174	208	175	209
rect	174	209	175	210
rect	174	210	175	211
rect	174	211	175	212
rect	174	212	175	213
rect	174	213	175	214
rect	174	214	175	215
rect	174	215	175	216
rect	174	216	175	217
rect	174	217	175	218
rect	174	218	175	219
rect	174	219	175	220
rect	174	220	175	221
rect	174	221	175	222
rect	174	222	175	223
rect	174	223	175	224
rect	174	224	175	225
rect	174	225	175	226
rect	174	226	175	227
rect	174	227	175	228
rect	174	228	175	229
rect	174	229	175	230
rect	174	230	175	231
rect	174	231	175	232
rect	174	232	175	233
rect	174	233	175	234
rect	174	234	175	235
rect	174	235	175	236
rect	174	236	175	237
rect	174	237	175	238
rect	174	238	175	239
rect	174	239	175	240
rect	174	240	175	241
rect	174	241	175	242
rect	174	242	175	243
rect	174	243	175	244
rect	174	244	175	245
rect	174	245	175	246
rect	174	246	175	247
rect	174	247	175	248
rect	174	248	175	249
rect	174	249	175	250
rect	174	250	175	251
rect	174	251	175	252
rect	174	252	175	253
rect	174	253	175	254
rect	174	254	175	255
rect	174	255	175	256
rect	174	256	175	257
rect	174	257	175	258
rect	174	258	175	259
rect	174	259	175	260
rect	174	260	175	261
rect	174	261	175	262
rect	174	262	175	263
rect	174	263	175	264
rect	174	264	175	265
rect	174	265	175	266
rect	174	266	175	267
rect	174	267	175	268
rect	174	268	175	269
rect	174	269	175	270
rect	174	270	175	271
rect	174	271	175	272
rect	174	272	175	273
rect	174	273	175	274
rect	174	274	175	275
rect	174	275	175	276
rect	174	276	175	277
rect	174	277	175	278
rect	174	278	175	279
rect	174	279	175	280
rect	174	280	175	281
rect	174	281	175	282
rect	174	282	175	283
rect	174	283	175	284
rect	174	284	175	285
rect	174	285	175	286
rect	174	286	175	287
rect	174	287	175	288
rect	174	288	175	289
rect	174	289	175	290
rect	174	290	175	291
rect	174	291	175	292
rect	174	292	175	293
rect	174	293	175	294
rect	174	294	175	295
rect	174	295	175	296
rect	174	296	175	297
rect	174	297	175	298
rect	174	298	175	299
rect	174	299	175	300
rect	174	300	175	301
rect	174	301	175	302
rect	174	302	175	303
rect	174	303	175	304
rect	174	304	175	305
rect	174	305	175	306
rect	174	306	175	307
rect	174	307	175	308
rect	174	308	175	309
rect	174	309	175	310
rect	174	310	175	311
rect	174	311	175	312
rect	174	312	175	313
rect	174	313	175	314
rect	174	314	175	315
rect	174	315	175	316
rect	174	316	175	317
rect	174	317	175	318
rect	174	318	175	319
rect	174	319	175	320
rect	174	320	175	321
rect	174	321	175	322
rect	174	322	175	323
rect	174	323	175	324
rect	174	324	175	325
rect	174	325	175	326
rect	174	326	175	327
rect	174	327	175	328
rect	174	328	175	329
rect	174	329	175	330
rect	175	0	176	1
rect	175	1	176	2
rect	175	2	176	3
rect	175	3	176	4
rect	175	4	176	5
rect	175	5	176	6
rect	175	6	176	7
rect	175	7	176	8
rect	175	8	176	9
rect	175	9	176	10
rect	175	10	176	11
rect	175	11	176	12
rect	175	12	176	13
rect	175	13	176	14
rect	175	14	176	15
rect	175	15	176	16
rect	175	16	176	17
rect	175	17	176	18
rect	175	18	176	19
rect	175	19	176	20
rect	175	20	176	21
rect	175	21	176	22
rect	175	22	176	23
rect	175	23	176	24
rect	175	24	176	25
rect	175	25	176	26
rect	175	26	176	27
rect	175	27	176	28
rect	175	28	176	29
rect	175	29	176	30
rect	175	30	176	31
rect	175	31	176	32
rect	175	32	176	33
rect	175	33	176	34
rect	175	34	176	35
rect	175	35	176	36
rect	175	36	176	37
rect	175	37	176	38
rect	175	38	176	39
rect	175	39	176	40
rect	175	40	176	41
rect	175	41	176	42
rect	175	42	176	43
rect	175	43	176	44
rect	175	44	176	45
rect	175	45	176	46
rect	175	46	176	47
rect	175	47	176	48
rect	175	48	176	49
rect	175	49	176	50
rect	175	50	176	51
rect	175	51	176	52
rect	175	52	176	53
rect	175	53	176	54
rect	175	54	176	55
rect	175	55	176	56
rect	175	56	176	57
rect	175	57	176	58
rect	175	58	176	59
rect	175	59	176	60
rect	175	60	176	61
rect	175	61	176	62
rect	175	62	176	63
rect	175	63	176	64
rect	175	64	176	65
rect	175	65	176	66
rect	175	66	176	67
rect	175	67	176	68
rect	175	68	176	69
rect	175	69	176	70
rect	175	70	176	71
rect	175	71	176	72
rect	175	72	176	73
rect	175	73	176	74
rect	175	74	176	75
rect	175	75	176	76
rect	175	76	176	77
rect	175	77	176	78
rect	175	78	176	79
rect	175	79	176	80
rect	175	80	176	81
rect	175	81	176	82
rect	175	82	176	83
rect	175	83	176	84
rect	175	84	176	85
rect	175	85	176	86
rect	175	86	176	87
rect	175	87	176	88
rect	175	88	176	89
rect	175	89	176	90
rect	175	90	176	91
rect	175	91	176	92
rect	175	92	176	93
rect	175	93	176	94
rect	175	94	176	95
rect	175	95	176	96
rect	175	96	176	97
rect	175	97	176	98
rect	175	98	176	99
rect	175	99	176	100
rect	175	100	176	101
rect	175	101	176	102
rect	175	102	176	103
rect	175	103	176	104
rect	175	104	176	105
rect	175	105	176	106
rect	175	106	176	107
rect	175	107	176	108
rect	175	108	176	109
rect	175	109	176	110
rect	175	110	176	111
rect	175	111	176	112
rect	175	112	176	113
rect	175	113	176	114
rect	175	114	176	115
rect	175	115	176	116
rect	175	116	176	117
rect	175	117	176	118
rect	175	118	176	119
rect	175	119	176	120
rect	175	120	176	121
rect	175	121	176	122
rect	175	122	176	123
rect	175	123	176	124
rect	175	124	176	125
rect	175	125	176	126
rect	175	126	176	127
rect	175	127	176	128
rect	175	128	176	129
rect	175	129	176	130
rect	175	130	176	131
rect	175	131	176	132
rect	175	132	176	133
rect	175	133	176	134
rect	175	134	176	135
rect	175	135	176	136
rect	175	136	176	137
rect	175	137	176	138
rect	175	138	176	139
rect	175	139	176	140
rect	175	140	176	141
rect	175	141	176	142
rect	175	142	176	143
rect	175	143	176	144
rect	175	144	176	145
rect	175	145	176	146
rect	175	146	176	147
rect	175	147	176	148
rect	175	148	176	149
rect	175	149	176	150
rect	175	150	176	151
rect	175	151	176	152
rect	175	152	176	153
rect	175	153	176	154
rect	175	154	176	155
rect	175	155	176	156
rect	175	156	176	157
rect	175	157	176	158
rect	175	158	176	159
rect	175	159	176	160
rect	175	160	176	161
rect	175	161	176	162
rect	175	162	176	163
rect	175	163	176	164
rect	175	164	176	165
rect	175	165	176	166
rect	175	166	176	167
rect	175	167	176	168
rect	175	168	176	169
rect	175	169	176	170
rect	175	170	176	171
rect	175	171	176	172
rect	175	172	176	173
rect	175	173	176	174
rect	175	174	176	175
rect	175	175	176	176
rect	175	176	176	177
rect	175	177	176	178
rect	175	178	176	179
rect	175	179	176	180
rect	175	180	176	181
rect	175	181	176	182
rect	175	182	176	183
rect	175	183	176	184
rect	175	184	176	185
rect	175	185	176	186
rect	175	186	176	187
rect	175	187	176	188
rect	175	188	176	189
rect	175	189	176	190
rect	175	190	176	191
rect	175	191	176	192
rect	175	192	176	193
rect	175	193	176	194
rect	175	194	176	195
rect	175	195	176	196
rect	175	196	176	197
rect	175	197	176	198
rect	175	198	176	199
rect	175	199	176	200
rect	175	200	176	201
rect	175	201	176	202
rect	175	202	176	203
rect	175	203	176	204
rect	175	204	176	205
rect	175	205	176	206
rect	175	206	176	207
rect	175	207	176	208
rect	175	208	176	209
rect	175	209	176	210
rect	175	210	176	211
rect	175	211	176	212
rect	175	212	176	213
rect	175	213	176	214
rect	175	214	176	215
rect	175	215	176	216
rect	175	216	176	217
rect	175	217	176	218
rect	175	218	176	219
rect	175	219	176	220
rect	175	220	176	221
rect	175	221	176	222
rect	175	222	176	223
rect	175	223	176	224
rect	175	224	176	225
rect	175	225	176	226
rect	175	226	176	227
rect	175	227	176	228
rect	175	228	176	229
rect	175	229	176	230
rect	175	230	176	231
rect	175	231	176	232
rect	175	232	176	233
rect	175	233	176	234
rect	175	234	176	235
rect	175	235	176	236
rect	175	236	176	237
rect	175	237	176	238
rect	175	238	176	239
rect	175	239	176	240
rect	175	240	176	241
rect	175	241	176	242
rect	175	242	176	243
rect	175	243	176	244
rect	175	244	176	245
rect	175	245	176	246
rect	175	246	176	247
rect	175	247	176	248
rect	175	248	176	249
rect	175	249	176	250
rect	175	250	176	251
rect	175	251	176	252
rect	175	252	176	253
rect	175	253	176	254
rect	175	254	176	255
rect	175	255	176	256
rect	175	256	176	257
rect	175	257	176	258
rect	175	258	176	259
rect	175	259	176	260
rect	175	260	176	261
rect	175	261	176	262
rect	175	262	176	263
rect	175	263	176	264
rect	175	264	176	265
rect	175	265	176	266
rect	175	266	176	267
rect	175	267	176	268
rect	175	268	176	269
rect	175	269	176	270
rect	175	270	176	271
rect	175	271	176	272
rect	175	272	176	273
rect	175	273	176	274
rect	175	274	176	275
rect	175	275	176	276
rect	175	276	176	277
rect	175	277	176	278
rect	175	278	176	279
rect	175	279	176	280
rect	175	280	176	281
rect	175	281	176	282
rect	175	282	176	283
rect	175	283	176	284
rect	175	284	176	285
rect	175	285	176	286
rect	175	286	176	287
rect	175	287	176	288
rect	175	288	176	289
rect	175	289	176	290
rect	175	290	176	291
rect	175	291	176	292
rect	175	292	176	293
rect	175	293	176	294
rect	175	294	176	295
rect	175	295	176	296
rect	175	296	176	297
rect	175	297	176	298
rect	175	298	176	299
rect	175	299	176	300
rect	175	300	176	301
rect	175	301	176	302
rect	175	302	176	303
rect	175	303	176	304
rect	175	304	176	305
rect	175	305	176	306
rect	175	306	176	307
rect	175	307	176	308
rect	175	308	176	309
rect	175	309	176	310
rect	175	310	176	311
rect	175	311	176	312
rect	175	312	176	313
rect	175	313	176	314
rect	175	314	176	315
rect	175	315	176	316
rect	175	316	176	317
rect	175	317	176	318
rect	175	318	176	319
rect	175	319	176	320
rect	175	320	176	321
rect	175	321	176	322
rect	175	322	176	323
rect	175	323	176	324
rect	175	324	176	325
rect	175	325	176	326
rect	175	326	176	327
rect	175	327	176	328
rect	175	328	176	329
rect	175	329	176	330
rect	176	0	177	1
rect	176	1	177	2
rect	176	2	177	3
rect	176	3	177	4
rect	176	4	177	5
rect	176	5	177	6
rect	176	6	177	7
rect	176	7	177	8
rect	176	8	177	9
rect	176	9	177	10
rect	176	10	177	11
rect	176	11	177	12
rect	176	12	177	13
rect	176	13	177	14
rect	176	14	177	15
rect	176	15	177	16
rect	176	16	177	17
rect	176	17	177	18
rect	176	18	177	19
rect	176	19	177	20
rect	176	20	177	21
rect	176	21	177	22
rect	176	22	177	23
rect	176	23	177	24
rect	176	24	177	25
rect	176	25	177	26
rect	176	26	177	27
rect	176	27	177	28
rect	176	28	177	29
rect	176	29	177	30
rect	176	30	177	31
rect	176	31	177	32
rect	176	32	177	33
rect	176	33	177	34
rect	176	34	177	35
rect	176	35	177	36
rect	176	36	177	37
rect	176	37	177	38
rect	176	38	177	39
rect	176	39	177	40
rect	176	40	177	41
rect	176	41	177	42
rect	176	42	177	43
rect	176	43	177	44
rect	176	44	177	45
rect	176	45	177	46
rect	176	46	177	47
rect	176	47	177	48
rect	176	48	177	49
rect	176	49	177	50
rect	176	50	177	51
rect	176	51	177	52
rect	176	52	177	53
rect	176	53	177	54
rect	176	54	177	55
rect	176	55	177	56
rect	176	56	177	57
rect	176	57	177	58
rect	176	58	177	59
rect	176	59	177	60
rect	176	60	177	61
rect	176	61	177	62
rect	176	62	177	63
rect	176	63	177	64
rect	176	64	177	65
rect	176	65	177	66
rect	176	66	177	67
rect	176	67	177	68
rect	176	68	177	69
rect	176	69	177	70
rect	176	70	177	71
rect	176	71	177	72
rect	176	72	177	73
rect	176	73	177	74
rect	176	74	177	75
rect	176	75	177	76
rect	176	76	177	77
rect	176	77	177	78
rect	176	78	177	79
rect	176	79	177	80
rect	176	80	177	81
rect	176	81	177	82
rect	176	82	177	83
rect	176	83	177	84
rect	176	84	177	85
rect	176	85	177	86
rect	176	86	177	87
rect	176	87	177	88
rect	176	88	177	89
rect	176	89	177	90
rect	176	90	177	91
rect	176	91	177	92
rect	176	92	177	93
rect	176	93	177	94
rect	176	94	177	95
rect	176	95	177	96
rect	176	96	177	97
rect	176	97	177	98
rect	176	98	177	99
rect	176	99	177	100
rect	176	100	177	101
rect	176	101	177	102
rect	176	102	177	103
rect	176	103	177	104
rect	176	104	177	105
rect	176	105	177	106
rect	176	106	177	107
rect	176	107	177	108
rect	176	108	177	109
rect	176	109	177	110
rect	176	110	177	111
rect	176	111	177	112
rect	176	112	177	113
rect	176	113	177	114
rect	176	114	177	115
rect	176	115	177	116
rect	176	116	177	117
rect	176	117	177	118
rect	176	118	177	119
rect	176	119	177	120
rect	176	120	177	121
rect	176	121	177	122
rect	176	122	177	123
rect	176	123	177	124
rect	176	124	177	125
rect	176	125	177	126
rect	176	126	177	127
rect	176	127	177	128
rect	176	128	177	129
rect	176	129	177	130
rect	176	130	177	131
rect	176	131	177	132
rect	176	132	177	133
rect	176	133	177	134
rect	176	134	177	135
rect	176	135	177	136
rect	176	136	177	137
rect	176	137	177	138
rect	176	138	177	139
rect	176	139	177	140
rect	176	140	177	141
rect	176	141	177	142
rect	176	142	177	143
rect	176	143	177	144
rect	176	144	177	145
rect	176	145	177	146
rect	176	146	177	147
rect	176	147	177	148
rect	176	148	177	149
rect	176	149	177	150
rect	176	150	177	151
rect	176	151	177	152
rect	176	152	177	153
rect	176	153	177	154
rect	176	154	177	155
rect	176	155	177	156
rect	176	156	177	157
rect	176	157	177	158
rect	176	158	177	159
rect	176	159	177	160
rect	176	160	177	161
rect	176	161	177	162
rect	176	162	177	163
rect	176	163	177	164
rect	176	164	177	165
rect	176	165	177	166
rect	176	166	177	167
rect	176	167	177	168
rect	176	168	177	169
rect	176	169	177	170
rect	176	170	177	171
rect	176	171	177	172
rect	176	172	177	173
rect	176	173	177	174
rect	176	174	177	175
rect	176	175	177	176
rect	176	176	177	177
rect	176	177	177	178
rect	176	178	177	179
rect	176	179	177	180
rect	176	180	177	181
rect	176	181	177	182
rect	176	182	177	183
rect	176	183	177	184
rect	176	184	177	185
rect	176	185	177	186
rect	176	186	177	187
rect	176	187	177	188
rect	176	188	177	189
rect	176	189	177	190
rect	176	190	177	191
rect	176	191	177	192
rect	176	192	177	193
rect	176	193	177	194
rect	176	194	177	195
rect	176	195	177	196
rect	176	196	177	197
rect	176	197	177	198
rect	176	198	177	199
rect	176	199	177	200
rect	176	200	177	201
rect	176	201	177	202
rect	176	202	177	203
rect	176	203	177	204
rect	176	204	177	205
rect	176	205	177	206
rect	176	206	177	207
rect	176	207	177	208
rect	176	208	177	209
rect	176	209	177	210
rect	176	210	177	211
rect	176	211	177	212
rect	176	212	177	213
rect	176	213	177	214
rect	176	214	177	215
rect	176	215	177	216
rect	176	216	177	217
rect	176	217	177	218
rect	176	218	177	219
rect	176	219	177	220
rect	176	220	177	221
rect	176	221	177	222
rect	176	222	177	223
rect	176	223	177	224
rect	176	224	177	225
rect	176	225	177	226
rect	176	226	177	227
rect	176	227	177	228
rect	176	228	177	229
rect	176	229	177	230
rect	176	230	177	231
rect	176	231	177	232
rect	176	232	177	233
rect	176	233	177	234
rect	176	234	177	235
rect	176	235	177	236
rect	176	236	177	237
rect	176	237	177	238
rect	176	238	177	239
rect	176	239	177	240
rect	176	240	177	241
rect	176	241	177	242
rect	176	242	177	243
rect	176	243	177	244
rect	176	244	177	245
rect	176	245	177	246
rect	176	246	177	247
rect	176	247	177	248
rect	176	248	177	249
rect	176	249	177	250
rect	176	250	177	251
rect	176	251	177	252
rect	176	252	177	253
rect	176	253	177	254
rect	176	254	177	255
rect	176	255	177	256
rect	176	256	177	257
rect	176	257	177	258
rect	176	258	177	259
rect	176	259	177	260
rect	176	260	177	261
rect	176	261	177	262
rect	176	262	177	263
rect	176	263	177	264
rect	176	264	177	265
rect	176	265	177	266
rect	176	266	177	267
rect	176	267	177	268
rect	176	268	177	269
rect	176	269	177	270
rect	176	270	177	271
rect	176	271	177	272
rect	176	272	177	273
rect	176	273	177	274
rect	176	274	177	275
rect	176	275	177	276
rect	176	276	177	277
rect	176	277	177	278
rect	176	278	177	279
rect	176	279	177	280
rect	176	280	177	281
rect	176	281	177	282
rect	176	282	177	283
rect	176	283	177	284
rect	176	284	177	285
rect	176	285	177	286
rect	176	286	177	287
rect	176	287	177	288
rect	176	288	177	289
rect	176	289	177	290
rect	176	290	177	291
rect	176	291	177	292
rect	176	292	177	293
rect	176	293	177	294
rect	176	294	177	295
rect	176	295	177	296
rect	176	296	177	297
rect	176	297	177	298
rect	176	298	177	299
rect	176	299	177	300
rect	176	300	177	301
rect	176	301	177	302
rect	176	302	177	303
rect	176	303	177	304
rect	176	304	177	305
rect	176	305	177	306
rect	176	306	177	307
rect	176	307	177	308
rect	176	308	177	309
rect	176	309	177	310
rect	176	310	177	311
rect	176	311	177	312
rect	176	312	177	313
rect	176	313	177	314
rect	176	314	177	315
rect	176	315	177	316
rect	176	316	177	317
rect	176	317	177	318
rect	176	318	177	319
rect	176	319	177	320
rect	176	320	177	321
rect	176	321	177	322
rect	176	322	177	323
rect	176	323	177	324
rect	176	324	177	325
rect	176	325	177	326
rect	176	326	177	327
rect	176	327	177	328
rect	176	328	177	329
rect	176	329	177	330
rect	177	0	178	1
rect	177	1	178	2
rect	177	2	178	3
rect	177	3	178	4
rect	177	4	178	5
rect	177	5	178	6
rect	177	6	178	7
rect	177	7	178	8
rect	177	8	178	9
rect	177	9	178	10
rect	177	10	178	11
rect	177	11	178	12
rect	177	12	178	13
rect	177	13	178	14
rect	177	14	178	15
rect	177	15	178	16
rect	177	16	178	17
rect	177	17	178	18
rect	177	18	178	19
rect	177	19	178	20
rect	177	20	178	21
rect	177	21	178	22
rect	177	22	178	23
rect	177	23	178	24
rect	177	24	178	25
rect	177	25	178	26
rect	177	26	178	27
rect	177	27	178	28
rect	177	28	178	29
rect	177	29	178	30
rect	177	30	178	31
rect	177	31	178	32
rect	177	32	178	33
rect	177	33	178	34
rect	177	34	178	35
rect	177	35	178	36
rect	177	36	178	37
rect	177	37	178	38
rect	177	38	178	39
rect	177	39	178	40
rect	177	40	178	41
rect	177	41	178	42
rect	177	42	178	43
rect	177	43	178	44
rect	177	44	178	45
rect	177	45	178	46
rect	177	46	178	47
rect	177	47	178	48
rect	177	48	178	49
rect	177	49	178	50
rect	177	50	178	51
rect	177	51	178	52
rect	177	52	178	53
rect	177	53	178	54
rect	177	54	178	55
rect	177	55	178	56
rect	177	56	178	57
rect	177	57	178	58
rect	177	58	178	59
rect	177	59	178	60
rect	177	60	178	61
rect	177	61	178	62
rect	177	62	178	63
rect	177	63	178	64
rect	177	64	178	65
rect	177	65	178	66
rect	177	66	178	67
rect	177	67	178	68
rect	177	68	178	69
rect	177	69	178	70
rect	177	70	178	71
rect	177	71	178	72
rect	177	72	178	73
rect	177	73	178	74
rect	177	74	178	75
rect	177	75	178	76
rect	177	76	178	77
rect	177	77	178	78
rect	177	78	178	79
rect	177	79	178	80
rect	177	80	178	81
rect	177	81	178	82
rect	177	82	178	83
rect	177	83	178	84
rect	177	84	178	85
rect	177	85	178	86
rect	177	86	178	87
rect	177	87	178	88
rect	177	88	178	89
rect	177	89	178	90
rect	177	90	178	91
rect	177	91	178	92
rect	177	92	178	93
rect	177	93	178	94
rect	177	94	178	95
rect	177	95	178	96
rect	177	96	178	97
rect	177	97	178	98
rect	177	98	178	99
rect	177	99	178	100
rect	177	100	178	101
rect	177	101	178	102
rect	177	102	178	103
rect	177	103	178	104
rect	177	104	178	105
rect	177	105	178	106
rect	177	106	178	107
rect	177	107	178	108
rect	177	108	178	109
rect	177	109	178	110
rect	177	110	178	111
rect	177	111	178	112
rect	177	112	178	113
rect	177	113	178	114
rect	177	114	178	115
rect	177	115	178	116
rect	177	116	178	117
rect	177	117	178	118
rect	177	118	178	119
rect	177	119	178	120
rect	177	120	178	121
rect	177	121	178	122
rect	177	122	178	123
rect	177	123	178	124
rect	177	124	178	125
rect	177	125	178	126
rect	177	126	178	127
rect	177	127	178	128
rect	177	128	178	129
rect	177	129	178	130
rect	177	130	178	131
rect	177	131	178	132
rect	177	132	178	133
rect	177	133	178	134
rect	177	134	178	135
rect	177	135	178	136
rect	177	136	178	137
rect	177	137	178	138
rect	177	138	178	139
rect	177	139	178	140
rect	177	140	178	141
rect	177	141	178	142
rect	177	142	178	143
rect	177	143	178	144
rect	177	144	178	145
rect	177	145	178	146
rect	177	146	178	147
rect	177	147	178	148
rect	177	148	178	149
rect	177	149	178	150
rect	177	150	178	151
rect	177	151	178	152
rect	177	152	178	153
rect	177	153	178	154
rect	177	154	178	155
rect	177	155	178	156
rect	177	156	178	157
rect	177	157	178	158
rect	177	158	178	159
rect	177	159	178	160
rect	177	160	178	161
rect	177	161	178	162
rect	177	162	178	163
rect	177	163	178	164
rect	177	164	178	165
rect	177	165	178	166
rect	177	166	178	167
rect	177	167	178	168
rect	177	168	178	169
rect	177	169	178	170
rect	177	170	178	171
rect	177	171	178	172
rect	177	172	178	173
rect	177	173	178	174
rect	177	174	178	175
rect	177	175	178	176
rect	177	176	178	177
rect	177	177	178	178
rect	177	178	178	179
rect	177	179	178	180
rect	177	180	178	181
rect	177	181	178	182
rect	177	182	178	183
rect	177	183	178	184
rect	177	184	178	185
rect	177	185	178	186
rect	177	186	178	187
rect	177	187	178	188
rect	177	188	178	189
rect	177	189	178	190
rect	177	190	178	191
rect	177	191	178	192
rect	177	192	178	193
rect	177	193	178	194
rect	177	194	178	195
rect	177	195	178	196
rect	177	196	178	197
rect	177	197	178	198
rect	177	198	178	199
rect	177	199	178	200
rect	177	200	178	201
rect	177	201	178	202
rect	177	202	178	203
rect	177	203	178	204
rect	177	204	178	205
rect	177	205	178	206
rect	177	206	178	207
rect	177	207	178	208
rect	177	208	178	209
rect	177	209	178	210
rect	177	210	178	211
rect	177	211	178	212
rect	177	212	178	213
rect	177	213	178	214
rect	177	214	178	215
rect	177	215	178	216
rect	177	216	178	217
rect	177	217	178	218
rect	177	218	178	219
rect	177	219	178	220
rect	177	220	178	221
rect	177	221	178	222
rect	177	222	178	223
rect	177	223	178	224
rect	177	224	178	225
rect	177	225	178	226
rect	177	226	178	227
rect	177	227	178	228
rect	177	228	178	229
rect	177	229	178	230
rect	177	230	178	231
rect	177	231	178	232
rect	177	232	178	233
rect	177	233	178	234
rect	177	234	178	235
rect	177	235	178	236
rect	177	236	178	237
rect	177	237	178	238
rect	177	238	178	239
rect	177	239	178	240
rect	177	240	178	241
rect	177	241	178	242
rect	177	242	178	243
rect	177	243	178	244
rect	177	244	178	245
rect	177	245	178	246
rect	177	246	178	247
rect	177	247	178	248
rect	177	248	178	249
rect	177	249	178	250
rect	177	250	178	251
rect	177	251	178	252
rect	177	252	178	253
rect	177	253	178	254
rect	177	254	178	255
rect	177	255	178	256
rect	177	256	178	257
rect	177	257	178	258
rect	177	258	178	259
rect	177	259	178	260
rect	177	260	178	261
rect	177	261	178	262
rect	177	262	178	263
rect	177	263	178	264
rect	177	264	178	265
rect	177	265	178	266
rect	177	266	178	267
rect	177	267	178	268
rect	177	268	178	269
rect	177	269	178	270
rect	177	270	178	271
rect	177	271	178	272
rect	177	272	178	273
rect	177	273	178	274
rect	177	274	178	275
rect	177	275	178	276
rect	177	276	178	277
rect	177	277	178	278
rect	177	278	178	279
rect	177	279	178	280
rect	177	280	178	281
rect	177	281	178	282
rect	177	282	178	283
rect	177	283	178	284
rect	177	284	178	285
rect	177	285	178	286
rect	177	286	178	287
rect	177	287	178	288
rect	177	288	178	289
rect	177	289	178	290
rect	177	290	178	291
rect	177	291	178	292
rect	177	292	178	293
rect	177	293	178	294
rect	177	294	178	295
rect	177	295	178	296
rect	177	296	178	297
rect	177	297	178	298
rect	177	298	178	299
rect	177	299	178	300
rect	177	300	178	301
rect	177	301	178	302
rect	177	302	178	303
rect	177	303	178	304
rect	177	304	178	305
rect	177	305	178	306
rect	177	306	178	307
rect	177	307	178	308
rect	177	308	178	309
rect	177	309	178	310
rect	177	310	178	311
rect	177	311	178	312
rect	177	312	178	313
rect	177	313	178	314
rect	177	314	178	315
rect	177	315	178	316
rect	177	316	178	317
rect	177	317	178	318
rect	177	318	178	319
rect	177	319	178	320
rect	177	320	178	321
rect	177	321	178	322
rect	177	322	178	323
rect	177	323	178	324
rect	177	324	178	325
rect	177	325	178	326
rect	177	326	178	327
rect	177	327	178	328
rect	177	328	178	329
rect	177	329	178	330
rect	197	0	198	1
rect	197	1	198	2
rect	197	2	198	3
rect	197	3	198	4
rect	197	4	198	5
rect	197	5	198	6
rect	197	6	198	7
rect	197	7	198	8
rect	197	8	198	9
rect	197	9	198	10
rect	197	10	198	11
rect	197	11	198	12
rect	197	12	198	13
rect	197	13	198	14
rect	197	14	198	15
rect	197	15	198	16
rect	197	16	198	17
rect	197	17	198	18
rect	197	18	198	19
rect	197	19	198	20
rect	197	20	198	21
rect	197	21	198	22
rect	197	22	198	23
rect	197	23	198	24
rect	197	24	198	25
rect	197	25	198	26
rect	197	26	198	27
rect	197	27	198	28
rect	197	28	198	29
rect	197	29	198	30
rect	197	30	198	31
rect	197	31	198	32
rect	197	32	198	33
rect	197	33	198	34
rect	197	34	198	35
rect	197	35	198	36
rect	197	36	198	37
rect	197	37	198	38
rect	197	38	198	39
rect	197	39	198	40
rect	197	40	198	41
rect	197	41	198	42
rect	197	42	198	43
rect	197	43	198	44
rect	197	44	198	45
rect	197	45	198	46
rect	197	46	198	47
rect	197	47	198	48
rect	197	48	198	49
rect	197	49	198	50
rect	197	50	198	51
rect	197	51	198	52
rect	197	52	198	53
rect	197	53	198	54
rect	197	54	198	55
rect	197	55	198	56
rect	197	56	198	57
rect	197	57	198	58
rect	197	58	198	59
rect	197	59	198	60
rect	197	60	198	61
rect	197	61	198	62
rect	197	62	198	63
rect	197	63	198	64
rect	197	64	198	65
rect	197	65	198	66
rect	197	66	198	67
rect	197	67	198	68
rect	197	68	198	69
rect	197	69	198	70
rect	197	70	198	71
rect	197	71	198	72
rect	197	72	198	73
rect	197	73	198	74
rect	197	74	198	75
rect	197	75	198	76
rect	197	76	198	77
rect	197	77	198	78
rect	197	78	198	79
rect	197	79	198	80
rect	197	80	198	81
rect	197	81	198	82
rect	197	82	198	83
rect	197	83	198	84
rect	197	84	198	85
rect	197	85	198	86
rect	197	86	198	87
rect	197	87	198	88
rect	197	88	198	89
rect	197	89	198	90
rect	197	90	198	91
rect	197	91	198	92
rect	197	92	198	93
rect	197	93	198	94
rect	197	94	198	95
rect	197	95	198	96
rect	197	96	198	97
rect	197	97	198	98
rect	197	98	198	99
rect	197	99	198	100
rect	197	100	198	101
rect	197	101	198	102
rect	197	102	198	103
rect	197	103	198	104
rect	197	104	198	105
rect	197	105	198	106
rect	197	106	198	107
rect	197	107	198	108
rect	197	108	198	109
rect	197	109	198	110
rect	197	110	198	111
rect	197	111	198	112
rect	197	112	198	113
rect	197	113	198	114
rect	197	114	198	115
rect	197	115	198	116
rect	197	116	198	117
rect	197	117	198	118
rect	197	118	198	119
rect	197	119	198	120
rect	197	120	198	121
rect	197	121	198	122
rect	197	122	198	123
rect	197	123	198	124
rect	197	124	198	125
rect	197	125	198	126
rect	197	126	198	127
rect	197	127	198	128
rect	197	128	198	129
rect	197	129	198	130
rect	197	130	198	131
rect	197	131	198	132
rect	197	132	198	133
rect	197	133	198	134
rect	197	134	198	135
rect	197	135	198	136
rect	197	136	198	137
rect	197	137	198	138
rect	197	138	198	139
rect	197	139	198	140
rect	197	140	198	141
rect	197	141	198	142
rect	197	142	198	143
rect	197	143	198	144
rect	197	144	198	145
rect	197	145	198	146
rect	197	146	198	147
rect	197	147	198	148
rect	197	148	198	149
rect	197	149	198	150
rect	197	150	198	151
rect	197	151	198	152
rect	197	152	198	153
rect	197	153	198	154
rect	197	154	198	155
rect	197	155	198	156
rect	197	156	198	157
rect	197	157	198	158
rect	197	158	198	159
rect	197	159	198	160
rect	197	160	198	161
rect	197	161	198	162
rect	197	162	198	163
rect	197	163	198	164
rect	197	164	198	165
rect	197	165	198	166
rect	197	166	198	167
rect	197	167	198	168
rect	197	168	198	169
rect	197	169	198	170
rect	197	170	198	171
rect	197	171	198	172
rect	197	172	198	173
rect	197	173	198	174
rect	197	174	198	175
rect	197	175	198	176
rect	197	176	198	177
rect	197	177	198	178
rect	197	178	198	179
rect	197	179	198	180
rect	197	180	198	181
rect	197	181	198	182
rect	197	182	198	183
rect	197	183	198	184
rect	197	184	198	185
rect	197	185	198	186
rect	197	186	198	187
rect	197	187	198	188
rect	197	188	198	189
rect	197	189	198	190
rect	197	190	198	191
rect	197	191	198	192
rect	197	192	198	193
rect	197	193	198	194
rect	197	194	198	195
rect	197	195	198	196
rect	197	196	198	197
rect	197	197	198	198
rect	197	198	198	199
rect	197	199	198	200
rect	197	200	198	201
rect	197	201	198	202
rect	197	202	198	203
rect	197	203	198	204
rect	197	204	198	205
rect	197	205	198	206
rect	197	206	198	207
rect	197	207	198	208
rect	197	208	198	209
rect	197	209	198	210
rect	197	210	198	211
rect	197	211	198	212
rect	197	212	198	213
rect	197	213	198	214
rect	197	214	198	215
rect	197	215	198	216
rect	197	216	198	217
rect	197	217	198	218
rect	197	218	198	219
rect	197	219	198	220
rect	197	220	198	221
rect	197	221	198	222
rect	197	222	198	223
rect	197	223	198	224
rect	197	224	198	225
rect	197	225	198	226
rect	197	226	198	227
rect	197	227	198	228
rect	197	228	198	229
rect	197	229	198	230
rect	197	230	198	231
rect	197	231	198	232
rect	197	232	198	233
rect	197	233	198	234
rect	197	234	198	235
rect	197	235	198	236
rect	197	236	198	237
rect	197	237	198	238
rect	197	238	198	239
rect	197	239	198	240
rect	197	240	198	241
rect	197	241	198	242
rect	197	242	198	243
rect	197	243	198	244
rect	197	244	198	245
rect	197	245	198	246
rect	197	246	198	247
rect	197	247	198	248
rect	197	248	198	249
rect	197	249	198	250
rect	197	250	198	251
rect	197	251	198	252
rect	197	252	198	253
rect	197	253	198	254
rect	197	254	198	255
rect	197	255	198	256
rect	197	256	198	257
rect	197	257	198	258
rect	197	258	198	259
rect	197	259	198	260
rect	197	260	198	261
rect	197	261	198	262
rect	197	262	198	263
rect	197	263	198	264
rect	197	264	198	265
rect	197	265	198	266
rect	197	266	198	267
rect	197	267	198	268
rect	197	268	198	269
rect	197	269	198	270
rect	197	270	198	271
rect	197	271	198	272
rect	197	272	198	273
rect	197	273	198	274
rect	197	274	198	275
rect	197	275	198	276
rect	197	276	198	277
rect	197	277	198	278
rect	197	278	198	279
rect	197	279	198	280
rect	197	280	198	281
rect	197	281	198	282
rect	197	282	198	283
rect	197	283	198	284
rect	197	284	198	285
rect	197	285	198	286
rect	197	286	198	287
rect	197	287	198	288
rect	197	288	198	289
rect	197	289	198	290
rect	197	290	198	291
rect	197	291	198	292
rect	197	292	198	293
rect	197	293	198	294
rect	197	294	198	295
rect	197	295	198	296
rect	197	296	198	297
rect	197	297	198	298
rect	197	298	198	299
rect	197	299	198	300
rect	197	300	198	301
rect	197	301	198	302
rect	197	302	198	303
rect	197	303	198	304
rect	197	304	198	305
rect	197	305	198	306
rect	197	306	198	307
rect	197	307	198	308
rect	197	308	198	309
rect	197	309	198	310
rect	197	310	198	311
rect	197	311	198	312
rect	197	312	198	313
rect	197	313	198	314
rect	197	314	198	315
rect	197	315	198	316
rect	197	316	198	317
rect	197	317	198	318
rect	197	318	198	319
rect	197	319	198	320
rect	197	320	198	321
rect	197	321	198	322
rect	197	322	198	323
rect	197	323	198	324
rect	197	324	198	325
rect	197	325	198	326
rect	197	326	198	327
rect	197	327	198	328
rect	197	328	198	329
rect	197	329	198	330
rect	197	330	198	331
rect	197	331	198	332
rect	197	332	198	333
rect	197	333	198	334
rect	197	334	198	335
rect	197	335	198	336
rect	198	0	199	1
rect	198	1	199	2
rect	198	2	199	3
rect	198	3	199	4
rect	198	4	199	5
rect	198	5	199	6
rect	198	6	199	7
rect	198	7	199	8
rect	198	8	199	9
rect	198	9	199	10
rect	198	10	199	11
rect	198	11	199	12
rect	198	12	199	13
rect	198	13	199	14
rect	198	14	199	15
rect	198	15	199	16
rect	198	16	199	17
rect	198	17	199	18
rect	198	18	199	19
rect	198	19	199	20
rect	198	20	199	21
rect	198	21	199	22
rect	198	22	199	23
rect	198	23	199	24
rect	198	24	199	25
rect	198	25	199	26
rect	198	26	199	27
rect	198	27	199	28
rect	198	28	199	29
rect	198	29	199	30
rect	198	30	199	31
rect	198	31	199	32
rect	198	32	199	33
rect	198	33	199	34
rect	198	34	199	35
rect	198	35	199	36
rect	198	36	199	37
rect	198	37	199	38
rect	198	38	199	39
rect	198	39	199	40
rect	198	40	199	41
rect	198	41	199	42
rect	198	42	199	43
rect	198	43	199	44
rect	198	44	199	45
rect	198	45	199	46
rect	198	46	199	47
rect	198	47	199	48
rect	198	48	199	49
rect	198	49	199	50
rect	198	50	199	51
rect	198	51	199	52
rect	198	52	199	53
rect	198	53	199	54
rect	198	54	199	55
rect	198	55	199	56
rect	198	56	199	57
rect	198	57	199	58
rect	198	58	199	59
rect	198	59	199	60
rect	198	60	199	61
rect	198	61	199	62
rect	198	62	199	63
rect	198	63	199	64
rect	198	64	199	65
rect	198	65	199	66
rect	198	66	199	67
rect	198	67	199	68
rect	198	68	199	69
rect	198	69	199	70
rect	198	70	199	71
rect	198	71	199	72
rect	198	72	199	73
rect	198	73	199	74
rect	198	74	199	75
rect	198	75	199	76
rect	198	76	199	77
rect	198	77	199	78
rect	198	78	199	79
rect	198	79	199	80
rect	198	80	199	81
rect	198	81	199	82
rect	198	82	199	83
rect	198	83	199	84
rect	198	84	199	85
rect	198	85	199	86
rect	198	86	199	87
rect	198	87	199	88
rect	198	88	199	89
rect	198	89	199	90
rect	198	90	199	91
rect	198	91	199	92
rect	198	92	199	93
rect	198	93	199	94
rect	198	94	199	95
rect	198	95	199	96
rect	198	96	199	97
rect	198	97	199	98
rect	198	98	199	99
rect	198	99	199	100
rect	198	100	199	101
rect	198	101	199	102
rect	198	102	199	103
rect	198	103	199	104
rect	198	104	199	105
rect	198	105	199	106
rect	198	106	199	107
rect	198	107	199	108
rect	198	108	199	109
rect	198	109	199	110
rect	198	110	199	111
rect	198	111	199	112
rect	198	112	199	113
rect	198	113	199	114
rect	198	114	199	115
rect	198	115	199	116
rect	198	116	199	117
rect	198	117	199	118
rect	198	118	199	119
rect	198	119	199	120
rect	198	120	199	121
rect	198	121	199	122
rect	198	122	199	123
rect	198	123	199	124
rect	198	124	199	125
rect	198	125	199	126
rect	198	126	199	127
rect	198	127	199	128
rect	198	128	199	129
rect	198	129	199	130
rect	198	130	199	131
rect	198	131	199	132
rect	198	132	199	133
rect	198	133	199	134
rect	198	134	199	135
rect	198	135	199	136
rect	198	136	199	137
rect	198	137	199	138
rect	198	138	199	139
rect	198	139	199	140
rect	198	140	199	141
rect	198	141	199	142
rect	198	142	199	143
rect	198	143	199	144
rect	198	144	199	145
rect	198	145	199	146
rect	198	146	199	147
rect	198	147	199	148
rect	198	148	199	149
rect	198	149	199	150
rect	198	150	199	151
rect	198	151	199	152
rect	198	152	199	153
rect	198	153	199	154
rect	198	154	199	155
rect	198	155	199	156
rect	198	156	199	157
rect	198	157	199	158
rect	198	158	199	159
rect	198	159	199	160
rect	198	160	199	161
rect	198	161	199	162
rect	198	162	199	163
rect	198	163	199	164
rect	198	164	199	165
rect	198	165	199	166
rect	198	166	199	167
rect	198	167	199	168
rect	198	168	199	169
rect	198	169	199	170
rect	198	170	199	171
rect	198	171	199	172
rect	198	172	199	173
rect	198	173	199	174
rect	198	174	199	175
rect	198	175	199	176
rect	198	176	199	177
rect	198	177	199	178
rect	198	178	199	179
rect	198	179	199	180
rect	198	180	199	181
rect	198	181	199	182
rect	198	182	199	183
rect	198	183	199	184
rect	198	184	199	185
rect	198	185	199	186
rect	198	186	199	187
rect	198	187	199	188
rect	198	188	199	189
rect	198	189	199	190
rect	198	190	199	191
rect	198	191	199	192
rect	198	192	199	193
rect	198	193	199	194
rect	198	194	199	195
rect	198	195	199	196
rect	198	196	199	197
rect	198	197	199	198
rect	198	198	199	199
rect	198	199	199	200
rect	198	200	199	201
rect	198	201	199	202
rect	198	202	199	203
rect	198	203	199	204
rect	198	204	199	205
rect	198	205	199	206
rect	198	206	199	207
rect	198	207	199	208
rect	198	208	199	209
rect	198	209	199	210
rect	198	210	199	211
rect	198	211	199	212
rect	198	212	199	213
rect	198	213	199	214
rect	198	214	199	215
rect	198	215	199	216
rect	198	216	199	217
rect	198	217	199	218
rect	198	218	199	219
rect	198	219	199	220
rect	198	220	199	221
rect	198	221	199	222
rect	198	222	199	223
rect	198	223	199	224
rect	198	224	199	225
rect	198	225	199	226
rect	198	226	199	227
rect	198	227	199	228
rect	198	228	199	229
rect	198	229	199	230
rect	198	230	199	231
rect	198	231	199	232
rect	198	232	199	233
rect	198	233	199	234
rect	198	234	199	235
rect	198	235	199	236
rect	198	236	199	237
rect	198	237	199	238
rect	198	238	199	239
rect	198	239	199	240
rect	198	240	199	241
rect	198	241	199	242
rect	198	242	199	243
rect	198	243	199	244
rect	198	244	199	245
rect	198	245	199	246
rect	198	246	199	247
rect	198	247	199	248
rect	198	248	199	249
rect	198	249	199	250
rect	198	250	199	251
rect	198	251	199	252
rect	198	252	199	253
rect	198	253	199	254
rect	198	254	199	255
rect	198	255	199	256
rect	198	256	199	257
rect	198	257	199	258
rect	198	258	199	259
rect	198	259	199	260
rect	198	260	199	261
rect	198	261	199	262
rect	198	262	199	263
rect	198	263	199	264
rect	198	264	199	265
rect	198	265	199	266
rect	198	266	199	267
rect	198	267	199	268
rect	198	268	199	269
rect	198	269	199	270
rect	198	270	199	271
rect	198	271	199	272
rect	198	272	199	273
rect	198	273	199	274
rect	198	274	199	275
rect	198	275	199	276
rect	198	276	199	277
rect	198	277	199	278
rect	198	278	199	279
rect	198	279	199	280
rect	198	280	199	281
rect	198	281	199	282
rect	198	282	199	283
rect	198	283	199	284
rect	198	284	199	285
rect	198	285	199	286
rect	198	286	199	287
rect	198	287	199	288
rect	198	288	199	289
rect	198	289	199	290
rect	198	290	199	291
rect	198	291	199	292
rect	198	292	199	293
rect	198	293	199	294
rect	198	294	199	295
rect	198	295	199	296
rect	198	296	199	297
rect	198	297	199	298
rect	198	298	199	299
rect	198	299	199	300
rect	198	300	199	301
rect	198	301	199	302
rect	198	302	199	303
rect	198	303	199	304
rect	198	304	199	305
rect	198	305	199	306
rect	198	306	199	307
rect	198	307	199	308
rect	198	308	199	309
rect	198	309	199	310
rect	198	310	199	311
rect	198	311	199	312
rect	198	312	199	313
rect	198	313	199	314
rect	198	314	199	315
rect	198	315	199	316
rect	198	316	199	317
rect	198	317	199	318
rect	198	318	199	319
rect	198	319	199	320
rect	198	320	199	321
rect	198	321	199	322
rect	198	322	199	323
rect	198	323	199	324
rect	198	324	199	325
rect	198	325	199	326
rect	198	326	199	327
rect	198	327	199	328
rect	198	328	199	329
rect	198	329	199	330
rect	198	330	199	331
rect	198	331	199	332
rect	198	332	199	333
rect	198	333	199	334
rect	198	334	199	335
rect	198	335	199	336
rect	199	0	200	1
rect	199	1	200	2
rect	199	2	200	3
rect	199	3	200	4
rect	199	4	200	5
rect	199	5	200	6
rect	199	6	200	7
rect	199	7	200	8
rect	199	8	200	9
rect	199	9	200	10
rect	199	10	200	11
rect	199	11	200	12
rect	199	12	200	13
rect	199	13	200	14
rect	199	14	200	15
rect	199	15	200	16
rect	199	16	200	17
rect	199	17	200	18
rect	199	18	200	19
rect	199	19	200	20
rect	199	20	200	21
rect	199	21	200	22
rect	199	22	200	23
rect	199	23	200	24
rect	199	24	200	25
rect	199	25	200	26
rect	199	26	200	27
rect	199	27	200	28
rect	199	28	200	29
rect	199	29	200	30
rect	199	30	200	31
rect	199	31	200	32
rect	199	32	200	33
rect	199	33	200	34
rect	199	34	200	35
rect	199	35	200	36
rect	199	36	200	37
rect	199	37	200	38
rect	199	38	200	39
rect	199	39	200	40
rect	199	40	200	41
rect	199	41	200	42
rect	199	42	200	43
rect	199	43	200	44
rect	199	44	200	45
rect	199	45	200	46
rect	199	46	200	47
rect	199	47	200	48
rect	199	48	200	49
rect	199	49	200	50
rect	199	50	200	51
rect	199	51	200	52
rect	199	52	200	53
rect	199	53	200	54
rect	199	54	200	55
rect	199	55	200	56
rect	199	56	200	57
rect	199	57	200	58
rect	199	58	200	59
rect	199	59	200	60
rect	199	60	200	61
rect	199	61	200	62
rect	199	62	200	63
rect	199	63	200	64
rect	199	64	200	65
rect	199	65	200	66
rect	199	66	200	67
rect	199	67	200	68
rect	199	68	200	69
rect	199	69	200	70
rect	199	70	200	71
rect	199	71	200	72
rect	199	72	200	73
rect	199	73	200	74
rect	199	74	200	75
rect	199	75	200	76
rect	199	76	200	77
rect	199	77	200	78
rect	199	78	200	79
rect	199	79	200	80
rect	199	80	200	81
rect	199	81	200	82
rect	199	82	200	83
rect	199	83	200	84
rect	199	84	200	85
rect	199	85	200	86
rect	199	86	200	87
rect	199	87	200	88
rect	199	88	200	89
rect	199	89	200	90
rect	199	90	200	91
rect	199	91	200	92
rect	199	92	200	93
rect	199	93	200	94
rect	199	94	200	95
rect	199	95	200	96
rect	199	96	200	97
rect	199	97	200	98
rect	199	98	200	99
rect	199	99	200	100
rect	199	100	200	101
rect	199	101	200	102
rect	199	102	200	103
rect	199	103	200	104
rect	199	104	200	105
rect	199	105	200	106
rect	199	106	200	107
rect	199	107	200	108
rect	199	108	200	109
rect	199	109	200	110
rect	199	110	200	111
rect	199	111	200	112
rect	199	112	200	113
rect	199	113	200	114
rect	199	114	200	115
rect	199	115	200	116
rect	199	116	200	117
rect	199	117	200	118
rect	199	118	200	119
rect	199	119	200	120
rect	199	120	200	121
rect	199	121	200	122
rect	199	122	200	123
rect	199	123	200	124
rect	199	124	200	125
rect	199	125	200	126
rect	199	126	200	127
rect	199	127	200	128
rect	199	128	200	129
rect	199	129	200	130
rect	199	130	200	131
rect	199	131	200	132
rect	199	132	200	133
rect	199	133	200	134
rect	199	134	200	135
rect	199	135	200	136
rect	199	136	200	137
rect	199	137	200	138
rect	199	138	200	139
rect	199	139	200	140
rect	199	140	200	141
rect	199	141	200	142
rect	199	142	200	143
rect	199	143	200	144
rect	199	144	200	145
rect	199	145	200	146
rect	199	146	200	147
rect	199	147	200	148
rect	199	148	200	149
rect	199	149	200	150
rect	199	150	200	151
rect	199	151	200	152
rect	199	152	200	153
rect	199	153	200	154
rect	199	154	200	155
rect	199	155	200	156
rect	199	156	200	157
rect	199	157	200	158
rect	199	158	200	159
rect	199	159	200	160
rect	199	160	200	161
rect	199	161	200	162
rect	199	162	200	163
rect	199	163	200	164
rect	199	164	200	165
rect	199	165	200	166
rect	199	166	200	167
rect	199	167	200	168
rect	199	168	200	169
rect	199	169	200	170
rect	199	170	200	171
rect	199	171	200	172
rect	199	172	200	173
rect	199	173	200	174
rect	199	174	200	175
rect	199	175	200	176
rect	199	176	200	177
rect	199	177	200	178
rect	199	178	200	179
rect	199	179	200	180
rect	199	180	200	181
rect	199	181	200	182
rect	199	182	200	183
rect	199	183	200	184
rect	199	184	200	185
rect	199	185	200	186
rect	199	186	200	187
rect	199	187	200	188
rect	199	188	200	189
rect	199	189	200	190
rect	199	190	200	191
rect	199	191	200	192
rect	199	192	200	193
rect	199	193	200	194
rect	199	194	200	195
rect	199	195	200	196
rect	199	196	200	197
rect	199	197	200	198
rect	199	198	200	199
rect	199	199	200	200
rect	199	200	200	201
rect	199	201	200	202
rect	199	202	200	203
rect	199	203	200	204
rect	199	204	200	205
rect	199	205	200	206
rect	199	206	200	207
rect	199	207	200	208
rect	199	208	200	209
rect	199	209	200	210
rect	199	210	200	211
rect	199	211	200	212
rect	199	212	200	213
rect	199	213	200	214
rect	199	214	200	215
rect	199	215	200	216
rect	199	216	200	217
rect	199	217	200	218
rect	199	218	200	219
rect	199	219	200	220
rect	199	220	200	221
rect	199	221	200	222
rect	199	222	200	223
rect	199	223	200	224
rect	199	224	200	225
rect	199	225	200	226
rect	199	226	200	227
rect	199	227	200	228
rect	199	228	200	229
rect	199	229	200	230
rect	199	230	200	231
rect	199	231	200	232
rect	199	232	200	233
rect	199	233	200	234
rect	199	234	200	235
rect	199	235	200	236
rect	199	236	200	237
rect	199	237	200	238
rect	199	238	200	239
rect	199	239	200	240
rect	199	240	200	241
rect	199	241	200	242
rect	199	242	200	243
rect	199	243	200	244
rect	199	244	200	245
rect	199	245	200	246
rect	199	246	200	247
rect	199	247	200	248
rect	199	248	200	249
rect	199	249	200	250
rect	199	250	200	251
rect	199	251	200	252
rect	199	252	200	253
rect	199	253	200	254
rect	199	254	200	255
rect	199	255	200	256
rect	199	256	200	257
rect	199	257	200	258
rect	199	258	200	259
rect	199	259	200	260
rect	199	260	200	261
rect	199	261	200	262
rect	199	262	200	263
rect	199	263	200	264
rect	199	264	200	265
rect	199	265	200	266
rect	199	266	200	267
rect	199	267	200	268
rect	199	268	200	269
rect	199	269	200	270
rect	199	270	200	271
rect	199	271	200	272
rect	199	272	200	273
rect	199	273	200	274
rect	199	274	200	275
rect	199	275	200	276
rect	199	276	200	277
rect	199	277	200	278
rect	199	278	200	279
rect	199	279	200	280
rect	199	280	200	281
rect	199	281	200	282
rect	199	282	200	283
rect	199	283	200	284
rect	199	284	200	285
rect	199	285	200	286
rect	199	286	200	287
rect	199	287	200	288
rect	199	288	200	289
rect	199	289	200	290
rect	199	290	200	291
rect	199	291	200	292
rect	199	292	200	293
rect	199	293	200	294
rect	199	294	200	295
rect	199	295	200	296
rect	199	296	200	297
rect	199	297	200	298
rect	199	298	200	299
rect	199	299	200	300
rect	199	300	200	301
rect	199	301	200	302
rect	199	302	200	303
rect	199	303	200	304
rect	199	304	200	305
rect	199	305	200	306
rect	199	306	200	307
rect	199	307	200	308
rect	199	308	200	309
rect	199	309	200	310
rect	199	310	200	311
rect	199	311	200	312
rect	199	312	200	313
rect	199	313	200	314
rect	199	314	200	315
rect	199	315	200	316
rect	199	316	200	317
rect	199	317	200	318
rect	199	318	200	319
rect	199	319	200	320
rect	199	320	200	321
rect	199	321	200	322
rect	199	322	200	323
rect	199	323	200	324
rect	199	324	200	325
rect	199	325	200	326
rect	199	326	200	327
rect	199	327	200	328
rect	199	328	200	329
rect	199	329	200	330
rect	199	330	200	331
rect	199	331	200	332
rect	199	332	200	333
rect	199	333	200	334
rect	199	334	200	335
rect	199	335	200	336
rect	200	0	201	1
rect	200	1	201	2
rect	200	2	201	3
rect	200	3	201	4
rect	200	4	201	5
rect	200	5	201	6
rect	200	6	201	7
rect	200	7	201	8
rect	200	8	201	9
rect	200	9	201	10
rect	200	10	201	11
rect	200	11	201	12
rect	200	12	201	13
rect	200	13	201	14
rect	200	14	201	15
rect	200	15	201	16
rect	200	16	201	17
rect	200	17	201	18
rect	200	18	201	19
rect	200	19	201	20
rect	200	20	201	21
rect	200	21	201	22
rect	200	22	201	23
rect	200	23	201	24
rect	200	24	201	25
rect	200	25	201	26
rect	200	26	201	27
rect	200	27	201	28
rect	200	28	201	29
rect	200	29	201	30
rect	200	30	201	31
rect	200	31	201	32
rect	200	32	201	33
rect	200	33	201	34
rect	200	34	201	35
rect	200	35	201	36
rect	200	36	201	37
rect	200	37	201	38
rect	200	38	201	39
rect	200	39	201	40
rect	200	40	201	41
rect	200	41	201	42
rect	200	42	201	43
rect	200	43	201	44
rect	200	44	201	45
rect	200	45	201	46
rect	200	46	201	47
rect	200	47	201	48
rect	200	48	201	49
rect	200	49	201	50
rect	200	50	201	51
rect	200	51	201	52
rect	200	52	201	53
rect	200	53	201	54
rect	200	54	201	55
rect	200	55	201	56
rect	200	56	201	57
rect	200	57	201	58
rect	200	58	201	59
rect	200	59	201	60
rect	200	60	201	61
rect	200	61	201	62
rect	200	62	201	63
rect	200	63	201	64
rect	200	64	201	65
rect	200	65	201	66
rect	200	66	201	67
rect	200	67	201	68
rect	200	68	201	69
rect	200	69	201	70
rect	200	70	201	71
rect	200	71	201	72
rect	200	72	201	73
rect	200	73	201	74
rect	200	74	201	75
rect	200	75	201	76
rect	200	76	201	77
rect	200	77	201	78
rect	200	78	201	79
rect	200	79	201	80
rect	200	80	201	81
rect	200	81	201	82
rect	200	82	201	83
rect	200	83	201	84
rect	200	84	201	85
rect	200	85	201	86
rect	200	86	201	87
rect	200	87	201	88
rect	200	88	201	89
rect	200	89	201	90
rect	200	90	201	91
rect	200	91	201	92
rect	200	92	201	93
rect	200	93	201	94
rect	200	94	201	95
rect	200	95	201	96
rect	200	96	201	97
rect	200	97	201	98
rect	200	98	201	99
rect	200	99	201	100
rect	200	100	201	101
rect	200	101	201	102
rect	200	102	201	103
rect	200	103	201	104
rect	200	104	201	105
rect	200	105	201	106
rect	200	106	201	107
rect	200	107	201	108
rect	200	108	201	109
rect	200	109	201	110
rect	200	110	201	111
rect	200	111	201	112
rect	200	112	201	113
rect	200	113	201	114
rect	200	114	201	115
rect	200	115	201	116
rect	200	116	201	117
rect	200	117	201	118
rect	200	118	201	119
rect	200	119	201	120
rect	200	120	201	121
rect	200	121	201	122
rect	200	122	201	123
rect	200	123	201	124
rect	200	124	201	125
rect	200	125	201	126
rect	200	126	201	127
rect	200	127	201	128
rect	200	128	201	129
rect	200	129	201	130
rect	200	130	201	131
rect	200	131	201	132
rect	200	132	201	133
rect	200	133	201	134
rect	200	134	201	135
rect	200	135	201	136
rect	200	136	201	137
rect	200	137	201	138
rect	200	138	201	139
rect	200	139	201	140
rect	200	140	201	141
rect	200	141	201	142
rect	200	142	201	143
rect	200	143	201	144
rect	200	144	201	145
rect	200	145	201	146
rect	200	146	201	147
rect	200	147	201	148
rect	200	148	201	149
rect	200	149	201	150
rect	200	150	201	151
rect	200	151	201	152
rect	200	152	201	153
rect	200	153	201	154
rect	200	154	201	155
rect	200	155	201	156
rect	200	156	201	157
rect	200	157	201	158
rect	200	158	201	159
rect	200	159	201	160
rect	200	160	201	161
rect	200	161	201	162
rect	200	162	201	163
rect	200	163	201	164
rect	200	164	201	165
rect	200	165	201	166
rect	200	166	201	167
rect	200	167	201	168
rect	200	168	201	169
rect	200	169	201	170
rect	200	170	201	171
rect	200	171	201	172
rect	200	172	201	173
rect	200	173	201	174
rect	200	174	201	175
rect	200	175	201	176
rect	200	176	201	177
rect	200	177	201	178
rect	200	178	201	179
rect	200	179	201	180
rect	200	180	201	181
rect	200	181	201	182
rect	200	182	201	183
rect	200	183	201	184
rect	200	184	201	185
rect	200	185	201	186
rect	200	186	201	187
rect	200	187	201	188
rect	200	188	201	189
rect	200	189	201	190
rect	200	190	201	191
rect	200	191	201	192
rect	200	192	201	193
rect	200	193	201	194
rect	200	194	201	195
rect	200	195	201	196
rect	200	196	201	197
rect	200	197	201	198
rect	200	198	201	199
rect	200	199	201	200
rect	200	200	201	201
rect	200	201	201	202
rect	200	202	201	203
rect	200	203	201	204
rect	200	204	201	205
rect	200	205	201	206
rect	200	206	201	207
rect	200	207	201	208
rect	200	208	201	209
rect	200	209	201	210
rect	200	210	201	211
rect	200	211	201	212
rect	200	212	201	213
rect	200	213	201	214
rect	200	214	201	215
rect	200	215	201	216
rect	200	216	201	217
rect	200	217	201	218
rect	200	218	201	219
rect	200	219	201	220
rect	200	220	201	221
rect	200	221	201	222
rect	200	222	201	223
rect	200	223	201	224
rect	200	224	201	225
rect	200	225	201	226
rect	200	226	201	227
rect	200	227	201	228
rect	200	228	201	229
rect	200	229	201	230
rect	200	230	201	231
rect	200	231	201	232
rect	200	232	201	233
rect	200	233	201	234
rect	200	234	201	235
rect	200	235	201	236
rect	200	236	201	237
rect	200	237	201	238
rect	200	238	201	239
rect	200	239	201	240
rect	200	240	201	241
rect	200	241	201	242
rect	200	242	201	243
rect	200	243	201	244
rect	200	244	201	245
rect	200	245	201	246
rect	200	246	201	247
rect	200	247	201	248
rect	200	248	201	249
rect	200	249	201	250
rect	200	250	201	251
rect	200	251	201	252
rect	200	252	201	253
rect	200	253	201	254
rect	200	254	201	255
rect	200	255	201	256
rect	200	256	201	257
rect	200	257	201	258
rect	200	258	201	259
rect	200	259	201	260
rect	200	260	201	261
rect	200	261	201	262
rect	200	262	201	263
rect	200	263	201	264
rect	200	264	201	265
rect	200	265	201	266
rect	200	266	201	267
rect	200	267	201	268
rect	200	268	201	269
rect	200	269	201	270
rect	200	270	201	271
rect	200	271	201	272
rect	200	272	201	273
rect	200	273	201	274
rect	200	274	201	275
rect	200	275	201	276
rect	200	276	201	277
rect	200	277	201	278
rect	200	278	201	279
rect	200	279	201	280
rect	200	280	201	281
rect	200	281	201	282
rect	200	282	201	283
rect	200	283	201	284
rect	200	284	201	285
rect	200	285	201	286
rect	200	286	201	287
rect	200	287	201	288
rect	200	288	201	289
rect	200	289	201	290
rect	200	290	201	291
rect	200	291	201	292
rect	200	292	201	293
rect	200	293	201	294
rect	200	294	201	295
rect	200	295	201	296
rect	200	296	201	297
rect	200	297	201	298
rect	200	298	201	299
rect	200	299	201	300
rect	200	300	201	301
rect	200	301	201	302
rect	200	302	201	303
rect	200	303	201	304
rect	200	304	201	305
rect	200	305	201	306
rect	200	306	201	307
rect	200	307	201	308
rect	200	308	201	309
rect	200	309	201	310
rect	200	310	201	311
rect	200	311	201	312
rect	200	312	201	313
rect	200	313	201	314
rect	200	314	201	315
rect	200	315	201	316
rect	200	316	201	317
rect	200	317	201	318
rect	200	318	201	319
rect	200	319	201	320
rect	200	320	201	321
rect	200	321	201	322
rect	200	322	201	323
rect	200	323	201	324
rect	200	324	201	325
rect	200	325	201	326
rect	200	326	201	327
rect	200	327	201	328
rect	200	328	201	329
rect	200	329	201	330
rect	200	330	201	331
rect	200	331	201	332
rect	200	332	201	333
rect	200	333	201	334
rect	200	334	201	335
rect	200	335	201	336
rect	201	0	202	1
rect	201	1	202	2
rect	201	2	202	3
rect	201	3	202	4
rect	201	4	202	5
rect	201	5	202	6
rect	201	6	202	7
rect	201	7	202	8
rect	201	8	202	9
rect	201	9	202	10
rect	201	10	202	11
rect	201	11	202	12
rect	201	12	202	13
rect	201	13	202	14
rect	201	14	202	15
rect	201	15	202	16
rect	201	16	202	17
rect	201	17	202	18
rect	201	18	202	19
rect	201	19	202	20
rect	201	20	202	21
rect	201	21	202	22
rect	201	22	202	23
rect	201	23	202	24
rect	201	24	202	25
rect	201	25	202	26
rect	201	26	202	27
rect	201	27	202	28
rect	201	28	202	29
rect	201	29	202	30
rect	201	30	202	31
rect	201	31	202	32
rect	201	32	202	33
rect	201	33	202	34
rect	201	34	202	35
rect	201	35	202	36
rect	201	36	202	37
rect	201	37	202	38
rect	201	38	202	39
rect	201	39	202	40
rect	201	40	202	41
rect	201	41	202	42
rect	201	42	202	43
rect	201	43	202	44
rect	201	44	202	45
rect	201	45	202	46
rect	201	46	202	47
rect	201	47	202	48
rect	201	48	202	49
rect	201	49	202	50
rect	201	50	202	51
rect	201	51	202	52
rect	201	52	202	53
rect	201	53	202	54
rect	201	54	202	55
rect	201	55	202	56
rect	201	56	202	57
rect	201	57	202	58
rect	201	58	202	59
rect	201	59	202	60
rect	201	60	202	61
rect	201	61	202	62
rect	201	62	202	63
rect	201	63	202	64
rect	201	64	202	65
rect	201	65	202	66
rect	201	66	202	67
rect	201	67	202	68
rect	201	68	202	69
rect	201	69	202	70
rect	201	70	202	71
rect	201	71	202	72
rect	201	72	202	73
rect	201	73	202	74
rect	201	74	202	75
rect	201	75	202	76
rect	201	76	202	77
rect	201	77	202	78
rect	201	78	202	79
rect	201	79	202	80
rect	201	80	202	81
rect	201	81	202	82
rect	201	82	202	83
rect	201	83	202	84
rect	201	84	202	85
rect	201	85	202	86
rect	201	86	202	87
rect	201	87	202	88
rect	201	88	202	89
rect	201	89	202	90
rect	201	90	202	91
rect	201	91	202	92
rect	201	92	202	93
rect	201	93	202	94
rect	201	94	202	95
rect	201	95	202	96
rect	201	96	202	97
rect	201	97	202	98
rect	201	98	202	99
rect	201	99	202	100
rect	201	100	202	101
rect	201	101	202	102
rect	201	102	202	103
rect	201	103	202	104
rect	201	104	202	105
rect	201	105	202	106
rect	201	106	202	107
rect	201	107	202	108
rect	201	108	202	109
rect	201	109	202	110
rect	201	110	202	111
rect	201	111	202	112
rect	201	112	202	113
rect	201	113	202	114
rect	201	114	202	115
rect	201	115	202	116
rect	201	116	202	117
rect	201	117	202	118
rect	201	118	202	119
rect	201	119	202	120
rect	201	120	202	121
rect	201	121	202	122
rect	201	122	202	123
rect	201	123	202	124
rect	201	124	202	125
rect	201	125	202	126
rect	201	126	202	127
rect	201	127	202	128
rect	201	128	202	129
rect	201	129	202	130
rect	201	130	202	131
rect	201	131	202	132
rect	201	132	202	133
rect	201	133	202	134
rect	201	134	202	135
rect	201	135	202	136
rect	201	136	202	137
rect	201	137	202	138
rect	201	138	202	139
rect	201	139	202	140
rect	201	140	202	141
rect	201	141	202	142
rect	201	142	202	143
rect	201	143	202	144
rect	201	144	202	145
rect	201	145	202	146
rect	201	146	202	147
rect	201	147	202	148
rect	201	148	202	149
rect	201	149	202	150
rect	201	150	202	151
rect	201	151	202	152
rect	201	152	202	153
rect	201	153	202	154
rect	201	154	202	155
rect	201	155	202	156
rect	201	156	202	157
rect	201	157	202	158
rect	201	158	202	159
rect	201	159	202	160
rect	201	160	202	161
rect	201	161	202	162
rect	201	162	202	163
rect	201	163	202	164
rect	201	164	202	165
rect	201	165	202	166
rect	201	166	202	167
rect	201	167	202	168
rect	201	168	202	169
rect	201	169	202	170
rect	201	170	202	171
rect	201	171	202	172
rect	201	172	202	173
rect	201	173	202	174
rect	201	174	202	175
rect	201	175	202	176
rect	201	176	202	177
rect	201	177	202	178
rect	201	178	202	179
rect	201	179	202	180
rect	201	180	202	181
rect	201	181	202	182
rect	201	182	202	183
rect	201	183	202	184
rect	201	184	202	185
rect	201	185	202	186
rect	201	186	202	187
rect	201	187	202	188
rect	201	188	202	189
rect	201	189	202	190
rect	201	190	202	191
rect	201	191	202	192
rect	201	192	202	193
rect	201	193	202	194
rect	201	194	202	195
rect	201	195	202	196
rect	201	196	202	197
rect	201	197	202	198
rect	201	198	202	199
rect	201	199	202	200
rect	201	200	202	201
rect	201	201	202	202
rect	201	202	202	203
rect	201	203	202	204
rect	201	204	202	205
rect	201	205	202	206
rect	201	206	202	207
rect	201	207	202	208
rect	201	208	202	209
rect	201	209	202	210
rect	201	210	202	211
rect	201	211	202	212
rect	201	212	202	213
rect	201	213	202	214
rect	201	214	202	215
rect	201	215	202	216
rect	201	216	202	217
rect	201	217	202	218
rect	201	218	202	219
rect	201	219	202	220
rect	201	220	202	221
rect	201	221	202	222
rect	201	222	202	223
rect	201	223	202	224
rect	201	224	202	225
rect	201	225	202	226
rect	201	226	202	227
rect	201	227	202	228
rect	201	228	202	229
rect	201	229	202	230
rect	201	230	202	231
rect	201	231	202	232
rect	201	232	202	233
rect	201	233	202	234
rect	201	234	202	235
rect	201	235	202	236
rect	201	236	202	237
rect	201	237	202	238
rect	201	238	202	239
rect	201	239	202	240
rect	201	240	202	241
rect	201	241	202	242
rect	201	242	202	243
rect	201	243	202	244
rect	201	244	202	245
rect	201	245	202	246
rect	201	246	202	247
rect	201	247	202	248
rect	201	248	202	249
rect	201	249	202	250
rect	201	250	202	251
rect	201	251	202	252
rect	201	252	202	253
rect	201	253	202	254
rect	201	254	202	255
rect	201	255	202	256
rect	201	256	202	257
rect	201	257	202	258
rect	201	258	202	259
rect	201	259	202	260
rect	201	260	202	261
rect	201	261	202	262
rect	201	262	202	263
rect	201	263	202	264
rect	201	264	202	265
rect	201	265	202	266
rect	201	266	202	267
rect	201	267	202	268
rect	201	268	202	269
rect	201	269	202	270
rect	201	270	202	271
rect	201	271	202	272
rect	201	272	202	273
rect	201	273	202	274
rect	201	274	202	275
rect	201	275	202	276
rect	201	276	202	277
rect	201	277	202	278
rect	201	278	202	279
rect	201	279	202	280
rect	201	280	202	281
rect	201	281	202	282
rect	201	282	202	283
rect	201	283	202	284
rect	201	284	202	285
rect	201	285	202	286
rect	201	286	202	287
rect	201	287	202	288
rect	201	288	202	289
rect	201	289	202	290
rect	201	290	202	291
rect	201	291	202	292
rect	201	292	202	293
rect	201	293	202	294
rect	201	294	202	295
rect	201	295	202	296
rect	201	296	202	297
rect	201	297	202	298
rect	201	298	202	299
rect	201	299	202	300
rect	201	300	202	301
rect	201	301	202	302
rect	201	302	202	303
rect	201	303	202	304
rect	201	304	202	305
rect	201	305	202	306
rect	201	306	202	307
rect	201	307	202	308
rect	201	308	202	309
rect	201	309	202	310
rect	201	310	202	311
rect	201	311	202	312
rect	201	312	202	313
rect	201	313	202	314
rect	201	314	202	315
rect	201	315	202	316
rect	201	316	202	317
rect	201	317	202	318
rect	201	318	202	319
rect	201	319	202	320
rect	201	320	202	321
rect	201	321	202	322
rect	201	322	202	323
rect	201	323	202	324
rect	201	324	202	325
rect	201	325	202	326
rect	201	326	202	327
rect	201	327	202	328
rect	201	328	202	329
rect	201	329	202	330
rect	201	330	202	331
rect	201	331	202	332
rect	201	332	202	333
rect	201	333	202	334
rect	201	334	202	335
rect	201	335	202	336
rect	202	0	203	1
rect	202	1	203	2
rect	202	2	203	3
rect	202	3	203	4
rect	202	4	203	5
rect	202	5	203	6
rect	202	6	203	7
rect	202	7	203	8
rect	202	8	203	9
rect	202	9	203	10
rect	202	10	203	11
rect	202	11	203	12
rect	202	12	203	13
rect	202	13	203	14
rect	202	14	203	15
rect	202	15	203	16
rect	202	16	203	17
rect	202	17	203	18
rect	202	18	203	19
rect	202	19	203	20
rect	202	20	203	21
rect	202	21	203	22
rect	202	22	203	23
rect	202	23	203	24
rect	202	24	203	25
rect	202	25	203	26
rect	202	26	203	27
rect	202	27	203	28
rect	202	28	203	29
rect	202	29	203	30
rect	202	30	203	31
rect	202	31	203	32
rect	202	32	203	33
rect	202	33	203	34
rect	202	34	203	35
rect	202	35	203	36
rect	202	36	203	37
rect	202	37	203	38
rect	202	38	203	39
rect	202	39	203	40
rect	202	40	203	41
rect	202	41	203	42
rect	202	42	203	43
rect	202	43	203	44
rect	202	44	203	45
rect	202	45	203	46
rect	202	46	203	47
rect	202	47	203	48
rect	202	48	203	49
rect	202	49	203	50
rect	202	50	203	51
rect	202	51	203	52
rect	202	52	203	53
rect	202	53	203	54
rect	202	54	203	55
rect	202	55	203	56
rect	202	56	203	57
rect	202	57	203	58
rect	202	58	203	59
rect	202	59	203	60
rect	202	60	203	61
rect	202	61	203	62
rect	202	62	203	63
rect	202	63	203	64
rect	202	64	203	65
rect	202	65	203	66
rect	202	66	203	67
rect	202	67	203	68
rect	202	68	203	69
rect	202	69	203	70
rect	202	70	203	71
rect	202	71	203	72
rect	202	72	203	73
rect	202	73	203	74
rect	202	74	203	75
rect	202	75	203	76
rect	202	76	203	77
rect	202	77	203	78
rect	202	78	203	79
rect	202	79	203	80
rect	202	80	203	81
rect	202	81	203	82
rect	202	82	203	83
rect	202	83	203	84
rect	202	84	203	85
rect	202	85	203	86
rect	202	86	203	87
rect	202	87	203	88
rect	202	88	203	89
rect	202	89	203	90
rect	202	90	203	91
rect	202	91	203	92
rect	202	92	203	93
rect	202	93	203	94
rect	202	94	203	95
rect	202	95	203	96
rect	202	96	203	97
rect	202	97	203	98
rect	202	98	203	99
rect	202	99	203	100
rect	202	100	203	101
rect	202	101	203	102
rect	202	102	203	103
rect	202	103	203	104
rect	202	104	203	105
rect	202	105	203	106
rect	202	106	203	107
rect	202	107	203	108
rect	202	108	203	109
rect	202	109	203	110
rect	202	110	203	111
rect	202	111	203	112
rect	202	112	203	113
rect	202	113	203	114
rect	202	114	203	115
rect	202	115	203	116
rect	202	116	203	117
rect	202	117	203	118
rect	202	118	203	119
rect	202	119	203	120
rect	202	120	203	121
rect	202	121	203	122
rect	202	122	203	123
rect	202	123	203	124
rect	202	124	203	125
rect	202	125	203	126
rect	202	126	203	127
rect	202	127	203	128
rect	202	128	203	129
rect	202	129	203	130
rect	202	130	203	131
rect	202	131	203	132
rect	202	132	203	133
rect	202	133	203	134
rect	202	134	203	135
rect	202	135	203	136
rect	202	136	203	137
rect	202	137	203	138
rect	202	138	203	139
rect	202	139	203	140
rect	202	140	203	141
rect	202	141	203	142
rect	202	142	203	143
rect	202	143	203	144
rect	202	144	203	145
rect	202	145	203	146
rect	202	146	203	147
rect	202	147	203	148
rect	202	148	203	149
rect	202	149	203	150
rect	202	150	203	151
rect	202	151	203	152
rect	202	152	203	153
rect	202	153	203	154
rect	202	154	203	155
rect	202	155	203	156
rect	202	156	203	157
rect	202	157	203	158
rect	202	158	203	159
rect	202	159	203	160
rect	202	160	203	161
rect	202	161	203	162
rect	202	162	203	163
rect	202	163	203	164
rect	202	164	203	165
rect	202	165	203	166
rect	202	166	203	167
rect	202	167	203	168
rect	202	168	203	169
rect	202	169	203	170
rect	202	170	203	171
rect	202	171	203	172
rect	202	172	203	173
rect	202	173	203	174
rect	202	174	203	175
rect	202	175	203	176
rect	202	176	203	177
rect	202	177	203	178
rect	202	178	203	179
rect	202	179	203	180
rect	202	180	203	181
rect	202	181	203	182
rect	202	182	203	183
rect	202	183	203	184
rect	202	184	203	185
rect	202	185	203	186
rect	202	186	203	187
rect	202	187	203	188
rect	202	188	203	189
rect	202	189	203	190
rect	202	190	203	191
rect	202	191	203	192
rect	202	192	203	193
rect	202	193	203	194
rect	202	194	203	195
rect	202	195	203	196
rect	202	196	203	197
rect	202	197	203	198
rect	202	198	203	199
rect	202	199	203	200
rect	202	200	203	201
rect	202	201	203	202
rect	202	202	203	203
rect	202	203	203	204
rect	202	204	203	205
rect	202	205	203	206
rect	202	206	203	207
rect	202	207	203	208
rect	202	208	203	209
rect	202	209	203	210
rect	202	210	203	211
rect	202	211	203	212
rect	202	212	203	213
rect	202	213	203	214
rect	202	214	203	215
rect	202	215	203	216
rect	202	216	203	217
rect	202	217	203	218
rect	202	218	203	219
rect	202	219	203	220
rect	202	220	203	221
rect	202	221	203	222
rect	202	222	203	223
rect	202	223	203	224
rect	202	224	203	225
rect	202	225	203	226
rect	202	226	203	227
rect	202	227	203	228
rect	202	228	203	229
rect	202	229	203	230
rect	202	230	203	231
rect	202	231	203	232
rect	202	232	203	233
rect	202	233	203	234
rect	202	234	203	235
rect	202	235	203	236
rect	202	236	203	237
rect	202	237	203	238
rect	202	238	203	239
rect	202	239	203	240
rect	202	240	203	241
rect	202	241	203	242
rect	202	242	203	243
rect	202	243	203	244
rect	202	244	203	245
rect	202	245	203	246
rect	202	246	203	247
rect	202	247	203	248
rect	202	248	203	249
rect	202	249	203	250
rect	202	250	203	251
rect	202	251	203	252
rect	202	252	203	253
rect	202	253	203	254
rect	202	254	203	255
rect	202	255	203	256
rect	202	256	203	257
rect	202	257	203	258
rect	202	258	203	259
rect	202	259	203	260
rect	202	260	203	261
rect	202	261	203	262
rect	202	262	203	263
rect	202	263	203	264
rect	202	264	203	265
rect	202	265	203	266
rect	202	266	203	267
rect	202	267	203	268
rect	202	268	203	269
rect	202	269	203	270
rect	202	270	203	271
rect	202	271	203	272
rect	202	272	203	273
rect	202	273	203	274
rect	202	274	203	275
rect	202	275	203	276
rect	202	276	203	277
rect	202	277	203	278
rect	202	278	203	279
rect	202	279	203	280
rect	202	280	203	281
rect	202	281	203	282
rect	202	282	203	283
rect	202	283	203	284
rect	202	284	203	285
rect	202	285	203	286
rect	202	286	203	287
rect	202	287	203	288
rect	202	288	203	289
rect	202	289	203	290
rect	202	290	203	291
rect	202	291	203	292
rect	202	292	203	293
rect	202	293	203	294
rect	202	294	203	295
rect	202	295	203	296
rect	202	296	203	297
rect	202	297	203	298
rect	202	298	203	299
rect	202	299	203	300
rect	202	300	203	301
rect	202	301	203	302
rect	202	302	203	303
rect	202	303	203	304
rect	202	304	203	305
rect	202	305	203	306
rect	202	306	203	307
rect	202	307	203	308
rect	202	308	203	309
rect	202	309	203	310
rect	202	310	203	311
rect	202	311	203	312
rect	202	312	203	313
rect	202	313	203	314
rect	202	314	203	315
rect	202	315	203	316
rect	202	316	203	317
rect	202	317	203	318
rect	202	318	203	319
rect	202	319	203	320
rect	202	320	203	321
rect	202	321	203	322
rect	202	322	203	323
rect	202	323	203	324
rect	202	324	203	325
rect	202	325	203	326
rect	202	326	203	327
rect	202	327	203	328
rect	202	328	203	329
rect	202	329	203	330
rect	202	330	203	331
rect	202	331	203	332
rect	202	332	203	333
rect	202	333	203	334
rect	202	334	203	335
rect	202	335	203	336
rect	228	0	229	1
rect	228	1	229	2
rect	228	2	229	3
rect	228	3	229	4
rect	228	4	229	5
rect	228	5	229	6
rect	228	6	229	7
rect	228	7	229	8
rect	228	8	229	9
rect	228	9	229	10
rect	228	10	229	11
rect	228	11	229	12
rect	228	12	229	13
rect	228	13	229	14
rect	228	14	229	15
rect	228	15	229	16
rect	228	16	229	17
rect	228	17	229	18
rect	228	18	229	19
rect	228	19	229	20
rect	228	20	229	21
rect	228	21	229	22
rect	228	22	229	23
rect	228	23	229	24
rect	228	24	229	25
rect	228	25	229	26
rect	228	26	229	27
rect	228	27	229	28
rect	228	28	229	29
rect	228	29	229	30
rect	228	30	229	31
rect	228	31	229	32
rect	228	32	229	33
rect	228	33	229	34
rect	228	34	229	35
rect	228	35	229	36
rect	228	36	229	37
rect	228	37	229	38
rect	228	38	229	39
rect	228	39	229	40
rect	228	40	229	41
rect	228	41	229	42
rect	228	42	229	43
rect	228	43	229	44
rect	228	44	229	45
rect	228	45	229	46
rect	228	46	229	47
rect	228	47	229	48
rect	228	48	229	49
rect	228	49	229	50
rect	228	50	229	51
rect	228	51	229	52
rect	228	52	229	53
rect	228	53	229	54
rect	228	54	229	55
rect	228	55	229	56
rect	228	56	229	57
rect	228	57	229	58
rect	228	58	229	59
rect	228	59	229	60
rect	228	60	229	61
rect	228	61	229	62
rect	228	62	229	63
rect	228	63	229	64
rect	228	64	229	65
rect	228	65	229	66
rect	228	66	229	67
rect	228	67	229	68
rect	228	68	229	69
rect	228	69	229	70
rect	228	70	229	71
rect	228	71	229	72
rect	228	72	229	73
rect	228	73	229	74
rect	228	74	229	75
rect	228	75	229	76
rect	228	76	229	77
rect	228	77	229	78
rect	228	78	229	79
rect	228	79	229	80
rect	228	80	229	81
rect	228	81	229	82
rect	228	82	229	83
rect	228	83	229	84
rect	228	84	229	85
rect	228	85	229	86
rect	228	86	229	87
rect	228	87	229	88
rect	228	88	229	89
rect	228	89	229	90
rect	228	90	229	91
rect	228	91	229	92
rect	228	92	229	93
rect	228	93	229	94
rect	228	94	229	95
rect	228	95	229	96
rect	228	96	229	97
rect	228	97	229	98
rect	228	98	229	99
rect	228	99	229	100
rect	228	100	229	101
rect	228	101	229	102
rect	228	102	229	103
rect	228	103	229	104
rect	228	104	229	105
rect	228	105	229	106
rect	228	106	229	107
rect	228	107	229	108
rect	228	108	229	109
rect	228	109	229	110
rect	228	110	229	111
rect	228	111	229	112
rect	228	112	229	113
rect	228	113	229	114
rect	228	114	229	115
rect	228	115	229	116
rect	228	116	229	117
rect	228	117	229	118
rect	228	118	229	119
rect	228	119	229	120
rect	228	120	229	121
rect	228	121	229	122
rect	228	122	229	123
rect	228	123	229	124
rect	228	124	229	125
rect	228	125	229	126
rect	228	126	229	127
rect	228	127	229	128
rect	228	128	229	129
rect	228	129	229	130
rect	228	130	229	131
rect	228	131	229	132
rect	228	132	229	133
rect	228	133	229	134
rect	228	134	229	135
rect	228	135	229	136
rect	228	136	229	137
rect	228	137	229	138
rect	228	138	229	139
rect	228	139	229	140
rect	228	140	229	141
rect	228	141	229	142
rect	228	142	229	143
rect	228	143	229	144
rect	228	144	229	145
rect	228	145	229	146
rect	228	146	229	147
rect	228	147	229	148
rect	228	148	229	149
rect	228	149	229	150
rect	228	150	229	151
rect	228	151	229	152
rect	228	152	229	153
rect	228	153	229	154
rect	228	154	229	155
rect	228	155	229	156
rect	228	156	229	157
rect	228	157	229	158
rect	228	158	229	159
rect	228	159	229	160
rect	228	160	229	161
rect	228	161	229	162
rect	228	162	229	163
rect	228	163	229	164
rect	228	164	229	165
rect	228	165	229	166
rect	228	166	229	167
rect	228	167	229	168
rect	228	168	229	169
rect	228	169	229	170
rect	228	170	229	171
rect	228	171	229	172
rect	228	172	229	173
rect	228	173	229	174
rect	228	174	229	175
rect	228	175	229	176
rect	228	176	229	177
rect	228	177	229	178
rect	228	178	229	179
rect	228	179	229	180
rect	228	180	229	181
rect	228	181	229	182
rect	228	182	229	183
rect	228	183	229	184
rect	228	184	229	185
rect	228	185	229	186
rect	228	186	229	187
rect	228	187	229	188
rect	228	188	229	189
rect	228	189	229	190
rect	228	190	229	191
rect	228	191	229	192
rect	228	192	229	193
rect	228	193	229	194
rect	228	194	229	195
rect	228	195	229	196
rect	228	196	229	197
rect	228	197	229	198
rect	228	198	229	199
rect	228	199	229	200
rect	228	200	229	201
rect	228	201	229	202
rect	228	202	229	203
rect	228	203	229	204
rect	228	204	229	205
rect	228	205	229	206
rect	228	206	229	207
rect	228	207	229	208
rect	228	208	229	209
rect	228	209	229	210
rect	228	210	229	211
rect	228	211	229	212
rect	228	212	229	213
rect	228	213	229	214
rect	228	214	229	215
rect	228	215	229	216
rect	228	216	229	217
rect	228	217	229	218
rect	228	218	229	219
rect	228	219	229	220
rect	228	220	229	221
rect	228	221	229	222
rect	228	222	229	223
rect	228	223	229	224
rect	228	224	229	225
rect	228	225	229	226
rect	228	226	229	227
rect	228	227	229	228
rect	228	228	229	229
rect	228	229	229	230
rect	228	230	229	231
rect	228	231	229	232
rect	228	232	229	233
rect	228	233	229	234
rect	228	234	229	235
rect	228	235	229	236
rect	228	236	229	237
rect	228	237	229	238
rect	228	238	229	239
rect	228	239	229	240
rect	228	240	229	241
rect	228	241	229	242
rect	228	242	229	243
rect	228	243	229	244
rect	228	244	229	245
rect	228	245	229	246
rect	228	246	229	247
rect	228	247	229	248
rect	228	248	229	249
rect	228	249	229	250
rect	228	250	229	251
rect	228	251	229	252
rect	228	252	229	253
rect	228	253	229	254
rect	228	254	229	255
rect	228	255	229	256
rect	228	256	229	257
rect	228	257	229	258
rect	228	258	229	259
rect	228	259	229	260
rect	228	260	229	261
rect	228	261	229	262
rect	228	262	229	263
rect	228	263	229	264
rect	228	264	229	265
rect	228	265	229	266
rect	228	266	229	267
rect	228	267	229	268
rect	228	268	229	269
rect	228	269	229	270
rect	228	270	229	271
rect	228	271	229	272
rect	228	272	229	273
rect	228	273	229	274
rect	228	274	229	275
rect	228	275	229	276
rect	228	276	229	277
rect	228	277	229	278
rect	228	278	229	279
rect	228	279	229	280
rect	228	280	229	281
rect	228	281	229	282
rect	228	282	229	283
rect	228	283	229	284
rect	228	284	229	285
rect	228	285	229	286
rect	228	286	229	287
rect	228	287	229	288
rect	228	288	229	289
rect	228	289	229	290
rect	228	290	229	291
rect	228	291	229	292
rect	228	292	229	293
rect	228	293	229	294
rect	228	294	229	295
rect	228	295	229	296
rect	228	296	229	297
rect	228	297	229	298
rect	228	298	229	299
rect	228	299	229	300
rect	228	300	229	301
rect	228	301	229	302
rect	228	302	229	303
rect	228	303	229	304
rect	228	304	229	305
rect	228	305	229	306
rect	228	306	229	307
rect	228	307	229	308
rect	228	308	229	309
rect	228	309	229	310
rect	228	310	229	311
rect	228	311	229	312
rect	228	312	229	313
rect	228	313	229	314
rect	228	314	229	315
rect	228	315	229	316
rect	228	316	229	317
rect	228	317	229	318
rect	228	318	229	319
rect	228	319	229	320
rect	228	320	229	321
rect	228	321	229	322
rect	228	322	229	323
rect	228	323	229	324
rect	228	324	229	325
rect	228	325	229	326
rect	228	326	229	327
rect	228	327	229	328
rect	228	328	229	329
rect	228	329	229	330
rect	228	330	229	331
rect	228	331	229	332
rect	228	332	229	333
rect	228	333	229	334
rect	228	334	229	335
rect	228	335	229	336
rect	229	0	230	1
rect	229	1	230	2
rect	229	2	230	3
rect	229	3	230	4
rect	229	4	230	5
rect	229	5	230	6
rect	229	6	230	7
rect	229	7	230	8
rect	229	8	230	9
rect	229	9	230	10
rect	229	10	230	11
rect	229	11	230	12
rect	229	12	230	13
rect	229	13	230	14
rect	229	14	230	15
rect	229	15	230	16
rect	229	16	230	17
rect	229	17	230	18
rect	229	18	230	19
rect	229	19	230	20
rect	229	20	230	21
rect	229	21	230	22
rect	229	22	230	23
rect	229	23	230	24
rect	229	24	230	25
rect	229	25	230	26
rect	229	26	230	27
rect	229	27	230	28
rect	229	28	230	29
rect	229	29	230	30
rect	229	30	230	31
rect	229	31	230	32
rect	229	32	230	33
rect	229	33	230	34
rect	229	34	230	35
rect	229	35	230	36
rect	229	36	230	37
rect	229	37	230	38
rect	229	38	230	39
rect	229	39	230	40
rect	229	40	230	41
rect	229	41	230	42
rect	229	42	230	43
rect	229	43	230	44
rect	229	44	230	45
rect	229	45	230	46
rect	229	46	230	47
rect	229	47	230	48
rect	229	48	230	49
rect	229	49	230	50
rect	229	50	230	51
rect	229	51	230	52
rect	229	52	230	53
rect	229	53	230	54
rect	229	54	230	55
rect	229	55	230	56
rect	229	56	230	57
rect	229	57	230	58
rect	229	58	230	59
rect	229	59	230	60
rect	229	60	230	61
rect	229	61	230	62
rect	229	62	230	63
rect	229	63	230	64
rect	229	64	230	65
rect	229	65	230	66
rect	229	66	230	67
rect	229	67	230	68
rect	229	68	230	69
rect	229	69	230	70
rect	229	70	230	71
rect	229	71	230	72
rect	229	72	230	73
rect	229	73	230	74
rect	229	74	230	75
rect	229	75	230	76
rect	229	76	230	77
rect	229	77	230	78
rect	229	78	230	79
rect	229	79	230	80
rect	229	80	230	81
rect	229	81	230	82
rect	229	82	230	83
rect	229	83	230	84
rect	229	84	230	85
rect	229	85	230	86
rect	229	86	230	87
rect	229	87	230	88
rect	229	88	230	89
rect	229	89	230	90
rect	229	90	230	91
rect	229	91	230	92
rect	229	92	230	93
rect	229	93	230	94
rect	229	94	230	95
rect	229	95	230	96
rect	229	96	230	97
rect	229	97	230	98
rect	229	98	230	99
rect	229	99	230	100
rect	229	100	230	101
rect	229	101	230	102
rect	229	102	230	103
rect	229	103	230	104
rect	229	104	230	105
rect	229	105	230	106
rect	229	106	230	107
rect	229	107	230	108
rect	229	108	230	109
rect	229	109	230	110
rect	229	110	230	111
rect	229	111	230	112
rect	229	112	230	113
rect	229	113	230	114
rect	229	114	230	115
rect	229	115	230	116
rect	229	116	230	117
rect	229	117	230	118
rect	229	118	230	119
rect	229	119	230	120
rect	229	120	230	121
rect	229	121	230	122
rect	229	122	230	123
rect	229	123	230	124
rect	229	124	230	125
rect	229	125	230	126
rect	229	126	230	127
rect	229	127	230	128
rect	229	128	230	129
rect	229	129	230	130
rect	229	130	230	131
rect	229	131	230	132
rect	229	132	230	133
rect	229	133	230	134
rect	229	134	230	135
rect	229	135	230	136
rect	229	136	230	137
rect	229	137	230	138
rect	229	138	230	139
rect	229	139	230	140
rect	229	140	230	141
rect	229	141	230	142
rect	229	142	230	143
rect	229	143	230	144
rect	229	144	230	145
rect	229	145	230	146
rect	229	146	230	147
rect	229	147	230	148
rect	229	148	230	149
rect	229	149	230	150
rect	229	150	230	151
rect	229	151	230	152
rect	229	152	230	153
rect	229	153	230	154
rect	229	154	230	155
rect	229	155	230	156
rect	229	156	230	157
rect	229	157	230	158
rect	229	158	230	159
rect	229	159	230	160
rect	229	160	230	161
rect	229	161	230	162
rect	229	162	230	163
rect	229	163	230	164
rect	229	164	230	165
rect	229	165	230	166
rect	229	166	230	167
rect	229	167	230	168
rect	229	168	230	169
rect	229	169	230	170
rect	229	170	230	171
rect	229	171	230	172
rect	229	172	230	173
rect	229	173	230	174
rect	229	174	230	175
rect	229	175	230	176
rect	229	176	230	177
rect	229	177	230	178
rect	229	178	230	179
rect	229	179	230	180
rect	229	180	230	181
rect	229	181	230	182
rect	229	182	230	183
rect	229	183	230	184
rect	229	184	230	185
rect	229	185	230	186
rect	229	186	230	187
rect	229	187	230	188
rect	229	188	230	189
rect	229	189	230	190
rect	229	190	230	191
rect	229	191	230	192
rect	229	192	230	193
rect	229	193	230	194
rect	229	194	230	195
rect	229	195	230	196
rect	229	196	230	197
rect	229	197	230	198
rect	229	198	230	199
rect	229	199	230	200
rect	229	200	230	201
rect	229	201	230	202
rect	229	202	230	203
rect	229	203	230	204
rect	229	204	230	205
rect	229	205	230	206
rect	229	206	230	207
rect	229	207	230	208
rect	229	208	230	209
rect	229	209	230	210
rect	229	210	230	211
rect	229	211	230	212
rect	229	212	230	213
rect	229	213	230	214
rect	229	214	230	215
rect	229	215	230	216
rect	229	216	230	217
rect	229	217	230	218
rect	229	218	230	219
rect	229	219	230	220
rect	229	220	230	221
rect	229	221	230	222
rect	229	222	230	223
rect	229	223	230	224
rect	229	224	230	225
rect	229	225	230	226
rect	229	226	230	227
rect	229	227	230	228
rect	229	228	230	229
rect	229	229	230	230
rect	229	230	230	231
rect	229	231	230	232
rect	229	232	230	233
rect	229	233	230	234
rect	229	234	230	235
rect	229	235	230	236
rect	229	236	230	237
rect	229	237	230	238
rect	229	238	230	239
rect	229	239	230	240
rect	229	240	230	241
rect	229	241	230	242
rect	229	242	230	243
rect	229	243	230	244
rect	229	244	230	245
rect	229	245	230	246
rect	229	246	230	247
rect	229	247	230	248
rect	229	248	230	249
rect	229	249	230	250
rect	229	250	230	251
rect	229	251	230	252
rect	229	252	230	253
rect	229	253	230	254
rect	229	254	230	255
rect	229	255	230	256
rect	229	256	230	257
rect	229	257	230	258
rect	229	258	230	259
rect	229	259	230	260
rect	229	260	230	261
rect	229	261	230	262
rect	229	262	230	263
rect	229	263	230	264
rect	229	264	230	265
rect	229	265	230	266
rect	229	266	230	267
rect	229	267	230	268
rect	229	268	230	269
rect	229	269	230	270
rect	229	270	230	271
rect	229	271	230	272
rect	229	272	230	273
rect	229	273	230	274
rect	229	274	230	275
rect	229	275	230	276
rect	229	276	230	277
rect	229	277	230	278
rect	229	278	230	279
rect	229	279	230	280
rect	229	280	230	281
rect	229	281	230	282
rect	229	282	230	283
rect	229	283	230	284
rect	229	284	230	285
rect	229	285	230	286
rect	229	286	230	287
rect	229	287	230	288
rect	229	288	230	289
rect	229	289	230	290
rect	229	290	230	291
rect	229	291	230	292
rect	229	292	230	293
rect	229	293	230	294
rect	229	294	230	295
rect	229	295	230	296
rect	229	296	230	297
rect	229	297	230	298
rect	229	298	230	299
rect	229	299	230	300
rect	229	300	230	301
rect	229	301	230	302
rect	229	302	230	303
rect	229	303	230	304
rect	229	304	230	305
rect	229	305	230	306
rect	229	306	230	307
rect	229	307	230	308
rect	229	308	230	309
rect	229	309	230	310
rect	229	310	230	311
rect	229	311	230	312
rect	229	312	230	313
rect	229	313	230	314
rect	229	314	230	315
rect	229	315	230	316
rect	229	316	230	317
rect	229	317	230	318
rect	229	318	230	319
rect	229	319	230	320
rect	229	320	230	321
rect	229	321	230	322
rect	229	322	230	323
rect	229	323	230	324
rect	229	324	230	325
rect	229	325	230	326
rect	229	326	230	327
rect	229	327	230	328
rect	229	328	230	329
rect	229	329	230	330
rect	229	330	230	331
rect	229	331	230	332
rect	229	332	230	333
rect	229	333	230	334
rect	229	334	230	335
rect	229	335	230	336
rect	230	0	231	1
rect	230	1	231	2
rect	230	2	231	3
rect	230	3	231	4
rect	230	4	231	5
rect	230	5	231	6
rect	230	6	231	7
rect	230	7	231	8
rect	230	8	231	9
rect	230	9	231	10
rect	230	10	231	11
rect	230	11	231	12
rect	230	12	231	13
rect	230	13	231	14
rect	230	14	231	15
rect	230	15	231	16
rect	230	16	231	17
rect	230	17	231	18
rect	230	18	231	19
rect	230	19	231	20
rect	230	20	231	21
rect	230	21	231	22
rect	230	22	231	23
rect	230	23	231	24
rect	230	24	231	25
rect	230	25	231	26
rect	230	26	231	27
rect	230	27	231	28
rect	230	28	231	29
rect	230	29	231	30
rect	230	30	231	31
rect	230	31	231	32
rect	230	32	231	33
rect	230	33	231	34
rect	230	34	231	35
rect	230	35	231	36
rect	230	36	231	37
rect	230	37	231	38
rect	230	38	231	39
rect	230	39	231	40
rect	230	40	231	41
rect	230	41	231	42
rect	230	42	231	43
rect	230	43	231	44
rect	230	44	231	45
rect	230	45	231	46
rect	230	46	231	47
rect	230	47	231	48
rect	230	48	231	49
rect	230	49	231	50
rect	230	50	231	51
rect	230	51	231	52
rect	230	52	231	53
rect	230	53	231	54
rect	230	54	231	55
rect	230	55	231	56
rect	230	56	231	57
rect	230	57	231	58
rect	230	58	231	59
rect	230	59	231	60
rect	230	60	231	61
rect	230	61	231	62
rect	230	62	231	63
rect	230	63	231	64
rect	230	64	231	65
rect	230	65	231	66
rect	230	66	231	67
rect	230	67	231	68
rect	230	68	231	69
rect	230	69	231	70
rect	230	70	231	71
rect	230	71	231	72
rect	230	72	231	73
rect	230	73	231	74
rect	230	74	231	75
rect	230	75	231	76
rect	230	76	231	77
rect	230	77	231	78
rect	230	78	231	79
rect	230	79	231	80
rect	230	80	231	81
rect	230	81	231	82
rect	230	82	231	83
rect	230	83	231	84
rect	230	84	231	85
rect	230	85	231	86
rect	230	86	231	87
rect	230	87	231	88
rect	230	88	231	89
rect	230	89	231	90
rect	230	90	231	91
rect	230	91	231	92
rect	230	92	231	93
rect	230	93	231	94
rect	230	94	231	95
rect	230	95	231	96
rect	230	96	231	97
rect	230	97	231	98
rect	230	98	231	99
rect	230	99	231	100
rect	230	100	231	101
rect	230	101	231	102
rect	230	102	231	103
rect	230	103	231	104
rect	230	104	231	105
rect	230	105	231	106
rect	230	106	231	107
rect	230	107	231	108
rect	230	108	231	109
rect	230	109	231	110
rect	230	110	231	111
rect	230	111	231	112
rect	230	112	231	113
rect	230	113	231	114
rect	230	114	231	115
rect	230	115	231	116
rect	230	116	231	117
rect	230	117	231	118
rect	230	118	231	119
rect	230	119	231	120
rect	230	120	231	121
rect	230	121	231	122
rect	230	122	231	123
rect	230	123	231	124
rect	230	124	231	125
rect	230	125	231	126
rect	230	126	231	127
rect	230	127	231	128
rect	230	128	231	129
rect	230	129	231	130
rect	230	130	231	131
rect	230	131	231	132
rect	230	132	231	133
rect	230	133	231	134
rect	230	134	231	135
rect	230	135	231	136
rect	230	136	231	137
rect	230	137	231	138
rect	230	138	231	139
rect	230	139	231	140
rect	230	140	231	141
rect	230	141	231	142
rect	230	142	231	143
rect	230	143	231	144
rect	230	144	231	145
rect	230	145	231	146
rect	230	146	231	147
rect	230	147	231	148
rect	230	148	231	149
rect	230	149	231	150
rect	230	150	231	151
rect	230	151	231	152
rect	230	152	231	153
rect	230	153	231	154
rect	230	154	231	155
rect	230	155	231	156
rect	230	156	231	157
rect	230	157	231	158
rect	230	158	231	159
rect	230	159	231	160
rect	230	160	231	161
rect	230	161	231	162
rect	230	162	231	163
rect	230	163	231	164
rect	230	164	231	165
rect	230	165	231	166
rect	230	166	231	167
rect	230	167	231	168
rect	230	168	231	169
rect	230	169	231	170
rect	230	170	231	171
rect	230	171	231	172
rect	230	172	231	173
rect	230	173	231	174
rect	230	174	231	175
rect	230	175	231	176
rect	230	176	231	177
rect	230	177	231	178
rect	230	178	231	179
rect	230	179	231	180
rect	230	180	231	181
rect	230	181	231	182
rect	230	182	231	183
rect	230	183	231	184
rect	230	184	231	185
rect	230	185	231	186
rect	230	186	231	187
rect	230	187	231	188
rect	230	188	231	189
rect	230	189	231	190
rect	230	190	231	191
rect	230	191	231	192
rect	230	192	231	193
rect	230	193	231	194
rect	230	194	231	195
rect	230	195	231	196
rect	230	196	231	197
rect	230	197	231	198
rect	230	198	231	199
rect	230	199	231	200
rect	230	200	231	201
rect	230	201	231	202
rect	230	202	231	203
rect	230	203	231	204
rect	230	204	231	205
rect	230	205	231	206
rect	230	206	231	207
rect	230	207	231	208
rect	230	208	231	209
rect	230	209	231	210
rect	230	210	231	211
rect	230	211	231	212
rect	230	212	231	213
rect	230	213	231	214
rect	230	214	231	215
rect	230	215	231	216
rect	230	216	231	217
rect	230	217	231	218
rect	230	218	231	219
rect	230	219	231	220
rect	230	220	231	221
rect	230	221	231	222
rect	230	222	231	223
rect	230	223	231	224
rect	230	224	231	225
rect	230	225	231	226
rect	230	226	231	227
rect	230	227	231	228
rect	230	228	231	229
rect	230	229	231	230
rect	230	230	231	231
rect	230	231	231	232
rect	230	232	231	233
rect	230	233	231	234
rect	230	234	231	235
rect	230	235	231	236
rect	230	236	231	237
rect	230	237	231	238
rect	230	238	231	239
rect	230	239	231	240
rect	230	240	231	241
rect	230	241	231	242
rect	230	242	231	243
rect	230	243	231	244
rect	230	244	231	245
rect	230	245	231	246
rect	230	246	231	247
rect	230	247	231	248
rect	230	248	231	249
rect	230	249	231	250
rect	230	250	231	251
rect	230	251	231	252
rect	230	252	231	253
rect	230	253	231	254
rect	230	254	231	255
rect	230	255	231	256
rect	230	256	231	257
rect	230	257	231	258
rect	230	258	231	259
rect	230	259	231	260
rect	230	260	231	261
rect	230	261	231	262
rect	230	262	231	263
rect	230	263	231	264
rect	230	264	231	265
rect	230	265	231	266
rect	230	266	231	267
rect	230	267	231	268
rect	230	268	231	269
rect	230	269	231	270
rect	230	270	231	271
rect	230	271	231	272
rect	230	272	231	273
rect	230	273	231	274
rect	230	274	231	275
rect	230	275	231	276
rect	230	276	231	277
rect	230	277	231	278
rect	230	278	231	279
rect	230	279	231	280
rect	230	280	231	281
rect	230	281	231	282
rect	230	282	231	283
rect	230	283	231	284
rect	230	284	231	285
rect	230	285	231	286
rect	230	286	231	287
rect	230	287	231	288
rect	230	288	231	289
rect	230	289	231	290
rect	230	290	231	291
rect	230	291	231	292
rect	230	292	231	293
rect	230	293	231	294
rect	230	294	231	295
rect	230	295	231	296
rect	230	296	231	297
rect	230	297	231	298
rect	230	298	231	299
rect	230	299	231	300
rect	230	300	231	301
rect	230	301	231	302
rect	230	302	231	303
rect	230	303	231	304
rect	230	304	231	305
rect	230	305	231	306
rect	230	306	231	307
rect	230	307	231	308
rect	230	308	231	309
rect	230	309	231	310
rect	230	310	231	311
rect	230	311	231	312
rect	230	312	231	313
rect	230	313	231	314
rect	230	314	231	315
rect	230	315	231	316
rect	230	316	231	317
rect	230	317	231	318
rect	230	318	231	319
rect	230	319	231	320
rect	230	320	231	321
rect	230	321	231	322
rect	230	322	231	323
rect	230	323	231	324
rect	230	324	231	325
rect	230	325	231	326
rect	230	326	231	327
rect	230	327	231	328
rect	230	328	231	329
rect	230	329	231	330
rect	230	330	231	331
rect	230	331	231	332
rect	230	332	231	333
rect	230	333	231	334
rect	230	334	231	335
rect	230	335	231	336
rect	231	0	232	1
rect	231	1	232	2
rect	231	2	232	3
rect	231	3	232	4
rect	231	4	232	5
rect	231	5	232	6
rect	231	6	232	7
rect	231	7	232	8
rect	231	8	232	9
rect	231	9	232	10
rect	231	10	232	11
rect	231	11	232	12
rect	231	12	232	13
rect	231	13	232	14
rect	231	14	232	15
rect	231	15	232	16
rect	231	16	232	17
rect	231	17	232	18
rect	231	18	232	19
rect	231	19	232	20
rect	231	20	232	21
rect	231	21	232	22
rect	231	22	232	23
rect	231	23	232	24
rect	231	24	232	25
rect	231	25	232	26
rect	231	26	232	27
rect	231	27	232	28
rect	231	28	232	29
rect	231	29	232	30
rect	231	30	232	31
rect	231	31	232	32
rect	231	32	232	33
rect	231	33	232	34
rect	231	34	232	35
rect	231	35	232	36
rect	231	36	232	37
rect	231	37	232	38
rect	231	38	232	39
rect	231	39	232	40
rect	231	40	232	41
rect	231	41	232	42
rect	231	42	232	43
rect	231	43	232	44
rect	231	44	232	45
rect	231	45	232	46
rect	231	46	232	47
rect	231	47	232	48
rect	231	48	232	49
rect	231	49	232	50
rect	231	50	232	51
rect	231	51	232	52
rect	231	52	232	53
rect	231	53	232	54
rect	231	54	232	55
rect	231	55	232	56
rect	231	56	232	57
rect	231	57	232	58
rect	231	58	232	59
rect	231	59	232	60
rect	231	60	232	61
rect	231	61	232	62
rect	231	62	232	63
rect	231	63	232	64
rect	231	64	232	65
rect	231	65	232	66
rect	231	66	232	67
rect	231	67	232	68
rect	231	68	232	69
rect	231	69	232	70
rect	231	70	232	71
rect	231	71	232	72
rect	231	72	232	73
rect	231	73	232	74
rect	231	74	232	75
rect	231	75	232	76
rect	231	76	232	77
rect	231	77	232	78
rect	231	78	232	79
rect	231	79	232	80
rect	231	80	232	81
rect	231	81	232	82
rect	231	82	232	83
rect	231	83	232	84
rect	231	84	232	85
rect	231	85	232	86
rect	231	86	232	87
rect	231	87	232	88
rect	231	88	232	89
rect	231	89	232	90
rect	231	90	232	91
rect	231	91	232	92
rect	231	92	232	93
rect	231	93	232	94
rect	231	94	232	95
rect	231	95	232	96
rect	231	96	232	97
rect	231	97	232	98
rect	231	98	232	99
rect	231	99	232	100
rect	231	100	232	101
rect	231	101	232	102
rect	231	102	232	103
rect	231	103	232	104
rect	231	104	232	105
rect	231	105	232	106
rect	231	106	232	107
rect	231	107	232	108
rect	231	108	232	109
rect	231	109	232	110
rect	231	110	232	111
rect	231	111	232	112
rect	231	112	232	113
rect	231	113	232	114
rect	231	114	232	115
rect	231	115	232	116
rect	231	116	232	117
rect	231	117	232	118
rect	231	118	232	119
rect	231	119	232	120
rect	231	120	232	121
rect	231	121	232	122
rect	231	122	232	123
rect	231	123	232	124
rect	231	124	232	125
rect	231	125	232	126
rect	231	126	232	127
rect	231	127	232	128
rect	231	128	232	129
rect	231	129	232	130
rect	231	130	232	131
rect	231	131	232	132
rect	231	132	232	133
rect	231	133	232	134
rect	231	134	232	135
rect	231	135	232	136
rect	231	136	232	137
rect	231	137	232	138
rect	231	138	232	139
rect	231	139	232	140
rect	231	140	232	141
rect	231	141	232	142
rect	231	142	232	143
rect	231	143	232	144
rect	231	144	232	145
rect	231	145	232	146
rect	231	146	232	147
rect	231	147	232	148
rect	231	148	232	149
rect	231	149	232	150
rect	231	150	232	151
rect	231	151	232	152
rect	231	152	232	153
rect	231	153	232	154
rect	231	154	232	155
rect	231	155	232	156
rect	231	156	232	157
rect	231	157	232	158
rect	231	158	232	159
rect	231	159	232	160
rect	231	160	232	161
rect	231	161	232	162
rect	231	162	232	163
rect	231	163	232	164
rect	231	164	232	165
rect	231	165	232	166
rect	231	166	232	167
rect	231	167	232	168
rect	231	168	232	169
rect	231	169	232	170
rect	231	170	232	171
rect	231	171	232	172
rect	231	172	232	173
rect	231	173	232	174
rect	231	174	232	175
rect	231	175	232	176
rect	231	176	232	177
rect	231	177	232	178
rect	231	178	232	179
rect	231	179	232	180
rect	231	180	232	181
rect	231	181	232	182
rect	231	182	232	183
rect	231	183	232	184
rect	231	184	232	185
rect	231	185	232	186
rect	231	186	232	187
rect	231	187	232	188
rect	231	188	232	189
rect	231	189	232	190
rect	231	190	232	191
rect	231	191	232	192
rect	231	192	232	193
rect	231	193	232	194
rect	231	194	232	195
rect	231	195	232	196
rect	231	196	232	197
rect	231	197	232	198
rect	231	198	232	199
rect	231	199	232	200
rect	231	200	232	201
rect	231	201	232	202
rect	231	202	232	203
rect	231	203	232	204
rect	231	204	232	205
rect	231	205	232	206
rect	231	206	232	207
rect	231	207	232	208
rect	231	208	232	209
rect	231	209	232	210
rect	231	210	232	211
rect	231	211	232	212
rect	231	212	232	213
rect	231	213	232	214
rect	231	214	232	215
rect	231	215	232	216
rect	231	216	232	217
rect	231	217	232	218
rect	231	218	232	219
rect	231	219	232	220
rect	231	220	232	221
rect	231	221	232	222
rect	231	222	232	223
rect	231	223	232	224
rect	231	224	232	225
rect	231	225	232	226
rect	231	226	232	227
rect	231	227	232	228
rect	231	228	232	229
rect	231	229	232	230
rect	231	230	232	231
rect	231	231	232	232
rect	231	232	232	233
rect	231	233	232	234
rect	231	234	232	235
rect	231	235	232	236
rect	231	236	232	237
rect	231	237	232	238
rect	231	238	232	239
rect	231	239	232	240
rect	231	240	232	241
rect	231	241	232	242
rect	231	242	232	243
rect	231	243	232	244
rect	231	244	232	245
rect	231	245	232	246
rect	231	246	232	247
rect	231	247	232	248
rect	231	248	232	249
rect	231	249	232	250
rect	231	250	232	251
rect	231	251	232	252
rect	231	252	232	253
rect	231	253	232	254
rect	231	254	232	255
rect	231	255	232	256
rect	231	256	232	257
rect	231	257	232	258
rect	231	258	232	259
rect	231	259	232	260
rect	231	260	232	261
rect	231	261	232	262
rect	231	262	232	263
rect	231	263	232	264
rect	231	264	232	265
rect	231	265	232	266
rect	231	266	232	267
rect	231	267	232	268
rect	231	268	232	269
rect	231	269	232	270
rect	231	270	232	271
rect	231	271	232	272
rect	231	272	232	273
rect	231	273	232	274
rect	231	274	232	275
rect	231	275	232	276
rect	231	276	232	277
rect	231	277	232	278
rect	231	278	232	279
rect	231	279	232	280
rect	231	280	232	281
rect	231	281	232	282
rect	231	282	232	283
rect	231	283	232	284
rect	231	284	232	285
rect	231	285	232	286
rect	231	286	232	287
rect	231	287	232	288
rect	231	288	232	289
rect	231	289	232	290
rect	231	290	232	291
rect	231	291	232	292
rect	231	292	232	293
rect	231	293	232	294
rect	231	294	232	295
rect	231	295	232	296
rect	231	296	232	297
rect	231	297	232	298
rect	231	298	232	299
rect	231	299	232	300
rect	231	300	232	301
rect	231	301	232	302
rect	231	302	232	303
rect	231	303	232	304
rect	231	304	232	305
rect	231	305	232	306
rect	231	306	232	307
rect	231	307	232	308
rect	231	308	232	309
rect	231	309	232	310
rect	231	310	232	311
rect	231	311	232	312
rect	231	312	232	313
rect	231	313	232	314
rect	231	314	232	315
rect	231	315	232	316
rect	231	316	232	317
rect	231	317	232	318
rect	231	318	232	319
rect	231	319	232	320
rect	231	320	232	321
rect	231	321	232	322
rect	231	322	232	323
rect	231	323	232	324
rect	231	324	232	325
rect	231	325	232	326
rect	231	326	232	327
rect	231	327	232	328
rect	231	328	232	329
rect	231	329	232	330
rect	231	330	232	331
rect	231	331	232	332
rect	231	332	232	333
rect	231	333	232	334
rect	231	334	232	335
rect	231	335	232	336
rect	232	0	233	1
rect	232	1	233	2
rect	232	2	233	3
rect	232	3	233	4
rect	232	4	233	5
rect	232	5	233	6
rect	232	6	233	7
rect	232	7	233	8
rect	232	8	233	9
rect	232	9	233	10
rect	232	10	233	11
rect	232	11	233	12
rect	232	12	233	13
rect	232	13	233	14
rect	232	14	233	15
rect	232	15	233	16
rect	232	16	233	17
rect	232	17	233	18
rect	232	18	233	19
rect	232	19	233	20
rect	232	20	233	21
rect	232	21	233	22
rect	232	22	233	23
rect	232	23	233	24
rect	232	24	233	25
rect	232	25	233	26
rect	232	26	233	27
rect	232	27	233	28
rect	232	28	233	29
rect	232	29	233	30
rect	232	30	233	31
rect	232	31	233	32
rect	232	32	233	33
rect	232	33	233	34
rect	232	34	233	35
rect	232	35	233	36
rect	232	36	233	37
rect	232	37	233	38
rect	232	38	233	39
rect	232	39	233	40
rect	232	40	233	41
rect	232	41	233	42
rect	232	42	233	43
rect	232	43	233	44
rect	232	44	233	45
rect	232	45	233	46
rect	232	46	233	47
rect	232	47	233	48
rect	232	48	233	49
rect	232	49	233	50
rect	232	50	233	51
rect	232	51	233	52
rect	232	52	233	53
rect	232	53	233	54
rect	232	54	233	55
rect	232	55	233	56
rect	232	56	233	57
rect	232	57	233	58
rect	232	58	233	59
rect	232	59	233	60
rect	232	60	233	61
rect	232	61	233	62
rect	232	62	233	63
rect	232	63	233	64
rect	232	64	233	65
rect	232	65	233	66
rect	232	66	233	67
rect	232	67	233	68
rect	232	68	233	69
rect	232	69	233	70
rect	232	70	233	71
rect	232	71	233	72
rect	232	72	233	73
rect	232	73	233	74
rect	232	74	233	75
rect	232	75	233	76
rect	232	76	233	77
rect	232	77	233	78
rect	232	78	233	79
rect	232	79	233	80
rect	232	80	233	81
rect	232	81	233	82
rect	232	82	233	83
rect	232	83	233	84
rect	232	84	233	85
rect	232	85	233	86
rect	232	86	233	87
rect	232	87	233	88
rect	232	88	233	89
rect	232	89	233	90
rect	232	90	233	91
rect	232	91	233	92
rect	232	92	233	93
rect	232	93	233	94
rect	232	94	233	95
rect	232	95	233	96
rect	232	96	233	97
rect	232	97	233	98
rect	232	98	233	99
rect	232	99	233	100
rect	232	100	233	101
rect	232	101	233	102
rect	232	102	233	103
rect	232	103	233	104
rect	232	104	233	105
rect	232	105	233	106
rect	232	106	233	107
rect	232	107	233	108
rect	232	108	233	109
rect	232	109	233	110
rect	232	110	233	111
rect	232	111	233	112
rect	232	112	233	113
rect	232	113	233	114
rect	232	114	233	115
rect	232	115	233	116
rect	232	116	233	117
rect	232	117	233	118
rect	232	118	233	119
rect	232	119	233	120
rect	232	120	233	121
rect	232	121	233	122
rect	232	122	233	123
rect	232	123	233	124
rect	232	124	233	125
rect	232	125	233	126
rect	232	126	233	127
rect	232	127	233	128
rect	232	128	233	129
rect	232	129	233	130
rect	232	130	233	131
rect	232	131	233	132
rect	232	132	233	133
rect	232	133	233	134
rect	232	134	233	135
rect	232	135	233	136
rect	232	136	233	137
rect	232	137	233	138
rect	232	138	233	139
rect	232	139	233	140
rect	232	140	233	141
rect	232	141	233	142
rect	232	142	233	143
rect	232	143	233	144
rect	232	144	233	145
rect	232	145	233	146
rect	232	146	233	147
rect	232	147	233	148
rect	232	148	233	149
rect	232	149	233	150
rect	232	150	233	151
rect	232	151	233	152
rect	232	152	233	153
rect	232	153	233	154
rect	232	154	233	155
rect	232	155	233	156
rect	232	156	233	157
rect	232	157	233	158
rect	232	158	233	159
rect	232	159	233	160
rect	232	160	233	161
rect	232	161	233	162
rect	232	162	233	163
rect	232	163	233	164
rect	232	164	233	165
rect	232	165	233	166
rect	232	166	233	167
rect	232	167	233	168
rect	232	168	233	169
rect	232	169	233	170
rect	232	170	233	171
rect	232	171	233	172
rect	232	172	233	173
rect	232	173	233	174
rect	232	174	233	175
rect	232	175	233	176
rect	232	176	233	177
rect	232	177	233	178
rect	232	178	233	179
rect	232	179	233	180
rect	232	180	233	181
rect	232	181	233	182
rect	232	182	233	183
rect	232	183	233	184
rect	232	184	233	185
rect	232	185	233	186
rect	232	186	233	187
rect	232	187	233	188
rect	232	188	233	189
rect	232	189	233	190
rect	232	190	233	191
rect	232	191	233	192
rect	232	192	233	193
rect	232	193	233	194
rect	232	194	233	195
rect	232	195	233	196
rect	232	196	233	197
rect	232	197	233	198
rect	232	198	233	199
rect	232	199	233	200
rect	232	200	233	201
rect	232	201	233	202
rect	232	202	233	203
rect	232	203	233	204
rect	232	204	233	205
rect	232	205	233	206
rect	232	206	233	207
rect	232	207	233	208
rect	232	208	233	209
rect	232	209	233	210
rect	232	210	233	211
rect	232	211	233	212
rect	232	212	233	213
rect	232	213	233	214
rect	232	214	233	215
rect	232	215	233	216
rect	232	216	233	217
rect	232	217	233	218
rect	232	218	233	219
rect	232	219	233	220
rect	232	220	233	221
rect	232	221	233	222
rect	232	222	233	223
rect	232	223	233	224
rect	232	224	233	225
rect	232	225	233	226
rect	232	226	233	227
rect	232	227	233	228
rect	232	228	233	229
rect	232	229	233	230
rect	232	230	233	231
rect	232	231	233	232
rect	232	232	233	233
rect	232	233	233	234
rect	232	234	233	235
rect	232	235	233	236
rect	232	236	233	237
rect	232	237	233	238
rect	232	238	233	239
rect	232	239	233	240
rect	232	240	233	241
rect	232	241	233	242
rect	232	242	233	243
rect	232	243	233	244
rect	232	244	233	245
rect	232	245	233	246
rect	232	246	233	247
rect	232	247	233	248
rect	232	248	233	249
rect	232	249	233	250
rect	232	250	233	251
rect	232	251	233	252
rect	232	252	233	253
rect	232	253	233	254
rect	232	254	233	255
rect	232	255	233	256
rect	232	256	233	257
rect	232	257	233	258
rect	232	258	233	259
rect	232	259	233	260
rect	232	260	233	261
rect	232	261	233	262
rect	232	262	233	263
rect	232	263	233	264
rect	232	264	233	265
rect	232	265	233	266
rect	232	266	233	267
rect	232	267	233	268
rect	232	268	233	269
rect	232	269	233	270
rect	232	270	233	271
rect	232	271	233	272
rect	232	272	233	273
rect	232	273	233	274
rect	232	274	233	275
rect	232	275	233	276
rect	232	276	233	277
rect	232	277	233	278
rect	232	278	233	279
rect	232	279	233	280
rect	232	280	233	281
rect	232	281	233	282
rect	232	282	233	283
rect	232	283	233	284
rect	232	284	233	285
rect	232	285	233	286
rect	232	286	233	287
rect	232	287	233	288
rect	232	288	233	289
rect	232	289	233	290
rect	232	290	233	291
rect	232	291	233	292
rect	232	292	233	293
rect	232	293	233	294
rect	232	294	233	295
rect	232	295	233	296
rect	232	296	233	297
rect	232	297	233	298
rect	232	298	233	299
rect	232	299	233	300
rect	232	300	233	301
rect	232	301	233	302
rect	232	302	233	303
rect	232	303	233	304
rect	232	304	233	305
rect	232	305	233	306
rect	232	306	233	307
rect	232	307	233	308
rect	232	308	233	309
rect	232	309	233	310
rect	232	310	233	311
rect	232	311	233	312
rect	232	312	233	313
rect	232	313	233	314
rect	232	314	233	315
rect	232	315	233	316
rect	232	316	233	317
rect	232	317	233	318
rect	232	318	233	319
rect	232	319	233	320
rect	232	320	233	321
rect	232	321	233	322
rect	232	322	233	323
rect	232	323	233	324
rect	232	324	233	325
rect	232	325	233	326
rect	232	326	233	327
rect	232	327	233	328
rect	232	328	233	329
rect	232	329	233	330
rect	232	330	233	331
rect	232	331	233	332
rect	232	332	233	333
rect	232	333	233	334
rect	232	334	233	335
rect	232	335	233	336
rect	233	0	234	1
rect	233	1	234	2
rect	233	2	234	3
rect	233	3	234	4
rect	233	4	234	5
rect	233	5	234	6
rect	233	6	234	7
rect	233	7	234	8
rect	233	8	234	9
rect	233	9	234	10
rect	233	10	234	11
rect	233	11	234	12
rect	233	12	234	13
rect	233	13	234	14
rect	233	14	234	15
rect	233	15	234	16
rect	233	16	234	17
rect	233	17	234	18
rect	233	18	234	19
rect	233	19	234	20
rect	233	20	234	21
rect	233	21	234	22
rect	233	22	234	23
rect	233	23	234	24
rect	233	24	234	25
rect	233	25	234	26
rect	233	26	234	27
rect	233	27	234	28
rect	233	28	234	29
rect	233	29	234	30
rect	233	30	234	31
rect	233	31	234	32
rect	233	32	234	33
rect	233	33	234	34
rect	233	34	234	35
rect	233	35	234	36
rect	233	36	234	37
rect	233	37	234	38
rect	233	38	234	39
rect	233	39	234	40
rect	233	40	234	41
rect	233	41	234	42
rect	233	42	234	43
rect	233	43	234	44
rect	233	44	234	45
rect	233	45	234	46
rect	233	46	234	47
rect	233	47	234	48
rect	233	48	234	49
rect	233	49	234	50
rect	233	50	234	51
rect	233	51	234	52
rect	233	52	234	53
rect	233	53	234	54
rect	233	54	234	55
rect	233	55	234	56
rect	233	56	234	57
rect	233	57	234	58
rect	233	58	234	59
rect	233	59	234	60
rect	233	60	234	61
rect	233	61	234	62
rect	233	62	234	63
rect	233	63	234	64
rect	233	64	234	65
rect	233	65	234	66
rect	233	66	234	67
rect	233	67	234	68
rect	233	68	234	69
rect	233	69	234	70
rect	233	70	234	71
rect	233	71	234	72
rect	233	72	234	73
rect	233	73	234	74
rect	233	74	234	75
rect	233	75	234	76
rect	233	76	234	77
rect	233	77	234	78
rect	233	78	234	79
rect	233	79	234	80
rect	233	80	234	81
rect	233	81	234	82
rect	233	82	234	83
rect	233	83	234	84
rect	233	84	234	85
rect	233	85	234	86
rect	233	86	234	87
rect	233	87	234	88
rect	233	88	234	89
rect	233	89	234	90
rect	233	90	234	91
rect	233	91	234	92
rect	233	92	234	93
rect	233	93	234	94
rect	233	94	234	95
rect	233	95	234	96
rect	233	96	234	97
rect	233	97	234	98
rect	233	98	234	99
rect	233	99	234	100
rect	233	100	234	101
rect	233	101	234	102
rect	233	102	234	103
rect	233	103	234	104
rect	233	104	234	105
rect	233	105	234	106
rect	233	106	234	107
rect	233	107	234	108
rect	233	108	234	109
rect	233	109	234	110
rect	233	110	234	111
rect	233	111	234	112
rect	233	112	234	113
rect	233	113	234	114
rect	233	114	234	115
rect	233	115	234	116
rect	233	116	234	117
rect	233	117	234	118
rect	233	118	234	119
rect	233	119	234	120
rect	233	120	234	121
rect	233	121	234	122
rect	233	122	234	123
rect	233	123	234	124
rect	233	124	234	125
rect	233	125	234	126
rect	233	126	234	127
rect	233	127	234	128
rect	233	128	234	129
rect	233	129	234	130
rect	233	130	234	131
rect	233	131	234	132
rect	233	132	234	133
rect	233	133	234	134
rect	233	134	234	135
rect	233	135	234	136
rect	233	136	234	137
rect	233	137	234	138
rect	233	138	234	139
rect	233	139	234	140
rect	233	140	234	141
rect	233	141	234	142
rect	233	142	234	143
rect	233	143	234	144
rect	233	144	234	145
rect	233	145	234	146
rect	233	146	234	147
rect	233	147	234	148
rect	233	148	234	149
rect	233	149	234	150
rect	233	150	234	151
rect	233	151	234	152
rect	233	152	234	153
rect	233	153	234	154
rect	233	154	234	155
rect	233	155	234	156
rect	233	156	234	157
rect	233	157	234	158
rect	233	158	234	159
rect	233	159	234	160
rect	233	160	234	161
rect	233	161	234	162
rect	233	162	234	163
rect	233	163	234	164
rect	233	164	234	165
rect	233	165	234	166
rect	233	166	234	167
rect	233	167	234	168
rect	233	168	234	169
rect	233	169	234	170
rect	233	170	234	171
rect	233	171	234	172
rect	233	172	234	173
rect	233	173	234	174
rect	233	174	234	175
rect	233	175	234	176
rect	233	176	234	177
rect	233	177	234	178
rect	233	178	234	179
rect	233	179	234	180
rect	233	180	234	181
rect	233	181	234	182
rect	233	182	234	183
rect	233	183	234	184
rect	233	184	234	185
rect	233	185	234	186
rect	233	186	234	187
rect	233	187	234	188
rect	233	188	234	189
rect	233	189	234	190
rect	233	190	234	191
rect	233	191	234	192
rect	233	192	234	193
rect	233	193	234	194
rect	233	194	234	195
rect	233	195	234	196
rect	233	196	234	197
rect	233	197	234	198
rect	233	198	234	199
rect	233	199	234	200
rect	233	200	234	201
rect	233	201	234	202
rect	233	202	234	203
rect	233	203	234	204
rect	233	204	234	205
rect	233	205	234	206
rect	233	206	234	207
rect	233	207	234	208
rect	233	208	234	209
rect	233	209	234	210
rect	233	210	234	211
rect	233	211	234	212
rect	233	212	234	213
rect	233	213	234	214
rect	233	214	234	215
rect	233	215	234	216
rect	233	216	234	217
rect	233	217	234	218
rect	233	218	234	219
rect	233	219	234	220
rect	233	220	234	221
rect	233	221	234	222
rect	233	222	234	223
rect	233	223	234	224
rect	233	224	234	225
rect	233	225	234	226
rect	233	226	234	227
rect	233	227	234	228
rect	233	228	234	229
rect	233	229	234	230
rect	233	230	234	231
rect	233	231	234	232
rect	233	232	234	233
rect	233	233	234	234
rect	233	234	234	235
rect	233	235	234	236
rect	233	236	234	237
rect	233	237	234	238
rect	233	238	234	239
rect	233	239	234	240
rect	233	240	234	241
rect	233	241	234	242
rect	233	242	234	243
rect	233	243	234	244
rect	233	244	234	245
rect	233	245	234	246
rect	233	246	234	247
rect	233	247	234	248
rect	233	248	234	249
rect	233	249	234	250
rect	233	250	234	251
rect	233	251	234	252
rect	233	252	234	253
rect	233	253	234	254
rect	233	254	234	255
rect	233	255	234	256
rect	233	256	234	257
rect	233	257	234	258
rect	233	258	234	259
rect	233	259	234	260
rect	233	260	234	261
rect	233	261	234	262
rect	233	262	234	263
rect	233	263	234	264
rect	233	264	234	265
rect	233	265	234	266
rect	233	266	234	267
rect	233	267	234	268
rect	233	268	234	269
rect	233	269	234	270
rect	233	270	234	271
rect	233	271	234	272
rect	233	272	234	273
rect	233	273	234	274
rect	233	274	234	275
rect	233	275	234	276
rect	233	276	234	277
rect	233	277	234	278
rect	233	278	234	279
rect	233	279	234	280
rect	233	280	234	281
rect	233	281	234	282
rect	233	282	234	283
rect	233	283	234	284
rect	233	284	234	285
rect	233	285	234	286
rect	233	286	234	287
rect	233	287	234	288
rect	233	288	234	289
rect	233	289	234	290
rect	233	290	234	291
rect	233	291	234	292
rect	233	292	234	293
rect	233	293	234	294
rect	233	294	234	295
rect	233	295	234	296
rect	233	296	234	297
rect	233	297	234	298
rect	233	298	234	299
rect	233	299	234	300
rect	233	300	234	301
rect	233	301	234	302
rect	233	302	234	303
rect	233	303	234	304
rect	233	304	234	305
rect	233	305	234	306
rect	233	306	234	307
rect	233	307	234	308
rect	233	308	234	309
rect	233	309	234	310
rect	233	310	234	311
rect	233	311	234	312
rect	233	312	234	313
rect	233	313	234	314
rect	233	314	234	315
rect	233	315	234	316
rect	233	316	234	317
rect	233	317	234	318
rect	233	318	234	319
rect	233	319	234	320
rect	233	320	234	321
rect	233	321	234	322
rect	233	322	234	323
rect	233	323	234	324
rect	233	324	234	325
rect	233	325	234	326
rect	233	326	234	327
rect	233	327	234	328
rect	233	328	234	329
rect	233	329	234	330
rect	233	330	234	331
rect	233	331	234	332
rect	233	332	234	333
rect	233	333	234	334
rect	233	334	234	335
rect	233	335	234	336
rect	245	323	246	324
rect	245	324	246	325
rect	245	325	246	326
rect	245	326	246	327
rect	245	327	246	328
rect	245	329	246	330
rect	245	330	246	331
rect	245	331	246	332
rect	245	332	246	333
rect	245	333	246	334
rect	245	334	246	335
rect	245	335	246	336
rect	245	336	246	337
rect	245	338	246	339
rect	245	339	246	340
rect	245	340	246	341
rect	245	341	246	342
rect	245	342	246	343
rect	245	343	246	344
rect	245	344	246	345
rect	245	345	246	346
rect	245	346	246	347
rect	245	347	246	348
rect	245	348	246	349
rect	245	349	246	350
rect	245	350	246	351
rect	245	351	246	352
rect	253	0	254	1
rect	253	1	254	2
rect	253	2	254	3
rect	253	3	254	4
rect	253	4	254	5
rect	253	5	254	6
rect	253	6	254	7
rect	253	7	254	8
rect	253	8	254	9
rect	253	9	254	10
rect	253	10	254	11
rect	253	11	254	12
rect	253	12	254	13
rect	253	13	254	14
rect	253	14	254	15
rect	253	15	254	16
rect	253	16	254	17
rect	253	17	254	18
rect	253	18	254	19
rect	253	19	254	20
rect	253	20	254	21
rect	253	21	254	22
rect	253	22	254	23
rect	253	23	254	24
rect	253	24	254	25
rect	253	25	254	26
rect	253	26	254	27
rect	253	27	254	28
rect	253	28	254	29
rect	253	29	254	30
rect	253	30	254	31
rect	253	31	254	32
rect	253	32	254	33
rect	253	33	254	34
rect	253	34	254	35
rect	253	35	254	36
rect	253	36	254	37
rect	253	37	254	38
rect	253	38	254	39
rect	253	39	254	40
rect	253	40	254	41
rect	253	41	254	42
rect	253	42	254	43
rect	253	43	254	44
rect	253	44	254	45
rect	253	45	254	46
rect	253	46	254	47
rect	253	47	254	48
rect	253	48	254	49
rect	253	49	254	50
rect	253	50	254	51
rect	253	51	254	52
rect	253	52	254	53
rect	253	53	254	54
rect	253	54	254	55
rect	253	55	254	56
rect	253	56	254	57
rect	253	57	254	58
rect	253	58	254	59
rect	253	59	254	60
rect	253	60	254	61
rect	253	61	254	62
rect	253	62	254	63
rect	253	63	254	64
rect	253	64	254	65
rect	253	65	254	66
rect	253	66	254	67
rect	253	67	254	68
rect	253	68	254	69
rect	253	69	254	70
rect	253	70	254	71
rect	253	71	254	72
rect	253	72	254	73
rect	253	73	254	74
rect	253	74	254	75
rect	253	75	254	76
rect	253	76	254	77
rect	253	77	254	78
rect	253	78	254	79
rect	253	79	254	80
rect	253	80	254	81
rect	253	81	254	82
rect	253	82	254	83
rect	253	83	254	84
rect	253	84	254	85
rect	253	85	254	86
rect	253	86	254	87
rect	253	87	254	88
rect	253	88	254	89
rect	253	89	254	90
rect	253	90	254	91
rect	253	91	254	92
rect	253	92	254	93
rect	253	93	254	94
rect	253	94	254	95
rect	253	95	254	96
rect	253	96	254	97
rect	253	97	254	98
rect	253	98	254	99
rect	253	99	254	100
rect	253	100	254	101
rect	253	101	254	102
rect	253	102	254	103
rect	253	103	254	104
rect	253	104	254	105
rect	253	105	254	106
rect	253	106	254	107
rect	253	107	254	108
rect	253	108	254	109
rect	253	109	254	110
rect	253	110	254	111
rect	253	111	254	112
rect	253	112	254	113
rect	253	113	254	114
rect	253	114	254	115
rect	253	115	254	116
rect	253	116	254	117
rect	253	117	254	118
rect	253	118	254	119
rect	253	119	254	120
rect	253	120	254	121
rect	253	121	254	122
rect	253	122	254	123
rect	253	123	254	124
rect	253	124	254	125
rect	253	125	254	126
rect	253	126	254	127
rect	253	127	254	128
rect	253	128	254	129
rect	253	129	254	130
rect	253	130	254	131
rect	253	131	254	132
rect	253	132	254	133
rect	253	133	254	134
rect	253	134	254	135
rect	253	135	254	136
rect	253	136	254	137
rect	253	137	254	138
rect	253	138	254	139
rect	253	139	254	140
rect	253	140	254	141
rect	253	141	254	142
rect	253	142	254	143
rect	253	143	254	144
rect	253	144	254	145
rect	253	145	254	146
rect	253	146	254	147
rect	253	147	254	148
rect	253	148	254	149
rect	253	149	254	150
rect	253	150	254	151
rect	253	151	254	152
rect	253	152	254	153
rect	253	153	254	154
rect	253	154	254	155
rect	253	155	254	156
rect	253	156	254	157
rect	253	157	254	158
rect	253	158	254	159
rect	253	159	254	160
rect	253	160	254	161
rect	253	161	254	162
rect	253	162	254	163
rect	253	163	254	164
rect	253	164	254	165
rect	253	165	254	166
rect	253	166	254	167
rect	253	167	254	168
rect	253	168	254	169
rect	253	169	254	170
rect	253	170	254	171
rect	253	171	254	172
rect	253	172	254	173
rect	253	173	254	174
rect	253	174	254	175
rect	253	175	254	176
rect	253	176	254	177
rect	253	177	254	178
rect	253	178	254	179
rect	253	179	254	180
rect	253	180	254	181
rect	253	181	254	182
rect	253	182	254	183
rect	253	183	254	184
rect	253	184	254	185
rect	253	185	254	186
rect	253	186	254	187
rect	253	187	254	188
rect	253	188	254	189
rect	253	189	254	190
rect	253	190	254	191
rect	253	191	254	192
rect	253	192	254	193
rect	253	193	254	194
rect	253	194	254	195
rect	253	195	254	196
rect	253	196	254	197
rect	253	197	254	198
rect	253	198	254	199
rect	253	199	254	200
rect	253	200	254	201
rect	253	201	254	202
rect	253	202	254	203
rect	253	203	254	204
rect	253	204	254	205
rect	253	205	254	206
rect	253	206	254	207
rect	253	207	254	208
rect	253	208	254	209
rect	253	209	254	210
rect	253	210	254	211
rect	253	211	254	212
rect	253	212	254	213
rect	253	213	254	214
rect	253	214	254	215
rect	253	215	254	216
rect	253	216	254	217
rect	253	217	254	218
rect	253	218	254	219
rect	253	219	254	220
rect	253	220	254	221
rect	253	221	254	222
rect	253	222	254	223
rect	253	223	254	224
rect	253	224	254	225
rect	253	225	254	226
rect	253	226	254	227
rect	253	227	254	228
rect	253	228	254	229
rect	253	229	254	230
rect	253	230	254	231
rect	253	231	254	232
rect	253	232	254	233
rect	253	233	254	234
rect	253	234	254	235
rect	253	235	254	236
rect	253	236	254	237
rect	253	237	254	238
rect	253	238	254	239
rect	253	239	254	240
rect	253	240	254	241
rect	253	241	254	242
rect	253	242	254	243
rect	253	243	254	244
rect	253	244	254	245
rect	253	245	254	246
rect	253	246	254	247
rect	253	247	254	248
rect	253	248	254	249
rect	253	249	254	250
rect	253	250	254	251
rect	253	251	254	252
rect	253	252	254	253
rect	253	253	254	254
rect	253	254	254	255
rect	253	255	254	256
rect	253	256	254	257
rect	253	257	254	258
rect	253	258	254	259
rect	253	259	254	260
rect	253	260	254	261
rect	253	261	254	262
rect	253	262	254	263
rect	253	263	254	264
rect	253	264	254	265
rect	253	265	254	266
rect	253	266	254	267
rect	253	267	254	268
rect	253	268	254	269
rect	253	269	254	270
rect	253	270	254	271
rect	253	271	254	272
rect	253	272	254	273
rect	253	273	254	274
rect	253	274	254	275
rect	253	275	254	276
rect	253	276	254	277
rect	253	277	254	278
rect	253	278	254	279
rect	253	279	254	280
rect	253	280	254	281
rect	253	281	254	282
rect	253	282	254	283
rect	253	283	254	284
rect	253	284	254	285
rect	253	285	254	286
rect	253	286	254	287
rect	253	287	254	288
rect	253	288	254	289
rect	253	289	254	290
rect	253	290	254	291
rect	253	291	254	292
rect	253	292	254	293
rect	253	293	254	294
rect	253	294	254	295
rect	253	295	254	296
rect	253	296	254	297
rect	253	297	254	298
rect	253	298	254	299
rect	253	299	254	300
rect	253	300	254	301
rect	253	301	254	302
rect	253	302	254	303
rect	253	303	254	304
rect	253	304	254	305
rect	253	305	254	306
rect	253	306	254	307
rect	253	307	254	308
rect	253	308	254	309
rect	253	309	254	310
rect	253	310	254	311
rect	253	311	254	312
rect	253	312	254	313
rect	253	313	254	314
rect	253	314	254	315
rect	253	315	254	316
rect	253	316	254	317
rect	253	317	254	318
rect	253	318	254	319
rect	253	319	254	320
rect	253	320	254	321
rect	253	321	254	322
rect	253	322	254	323
rect	253	323	254	324
rect	253	324	254	325
rect	253	325	254	326
rect	253	326	254	327
rect	253	327	254	328
rect	253	328	254	329
rect	253	329	254	330
rect	253	330	254	331
rect	253	331	254	332
rect	253	332	254	333
rect	253	333	254	334
rect	253	334	254	335
rect	253	335	254	336
rect	253	336	254	337
rect	253	337	254	338
rect	253	338	254	339
rect	253	339	254	340
rect	253	340	254	341
rect	253	341	254	342
rect	253	342	254	343
rect	253	343	254	344
rect	253	344	254	345
rect	253	345	254	346
rect	253	346	254	347
rect	253	347	254	348
rect	253	348	254	349
rect	253	349	254	350
rect	253	350	254	351
rect	253	351	254	352
rect	253	352	254	353
rect	253	353	254	354
rect	253	354	254	355
rect	253	355	254	356
rect	253	356	254	357
rect	253	357	254	358
rect	253	358	254	359
rect	253	359	254	360
rect	253	360	254	361
rect	253	361	254	362
rect	253	362	254	363
rect	253	363	254	364
rect	253	364	254	365
rect	253	365	254	366
rect	254	0	255	1
rect	254	1	255	2
rect	254	2	255	3
rect	254	3	255	4
rect	254	4	255	5
rect	254	5	255	6
rect	254	6	255	7
rect	254	7	255	8
rect	254	8	255	9
rect	254	9	255	10
rect	254	10	255	11
rect	254	11	255	12
rect	254	12	255	13
rect	254	13	255	14
rect	254	14	255	15
rect	254	15	255	16
rect	254	16	255	17
rect	254	17	255	18
rect	254	18	255	19
rect	254	19	255	20
rect	254	20	255	21
rect	254	21	255	22
rect	254	22	255	23
rect	254	23	255	24
rect	254	24	255	25
rect	254	25	255	26
rect	254	26	255	27
rect	254	27	255	28
rect	254	28	255	29
rect	254	29	255	30
rect	254	30	255	31
rect	254	31	255	32
rect	254	32	255	33
rect	254	33	255	34
rect	254	34	255	35
rect	254	35	255	36
rect	254	36	255	37
rect	254	37	255	38
rect	254	38	255	39
rect	254	39	255	40
rect	254	40	255	41
rect	254	41	255	42
rect	254	42	255	43
rect	254	43	255	44
rect	254	44	255	45
rect	254	45	255	46
rect	254	46	255	47
rect	254	47	255	48
rect	254	48	255	49
rect	254	49	255	50
rect	254	50	255	51
rect	254	51	255	52
rect	254	52	255	53
rect	254	53	255	54
rect	254	54	255	55
rect	254	55	255	56
rect	254	56	255	57
rect	254	57	255	58
rect	254	58	255	59
rect	254	59	255	60
rect	254	60	255	61
rect	254	61	255	62
rect	254	62	255	63
rect	254	63	255	64
rect	254	64	255	65
rect	254	65	255	66
rect	254	66	255	67
rect	254	67	255	68
rect	254	68	255	69
rect	254	69	255	70
rect	254	70	255	71
rect	254	71	255	72
rect	254	72	255	73
rect	254	73	255	74
rect	254	74	255	75
rect	254	75	255	76
rect	254	76	255	77
rect	254	77	255	78
rect	254	78	255	79
rect	254	79	255	80
rect	254	80	255	81
rect	254	81	255	82
rect	254	82	255	83
rect	254	83	255	84
rect	254	84	255	85
rect	254	85	255	86
rect	254	86	255	87
rect	254	87	255	88
rect	254	88	255	89
rect	254	89	255	90
rect	254	90	255	91
rect	254	91	255	92
rect	254	92	255	93
rect	254	93	255	94
rect	254	94	255	95
rect	254	95	255	96
rect	254	96	255	97
rect	254	97	255	98
rect	254	98	255	99
rect	254	99	255	100
rect	254	100	255	101
rect	254	101	255	102
rect	254	102	255	103
rect	254	103	255	104
rect	254	104	255	105
rect	254	105	255	106
rect	254	106	255	107
rect	254	107	255	108
rect	254	108	255	109
rect	254	109	255	110
rect	254	110	255	111
rect	254	111	255	112
rect	254	112	255	113
rect	254	113	255	114
rect	254	114	255	115
rect	254	115	255	116
rect	254	116	255	117
rect	254	117	255	118
rect	254	118	255	119
rect	254	119	255	120
rect	254	120	255	121
rect	254	121	255	122
rect	254	122	255	123
rect	254	123	255	124
rect	254	124	255	125
rect	254	125	255	126
rect	254	126	255	127
rect	254	127	255	128
rect	254	128	255	129
rect	254	129	255	130
rect	254	130	255	131
rect	254	131	255	132
rect	254	132	255	133
rect	254	133	255	134
rect	254	134	255	135
rect	254	135	255	136
rect	254	136	255	137
rect	254	137	255	138
rect	254	138	255	139
rect	254	139	255	140
rect	254	140	255	141
rect	254	141	255	142
rect	254	142	255	143
rect	254	143	255	144
rect	254	144	255	145
rect	254	145	255	146
rect	254	146	255	147
rect	254	147	255	148
rect	254	148	255	149
rect	254	149	255	150
rect	254	150	255	151
rect	254	151	255	152
rect	254	152	255	153
rect	254	153	255	154
rect	254	154	255	155
rect	254	155	255	156
rect	254	156	255	157
rect	254	157	255	158
rect	254	158	255	159
rect	254	159	255	160
rect	254	160	255	161
rect	254	161	255	162
rect	254	162	255	163
rect	254	163	255	164
rect	254	164	255	165
rect	254	165	255	166
rect	254	166	255	167
rect	254	167	255	168
rect	254	168	255	169
rect	254	169	255	170
rect	254	170	255	171
rect	254	171	255	172
rect	254	172	255	173
rect	254	173	255	174
rect	254	174	255	175
rect	254	175	255	176
rect	254	176	255	177
rect	254	177	255	178
rect	254	178	255	179
rect	254	179	255	180
rect	254	180	255	181
rect	254	181	255	182
rect	254	182	255	183
rect	254	183	255	184
rect	254	184	255	185
rect	254	185	255	186
rect	254	186	255	187
rect	254	187	255	188
rect	254	188	255	189
rect	254	189	255	190
rect	254	190	255	191
rect	254	191	255	192
rect	254	192	255	193
rect	254	193	255	194
rect	254	194	255	195
rect	254	195	255	196
rect	254	196	255	197
rect	254	197	255	198
rect	254	198	255	199
rect	254	199	255	200
rect	254	200	255	201
rect	254	201	255	202
rect	254	202	255	203
rect	254	203	255	204
rect	254	204	255	205
rect	254	205	255	206
rect	254	206	255	207
rect	254	207	255	208
rect	254	208	255	209
rect	254	209	255	210
rect	254	210	255	211
rect	254	211	255	212
rect	254	212	255	213
rect	254	213	255	214
rect	254	214	255	215
rect	254	215	255	216
rect	254	216	255	217
rect	254	217	255	218
rect	254	218	255	219
rect	254	219	255	220
rect	254	220	255	221
rect	254	221	255	222
rect	254	222	255	223
rect	254	223	255	224
rect	254	224	255	225
rect	254	225	255	226
rect	254	226	255	227
rect	254	227	255	228
rect	254	228	255	229
rect	254	229	255	230
rect	254	230	255	231
rect	254	231	255	232
rect	254	232	255	233
rect	254	233	255	234
rect	254	234	255	235
rect	254	235	255	236
rect	254	236	255	237
rect	254	237	255	238
rect	254	238	255	239
rect	254	239	255	240
rect	254	240	255	241
rect	254	241	255	242
rect	254	242	255	243
rect	254	243	255	244
rect	254	244	255	245
rect	254	245	255	246
rect	254	246	255	247
rect	254	247	255	248
rect	254	248	255	249
rect	254	249	255	250
rect	254	250	255	251
rect	254	251	255	252
rect	254	252	255	253
rect	254	253	255	254
rect	254	254	255	255
rect	254	255	255	256
rect	254	256	255	257
rect	254	257	255	258
rect	254	258	255	259
rect	254	259	255	260
rect	254	260	255	261
rect	254	261	255	262
rect	254	262	255	263
rect	254	263	255	264
rect	254	264	255	265
rect	254	265	255	266
rect	254	266	255	267
rect	254	267	255	268
rect	254	268	255	269
rect	254	269	255	270
rect	254	270	255	271
rect	254	271	255	272
rect	254	272	255	273
rect	254	273	255	274
rect	254	274	255	275
rect	254	275	255	276
rect	254	276	255	277
rect	254	277	255	278
rect	254	278	255	279
rect	254	279	255	280
rect	254	280	255	281
rect	254	281	255	282
rect	254	282	255	283
rect	254	283	255	284
rect	254	284	255	285
rect	254	285	255	286
rect	254	286	255	287
rect	254	287	255	288
rect	254	288	255	289
rect	254	289	255	290
rect	254	290	255	291
rect	254	291	255	292
rect	254	292	255	293
rect	254	293	255	294
rect	254	294	255	295
rect	254	295	255	296
rect	254	296	255	297
rect	254	297	255	298
rect	254	298	255	299
rect	254	299	255	300
rect	254	300	255	301
rect	254	301	255	302
rect	254	302	255	303
rect	254	303	255	304
rect	254	304	255	305
rect	254	305	255	306
rect	254	306	255	307
rect	254	307	255	308
rect	254	308	255	309
rect	254	309	255	310
rect	254	310	255	311
rect	254	311	255	312
rect	254	312	255	313
rect	254	313	255	314
rect	254	314	255	315
rect	254	315	255	316
rect	254	316	255	317
rect	254	317	255	318
rect	254	318	255	319
rect	254	319	255	320
rect	254	320	255	321
rect	254	321	255	322
rect	254	322	255	323
rect	254	323	255	324
rect	254	324	255	325
rect	254	325	255	326
rect	254	326	255	327
rect	254	327	255	328
rect	254	328	255	329
rect	254	329	255	330
rect	254	330	255	331
rect	254	331	255	332
rect	254	332	255	333
rect	254	333	255	334
rect	254	334	255	335
rect	254	335	255	336
rect	254	336	255	337
rect	254	337	255	338
rect	254	338	255	339
rect	254	339	255	340
rect	254	340	255	341
rect	254	341	255	342
rect	254	342	255	343
rect	254	343	255	344
rect	254	344	255	345
rect	254	345	255	346
rect	254	346	255	347
rect	254	347	255	348
rect	254	348	255	349
rect	254	349	255	350
rect	254	350	255	351
rect	254	351	255	352
rect	254	352	255	353
rect	254	353	255	354
rect	254	354	255	355
rect	254	355	255	356
rect	254	356	255	357
rect	254	357	255	358
rect	254	358	255	359
rect	254	359	255	360
rect	254	360	255	361
rect	254	361	255	362
rect	254	362	255	363
rect	254	363	255	364
rect	254	364	255	365
rect	254	365	255	366
rect	255	0	256	1
rect	255	1	256	2
rect	255	2	256	3
rect	255	3	256	4
rect	255	4	256	5
rect	255	5	256	6
rect	255	6	256	7
rect	255	7	256	8
rect	255	8	256	9
rect	255	9	256	10
rect	255	10	256	11
rect	255	11	256	12
rect	255	12	256	13
rect	255	13	256	14
rect	255	14	256	15
rect	255	15	256	16
rect	255	16	256	17
rect	255	17	256	18
rect	255	18	256	19
rect	255	19	256	20
rect	255	20	256	21
rect	255	21	256	22
rect	255	22	256	23
rect	255	23	256	24
rect	255	24	256	25
rect	255	25	256	26
rect	255	26	256	27
rect	255	27	256	28
rect	255	28	256	29
rect	255	29	256	30
rect	255	30	256	31
rect	255	31	256	32
rect	255	32	256	33
rect	255	33	256	34
rect	255	34	256	35
rect	255	35	256	36
rect	255	36	256	37
rect	255	37	256	38
rect	255	38	256	39
rect	255	39	256	40
rect	255	40	256	41
rect	255	41	256	42
rect	255	42	256	43
rect	255	43	256	44
rect	255	44	256	45
rect	255	45	256	46
rect	255	46	256	47
rect	255	47	256	48
rect	255	48	256	49
rect	255	49	256	50
rect	255	50	256	51
rect	255	51	256	52
rect	255	52	256	53
rect	255	53	256	54
rect	255	54	256	55
rect	255	55	256	56
rect	255	56	256	57
rect	255	57	256	58
rect	255	58	256	59
rect	255	59	256	60
rect	255	60	256	61
rect	255	61	256	62
rect	255	62	256	63
rect	255	63	256	64
rect	255	64	256	65
rect	255	65	256	66
rect	255	66	256	67
rect	255	67	256	68
rect	255	68	256	69
rect	255	69	256	70
rect	255	70	256	71
rect	255	71	256	72
rect	255	72	256	73
rect	255	73	256	74
rect	255	74	256	75
rect	255	75	256	76
rect	255	76	256	77
rect	255	77	256	78
rect	255	78	256	79
rect	255	79	256	80
rect	255	80	256	81
rect	255	81	256	82
rect	255	82	256	83
rect	255	83	256	84
rect	255	84	256	85
rect	255	85	256	86
rect	255	86	256	87
rect	255	87	256	88
rect	255	88	256	89
rect	255	89	256	90
rect	255	90	256	91
rect	255	91	256	92
rect	255	92	256	93
rect	255	93	256	94
rect	255	94	256	95
rect	255	95	256	96
rect	255	96	256	97
rect	255	97	256	98
rect	255	98	256	99
rect	255	99	256	100
rect	255	100	256	101
rect	255	101	256	102
rect	255	102	256	103
rect	255	103	256	104
rect	255	104	256	105
rect	255	105	256	106
rect	255	106	256	107
rect	255	107	256	108
rect	255	108	256	109
rect	255	109	256	110
rect	255	110	256	111
rect	255	111	256	112
rect	255	112	256	113
rect	255	113	256	114
rect	255	114	256	115
rect	255	115	256	116
rect	255	116	256	117
rect	255	117	256	118
rect	255	118	256	119
rect	255	119	256	120
rect	255	120	256	121
rect	255	121	256	122
rect	255	122	256	123
rect	255	123	256	124
rect	255	124	256	125
rect	255	125	256	126
rect	255	126	256	127
rect	255	127	256	128
rect	255	128	256	129
rect	255	129	256	130
rect	255	130	256	131
rect	255	131	256	132
rect	255	132	256	133
rect	255	133	256	134
rect	255	134	256	135
rect	255	135	256	136
rect	255	136	256	137
rect	255	137	256	138
rect	255	138	256	139
rect	255	139	256	140
rect	255	140	256	141
rect	255	141	256	142
rect	255	142	256	143
rect	255	143	256	144
rect	255	144	256	145
rect	255	145	256	146
rect	255	146	256	147
rect	255	147	256	148
rect	255	148	256	149
rect	255	149	256	150
rect	255	150	256	151
rect	255	151	256	152
rect	255	152	256	153
rect	255	153	256	154
rect	255	154	256	155
rect	255	155	256	156
rect	255	156	256	157
rect	255	157	256	158
rect	255	158	256	159
rect	255	159	256	160
rect	255	160	256	161
rect	255	161	256	162
rect	255	162	256	163
rect	255	163	256	164
rect	255	164	256	165
rect	255	165	256	166
rect	255	166	256	167
rect	255	167	256	168
rect	255	168	256	169
rect	255	169	256	170
rect	255	170	256	171
rect	255	171	256	172
rect	255	172	256	173
rect	255	173	256	174
rect	255	174	256	175
rect	255	175	256	176
rect	255	176	256	177
rect	255	177	256	178
rect	255	178	256	179
rect	255	179	256	180
rect	255	180	256	181
rect	255	181	256	182
rect	255	182	256	183
rect	255	183	256	184
rect	255	184	256	185
rect	255	185	256	186
rect	255	186	256	187
rect	255	187	256	188
rect	255	188	256	189
rect	255	189	256	190
rect	255	190	256	191
rect	255	191	256	192
rect	255	192	256	193
rect	255	193	256	194
rect	255	194	256	195
rect	255	195	256	196
rect	255	196	256	197
rect	255	197	256	198
rect	255	198	256	199
rect	255	199	256	200
rect	255	200	256	201
rect	255	201	256	202
rect	255	202	256	203
rect	255	203	256	204
rect	255	204	256	205
rect	255	205	256	206
rect	255	206	256	207
rect	255	207	256	208
rect	255	208	256	209
rect	255	209	256	210
rect	255	210	256	211
rect	255	211	256	212
rect	255	212	256	213
rect	255	213	256	214
rect	255	214	256	215
rect	255	215	256	216
rect	255	216	256	217
rect	255	217	256	218
rect	255	218	256	219
rect	255	219	256	220
rect	255	220	256	221
rect	255	221	256	222
rect	255	222	256	223
rect	255	223	256	224
rect	255	224	256	225
rect	255	225	256	226
rect	255	226	256	227
rect	255	227	256	228
rect	255	228	256	229
rect	255	229	256	230
rect	255	230	256	231
rect	255	231	256	232
rect	255	232	256	233
rect	255	233	256	234
rect	255	234	256	235
rect	255	235	256	236
rect	255	236	256	237
rect	255	237	256	238
rect	255	238	256	239
rect	255	239	256	240
rect	255	240	256	241
rect	255	241	256	242
rect	255	242	256	243
rect	255	243	256	244
rect	255	244	256	245
rect	255	245	256	246
rect	255	246	256	247
rect	255	247	256	248
rect	255	248	256	249
rect	255	249	256	250
rect	255	250	256	251
rect	255	251	256	252
rect	255	252	256	253
rect	255	253	256	254
rect	255	254	256	255
rect	255	255	256	256
rect	255	256	256	257
rect	255	257	256	258
rect	255	258	256	259
rect	255	259	256	260
rect	255	260	256	261
rect	255	261	256	262
rect	255	262	256	263
rect	255	263	256	264
rect	255	264	256	265
rect	255	265	256	266
rect	255	266	256	267
rect	255	267	256	268
rect	255	268	256	269
rect	255	269	256	270
rect	255	270	256	271
rect	255	271	256	272
rect	255	272	256	273
rect	255	273	256	274
rect	255	274	256	275
rect	255	275	256	276
rect	255	276	256	277
rect	255	277	256	278
rect	255	278	256	279
rect	255	279	256	280
rect	255	280	256	281
rect	255	281	256	282
rect	255	282	256	283
rect	255	283	256	284
rect	255	284	256	285
rect	255	285	256	286
rect	255	286	256	287
rect	255	287	256	288
rect	255	288	256	289
rect	255	289	256	290
rect	255	290	256	291
rect	255	291	256	292
rect	255	292	256	293
rect	255	293	256	294
rect	255	294	256	295
rect	255	295	256	296
rect	255	296	256	297
rect	255	297	256	298
rect	255	298	256	299
rect	255	299	256	300
rect	255	300	256	301
rect	255	301	256	302
rect	255	302	256	303
rect	255	303	256	304
rect	255	304	256	305
rect	255	305	256	306
rect	255	306	256	307
rect	255	307	256	308
rect	255	308	256	309
rect	255	309	256	310
rect	255	310	256	311
rect	255	311	256	312
rect	255	312	256	313
rect	255	313	256	314
rect	255	314	256	315
rect	255	315	256	316
rect	255	316	256	317
rect	255	317	256	318
rect	255	318	256	319
rect	255	319	256	320
rect	255	320	256	321
rect	255	321	256	322
rect	255	322	256	323
rect	255	323	256	324
rect	255	324	256	325
rect	255	325	256	326
rect	255	326	256	327
rect	255	327	256	328
rect	255	328	256	329
rect	255	329	256	330
rect	255	330	256	331
rect	255	331	256	332
rect	255	332	256	333
rect	255	333	256	334
rect	255	334	256	335
rect	255	335	256	336
rect	255	336	256	337
rect	255	337	256	338
rect	255	338	256	339
rect	255	339	256	340
rect	255	340	256	341
rect	255	341	256	342
rect	255	342	256	343
rect	255	343	256	344
rect	255	344	256	345
rect	255	345	256	346
rect	255	346	256	347
rect	255	347	256	348
rect	255	348	256	349
rect	255	349	256	350
rect	255	350	256	351
rect	255	351	256	352
rect	255	352	256	353
rect	255	353	256	354
rect	255	354	256	355
rect	255	355	256	356
rect	255	356	256	357
rect	255	357	256	358
rect	255	358	256	359
rect	255	359	256	360
rect	255	360	256	361
rect	255	361	256	362
rect	255	362	256	363
rect	255	363	256	364
rect	255	364	256	365
rect	255	365	256	366
rect	256	0	257	1
rect	256	1	257	2
rect	256	2	257	3
rect	256	3	257	4
rect	256	4	257	5
rect	256	5	257	6
rect	256	6	257	7
rect	256	7	257	8
rect	256	8	257	9
rect	256	9	257	10
rect	256	10	257	11
rect	256	11	257	12
rect	256	12	257	13
rect	256	13	257	14
rect	256	14	257	15
rect	256	15	257	16
rect	256	16	257	17
rect	256	17	257	18
rect	256	18	257	19
rect	256	19	257	20
rect	256	20	257	21
rect	256	21	257	22
rect	256	22	257	23
rect	256	23	257	24
rect	256	24	257	25
rect	256	25	257	26
rect	256	26	257	27
rect	256	27	257	28
rect	256	28	257	29
rect	256	29	257	30
rect	256	30	257	31
rect	256	31	257	32
rect	256	32	257	33
rect	256	33	257	34
rect	256	34	257	35
rect	256	35	257	36
rect	256	36	257	37
rect	256	37	257	38
rect	256	38	257	39
rect	256	39	257	40
rect	256	40	257	41
rect	256	41	257	42
rect	256	42	257	43
rect	256	43	257	44
rect	256	44	257	45
rect	256	45	257	46
rect	256	46	257	47
rect	256	47	257	48
rect	256	48	257	49
rect	256	49	257	50
rect	256	50	257	51
rect	256	51	257	52
rect	256	52	257	53
rect	256	53	257	54
rect	256	54	257	55
rect	256	55	257	56
rect	256	56	257	57
rect	256	57	257	58
rect	256	58	257	59
rect	256	59	257	60
rect	256	60	257	61
rect	256	61	257	62
rect	256	62	257	63
rect	256	63	257	64
rect	256	64	257	65
rect	256	65	257	66
rect	256	66	257	67
rect	256	67	257	68
rect	256	68	257	69
rect	256	69	257	70
rect	256	70	257	71
rect	256	71	257	72
rect	256	72	257	73
rect	256	73	257	74
rect	256	74	257	75
rect	256	75	257	76
rect	256	76	257	77
rect	256	77	257	78
rect	256	78	257	79
rect	256	79	257	80
rect	256	80	257	81
rect	256	81	257	82
rect	256	82	257	83
rect	256	83	257	84
rect	256	84	257	85
rect	256	85	257	86
rect	256	86	257	87
rect	256	87	257	88
rect	256	88	257	89
rect	256	89	257	90
rect	256	90	257	91
rect	256	91	257	92
rect	256	92	257	93
rect	256	93	257	94
rect	256	94	257	95
rect	256	95	257	96
rect	256	96	257	97
rect	256	97	257	98
rect	256	98	257	99
rect	256	99	257	100
rect	256	100	257	101
rect	256	101	257	102
rect	256	102	257	103
rect	256	103	257	104
rect	256	104	257	105
rect	256	105	257	106
rect	256	106	257	107
rect	256	107	257	108
rect	256	108	257	109
rect	256	109	257	110
rect	256	110	257	111
rect	256	111	257	112
rect	256	112	257	113
rect	256	113	257	114
rect	256	114	257	115
rect	256	115	257	116
rect	256	116	257	117
rect	256	117	257	118
rect	256	118	257	119
rect	256	119	257	120
rect	256	120	257	121
rect	256	121	257	122
rect	256	122	257	123
rect	256	123	257	124
rect	256	124	257	125
rect	256	125	257	126
rect	256	126	257	127
rect	256	127	257	128
rect	256	128	257	129
rect	256	129	257	130
rect	256	130	257	131
rect	256	131	257	132
rect	256	132	257	133
rect	256	133	257	134
rect	256	134	257	135
rect	256	135	257	136
rect	256	136	257	137
rect	256	137	257	138
rect	256	138	257	139
rect	256	139	257	140
rect	256	140	257	141
rect	256	141	257	142
rect	256	142	257	143
rect	256	143	257	144
rect	256	144	257	145
rect	256	145	257	146
rect	256	146	257	147
rect	256	147	257	148
rect	256	148	257	149
rect	256	149	257	150
rect	256	150	257	151
rect	256	151	257	152
rect	256	152	257	153
rect	256	153	257	154
rect	256	154	257	155
rect	256	155	257	156
rect	256	156	257	157
rect	256	157	257	158
rect	256	158	257	159
rect	256	159	257	160
rect	256	160	257	161
rect	256	161	257	162
rect	256	162	257	163
rect	256	163	257	164
rect	256	164	257	165
rect	256	165	257	166
rect	256	166	257	167
rect	256	167	257	168
rect	256	168	257	169
rect	256	169	257	170
rect	256	170	257	171
rect	256	171	257	172
rect	256	172	257	173
rect	256	173	257	174
rect	256	174	257	175
rect	256	175	257	176
rect	256	176	257	177
rect	256	177	257	178
rect	256	178	257	179
rect	256	179	257	180
rect	256	180	257	181
rect	256	181	257	182
rect	256	182	257	183
rect	256	183	257	184
rect	256	184	257	185
rect	256	185	257	186
rect	256	186	257	187
rect	256	187	257	188
rect	256	188	257	189
rect	256	189	257	190
rect	256	190	257	191
rect	256	191	257	192
rect	256	192	257	193
rect	256	193	257	194
rect	256	194	257	195
rect	256	195	257	196
rect	256	196	257	197
rect	256	197	257	198
rect	256	198	257	199
rect	256	199	257	200
rect	256	200	257	201
rect	256	201	257	202
rect	256	202	257	203
rect	256	203	257	204
rect	256	204	257	205
rect	256	205	257	206
rect	256	206	257	207
rect	256	207	257	208
rect	256	208	257	209
rect	256	209	257	210
rect	256	210	257	211
rect	256	211	257	212
rect	256	212	257	213
rect	256	213	257	214
rect	256	214	257	215
rect	256	215	257	216
rect	256	216	257	217
rect	256	217	257	218
rect	256	218	257	219
rect	256	219	257	220
rect	256	220	257	221
rect	256	221	257	222
rect	256	222	257	223
rect	256	223	257	224
rect	256	224	257	225
rect	256	225	257	226
rect	256	226	257	227
rect	256	227	257	228
rect	256	228	257	229
rect	256	229	257	230
rect	256	230	257	231
rect	256	231	257	232
rect	256	232	257	233
rect	256	233	257	234
rect	256	234	257	235
rect	256	235	257	236
rect	256	236	257	237
rect	256	237	257	238
rect	256	238	257	239
rect	256	239	257	240
rect	256	240	257	241
rect	256	241	257	242
rect	256	242	257	243
rect	256	243	257	244
rect	256	244	257	245
rect	256	245	257	246
rect	256	246	257	247
rect	256	247	257	248
rect	256	248	257	249
rect	256	249	257	250
rect	256	250	257	251
rect	256	251	257	252
rect	256	252	257	253
rect	256	253	257	254
rect	256	254	257	255
rect	256	255	257	256
rect	256	256	257	257
rect	256	257	257	258
rect	256	258	257	259
rect	256	259	257	260
rect	256	260	257	261
rect	256	261	257	262
rect	256	262	257	263
rect	256	263	257	264
rect	256	264	257	265
rect	256	265	257	266
rect	256	266	257	267
rect	256	267	257	268
rect	256	268	257	269
rect	256	269	257	270
rect	256	270	257	271
rect	256	271	257	272
rect	256	272	257	273
rect	256	273	257	274
rect	256	274	257	275
rect	256	275	257	276
rect	256	276	257	277
rect	256	277	257	278
rect	256	278	257	279
rect	256	279	257	280
rect	256	280	257	281
rect	256	281	257	282
rect	256	282	257	283
rect	256	283	257	284
rect	256	284	257	285
rect	256	285	257	286
rect	256	286	257	287
rect	256	287	257	288
rect	256	288	257	289
rect	256	289	257	290
rect	256	290	257	291
rect	256	291	257	292
rect	256	292	257	293
rect	256	293	257	294
rect	256	294	257	295
rect	256	295	257	296
rect	256	296	257	297
rect	256	297	257	298
rect	256	298	257	299
rect	256	299	257	300
rect	256	300	257	301
rect	256	301	257	302
rect	256	302	257	303
rect	256	303	257	304
rect	256	304	257	305
rect	256	305	257	306
rect	256	306	257	307
rect	256	307	257	308
rect	256	308	257	309
rect	256	309	257	310
rect	256	310	257	311
rect	256	311	257	312
rect	256	312	257	313
rect	256	313	257	314
rect	256	314	257	315
rect	256	315	257	316
rect	256	316	257	317
rect	256	317	257	318
rect	256	318	257	319
rect	256	319	257	320
rect	256	320	257	321
rect	256	321	257	322
rect	256	322	257	323
rect	256	323	257	324
rect	256	324	257	325
rect	256	325	257	326
rect	256	326	257	327
rect	256	327	257	328
rect	256	328	257	329
rect	256	329	257	330
rect	256	330	257	331
rect	256	331	257	332
rect	256	332	257	333
rect	256	333	257	334
rect	256	334	257	335
rect	256	335	257	336
rect	256	336	257	337
rect	256	337	257	338
rect	256	338	257	339
rect	256	339	257	340
rect	256	340	257	341
rect	256	341	257	342
rect	256	342	257	343
rect	256	343	257	344
rect	256	344	257	345
rect	256	345	257	346
rect	256	346	257	347
rect	256	347	257	348
rect	256	348	257	349
rect	256	349	257	350
rect	256	350	257	351
rect	256	351	257	352
rect	256	352	257	353
rect	256	353	257	354
rect	256	354	257	355
rect	256	355	257	356
rect	256	356	257	357
rect	256	357	257	358
rect	256	358	257	359
rect	256	359	257	360
rect	256	360	257	361
rect	256	361	257	362
rect	256	362	257	363
rect	256	363	257	364
rect	256	364	257	365
rect	256	365	257	366
rect	257	0	258	1
rect	257	1	258	2
rect	257	2	258	3
rect	257	3	258	4
rect	257	4	258	5
rect	257	5	258	6
rect	257	6	258	7
rect	257	7	258	8
rect	257	8	258	9
rect	257	9	258	10
rect	257	10	258	11
rect	257	11	258	12
rect	257	12	258	13
rect	257	13	258	14
rect	257	14	258	15
rect	257	15	258	16
rect	257	16	258	17
rect	257	17	258	18
rect	257	18	258	19
rect	257	19	258	20
rect	257	20	258	21
rect	257	21	258	22
rect	257	22	258	23
rect	257	23	258	24
rect	257	24	258	25
rect	257	25	258	26
rect	257	26	258	27
rect	257	27	258	28
rect	257	28	258	29
rect	257	29	258	30
rect	257	30	258	31
rect	257	31	258	32
rect	257	32	258	33
rect	257	33	258	34
rect	257	34	258	35
rect	257	35	258	36
rect	257	36	258	37
rect	257	37	258	38
rect	257	38	258	39
rect	257	39	258	40
rect	257	40	258	41
rect	257	41	258	42
rect	257	42	258	43
rect	257	43	258	44
rect	257	44	258	45
rect	257	45	258	46
rect	257	46	258	47
rect	257	47	258	48
rect	257	48	258	49
rect	257	49	258	50
rect	257	50	258	51
rect	257	51	258	52
rect	257	52	258	53
rect	257	53	258	54
rect	257	54	258	55
rect	257	55	258	56
rect	257	56	258	57
rect	257	57	258	58
rect	257	58	258	59
rect	257	59	258	60
rect	257	60	258	61
rect	257	61	258	62
rect	257	62	258	63
rect	257	63	258	64
rect	257	64	258	65
rect	257	65	258	66
rect	257	66	258	67
rect	257	67	258	68
rect	257	68	258	69
rect	257	69	258	70
rect	257	70	258	71
rect	257	71	258	72
rect	257	72	258	73
rect	257	73	258	74
rect	257	74	258	75
rect	257	75	258	76
rect	257	76	258	77
rect	257	77	258	78
rect	257	78	258	79
rect	257	79	258	80
rect	257	80	258	81
rect	257	81	258	82
rect	257	82	258	83
rect	257	83	258	84
rect	257	84	258	85
rect	257	85	258	86
rect	257	86	258	87
rect	257	87	258	88
rect	257	88	258	89
rect	257	89	258	90
rect	257	90	258	91
rect	257	91	258	92
rect	257	92	258	93
rect	257	93	258	94
rect	257	94	258	95
rect	257	95	258	96
rect	257	96	258	97
rect	257	97	258	98
rect	257	98	258	99
rect	257	99	258	100
rect	257	100	258	101
rect	257	101	258	102
rect	257	102	258	103
rect	257	103	258	104
rect	257	104	258	105
rect	257	105	258	106
rect	257	106	258	107
rect	257	107	258	108
rect	257	108	258	109
rect	257	109	258	110
rect	257	110	258	111
rect	257	111	258	112
rect	257	112	258	113
rect	257	113	258	114
rect	257	114	258	115
rect	257	115	258	116
rect	257	116	258	117
rect	257	117	258	118
rect	257	118	258	119
rect	257	119	258	120
rect	257	120	258	121
rect	257	121	258	122
rect	257	122	258	123
rect	257	123	258	124
rect	257	124	258	125
rect	257	125	258	126
rect	257	126	258	127
rect	257	127	258	128
rect	257	128	258	129
rect	257	129	258	130
rect	257	130	258	131
rect	257	131	258	132
rect	257	132	258	133
rect	257	133	258	134
rect	257	134	258	135
rect	257	135	258	136
rect	257	136	258	137
rect	257	137	258	138
rect	257	138	258	139
rect	257	139	258	140
rect	257	140	258	141
rect	257	141	258	142
rect	257	142	258	143
rect	257	143	258	144
rect	257	144	258	145
rect	257	145	258	146
rect	257	146	258	147
rect	257	147	258	148
rect	257	148	258	149
rect	257	149	258	150
rect	257	150	258	151
rect	257	151	258	152
rect	257	152	258	153
rect	257	153	258	154
rect	257	154	258	155
rect	257	155	258	156
rect	257	156	258	157
rect	257	157	258	158
rect	257	158	258	159
rect	257	159	258	160
rect	257	160	258	161
rect	257	161	258	162
rect	257	162	258	163
rect	257	163	258	164
rect	257	164	258	165
rect	257	165	258	166
rect	257	166	258	167
rect	257	167	258	168
rect	257	168	258	169
rect	257	169	258	170
rect	257	170	258	171
rect	257	171	258	172
rect	257	172	258	173
rect	257	173	258	174
rect	257	174	258	175
rect	257	175	258	176
rect	257	176	258	177
rect	257	177	258	178
rect	257	178	258	179
rect	257	179	258	180
rect	257	180	258	181
rect	257	181	258	182
rect	257	182	258	183
rect	257	183	258	184
rect	257	184	258	185
rect	257	185	258	186
rect	257	186	258	187
rect	257	187	258	188
rect	257	188	258	189
rect	257	189	258	190
rect	257	190	258	191
rect	257	191	258	192
rect	257	192	258	193
rect	257	193	258	194
rect	257	194	258	195
rect	257	195	258	196
rect	257	196	258	197
rect	257	197	258	198
rect	257	198	258	199
rect	257	199	258	200
rect	257	200	258	201
rect	257	201	258	202
rect	257	202	258	203
rect	257	203	258	204
rect	257	204	258	205
rect	257	205	258	206
rect	257	206	258	207
rect	257	207	258	208
rect	257	208	258	209
rect	257	209	258	210
rect	257	210	258	211
rect	257	211	258	212
rect	257	212	258	213
rect	257	213	258	214
rect	257	214	258	215
rect	257	215	258	216
rect	257	216	258	217
rect	257	217	258	218
rect	257	218	258	219
rect	257	219	258	220
rect	257	220	258	221
rect	257	221	258	222
rect	257	222	258	223
rect	257	223	258	224
rect	257	224	258	225
rect	257	225	258	226
rect	257	226	258	227
rect	257	227	258	228
rect	257	228	258	229
rect	257	229	258	230
rect	257	230	258	231
rect	257	231	258	232
rect	257	232	258	233
rect	257	233	258	234
rect	257	234	258	235
rect	257	235	258	236
rect	257	236	258	237
rect	257	237	258	238
rect	257	238	258	239
rect	257	239	258	240
rect	257	240	258	241
rect	257	241	258	242
rect	257	242	258	243
rect	257	243	258	244
rect	257	244	258	245
rect	257	245	258	246
rect	257	246	258	247
rect	257	247	258	248
rect	257	248	258	249
rect	257	249	258	250
rect	257	250	258	251
rect	257	251	258	252
rect	257	252	258	253
rect	257	253	258	254
rect	257	254	258	255
rect	257	255	258	256
rect	257	256	258	257
rect	257	257	258	258
rect	257	258	258	259
rect	257	259	258	260
rect	257	260	258	261
rect	257	261	258	262
rect	257	262	258	263
rect	257	263	258	264
rect	257	264	258	265
rect	257	265	258	266
rect	257	266	258	267
rect	257	267	258	268
rect	257	268	258	269
rect	257	269	258	270
rect	257	270	258	271
rect	257	271	258	272
rect	257	272	258	273
rect	257	273	258	274
rect	257	274	258	275
rect	257	275	258	276
rect	257	276	258	277
rect	257	277	258	278
rect	257	278	258	279
rect	257	279	258	280
rect	257	280	258	281
rect	257	281	258	282
rect	257	282	258	283
rect	257	283	258	284
rect	257	284	258	285
rect	257	285	258	286
rect	257	286	258	287
rect	257	287	258	288
rect	257	288	258	289
rect	257	289	258	290
rect	257	290	258	291
rect	257	291	258	292
rect	257	292	258	293
rect	257	293	258	294
rect	257	294	258	295
rect	257	295	258	296
rect	257	296	258	297
rect	257	297	258	298
rect	257	298	258	299
rect	257	299	258	300
rect	257	300	258	301
rect	257	301	258	302
rect	257	302	258	303
rect	257	303	258	304
rect	257	304	258	305
rect	257	305	258	306
rect	257	306	258	307
rect	257	307	258	308
rect	257	308	258	309
rect	257	309	258	310
rect	257	310	258	311
rect	257	311	258	312
rect	257	312	258	313
rect	257	313	258	314
rect	257	314	258	315
rect	257	315	258	316
rect	257	316	258	317
rect	257	317	258	318
rect	257	318	258	319
rect	257	319	258	320
rect	257	320	258	321
rect	257	321	258	322
rect	257	322	258	323
rect	257	323	258	324
rect	257	324	258	325
rect	257	325	258	326
rect	257	326	258	327
rect	257	327	258	328
rect	257	328	258	329
rect	257	329	258	330
rect	257	330	258	331
rect	257	331	258	332
rect	257	332	258	333
rect	257	333	258	334
rect	257	334	258	335
rect	257	335	258	336
rect	257	336	258	337
rect	257	337	258	338
rect	257	338	258	339
rect	257	339	258	340
rect	257	340	258	341
rect	257	341	258	342
rect	257	342	258	343
rect	257	343	258	344
rect	257	344	258	345
rect	257	345	258	346
rect	257	346	258	347
rect	257	347	258	348
rect	257	348	258	349
rect	257	349	258	350
rect	257	350	258	351
rect	257	351	258	352
rect	257	352	258	353
rect	257	353	258	354
rect	257	354	258	355
rect	257	355	258	356
rect	257	356	258	357
rect	257	357	258	358
rect	257	358	258	359
rect	257	359	258	360
rect	257	360	258	361
rect	257	361	258	362
rect	257	362	258	363
rect	257	363	258	364
rect	257	364	258	365
rect	257	365	258	366
rect	258	0	259	1
rect	258	1	259	2
rect	258	2	259	3
rect	258	3	259	4
rect	258	4	259	5
rect	258	5	259	6
rect	258	6	259	7
rect	258	7	259	8
rect	258	8	259	9
rect	258	9	259	10
rect	258	10	259	11
rect	258	11	259	12
rect	258	12	259	13
rect	258	13	259	14
rect	258	14	259	15
rect	258	15	259	16
rect	258	16	259	17
rect	258	17	259	18
rect	258	18	259	19
rect	258	19	259	20
rect	258	20	259	21
rect	258	21	259	22
rect	258	22	259	23
rect	258	23	259	24
rect	258	24	259	25
rect	258	25	259	26
rect	258	26	259	27
rect	258	27	259	28
rect	258	28	259	29
rect	258	29	259	30
rect	258	30	259	31
rect	258	31	259	32
rect	258	32	259	33
rect	258	33	259	34
rect	258	34	259	35
rect	258	35	259	36
rect	258	36	259	37
rect	258	37	259	38
rect	258	38	259	39
rect	258	39	259	40
rect	258	40	259	41
rect	258	41	259	42
rect	258	42	259	43
rect	258	43	259	44
rect	258	44	259	45
rect	258	45	259	46
rect	258	46	259	47
rect	258	47	259	48
rect	258	48	259	49
rect	258	49	259	50
rect	258	50	259	51
rect	258	51	259	52
rect	258	52	259	53
rect	258	53	259	54
rect	258	54	259	55
rect	258	55	259	56
rect	258	56	259	57
rect	258	57	259	58
rect	258	58	259	59
rect	258	59	259	60
rect	258	60	259	61
rect	258	61	259	62
rect	258	62	259	63
rect	258	63	259	64
rect	258	64	259	65
rect	258	65	259	66
rect	258	66	259	67
rect	258	67	259	68
rect	258	68	259	69
rect	258	69	259	70
rect	258	70	259	71
rect	258	71	259	72
rect	258	72	259	73
rect	258	73	259	74
rect	258	74	259	75
rect	258	75	259	76
rect	258	76	259	77
rect	258	77	259	78
rect	258	78	259	79
rect	258	79	259	80
rect	258	80	259	81
rect	258	81	259	82
rect	258	82	259	83
rect	258	83	259	84
rect	258	84	259	85
rect	258	85	259	86
rect	258	86	259	87
rect	258	87	259	88
rect	258	88	259	89
rect	258	89	259	90
rect	258	90	259	91
rect	258	91	259	92
rect	258	92	259	93
rect	258	93	259	94
rect	258	94	259	95
rect	258	95	259	96
rect	258	96	259	97
rect	258	97	259	98
rect	258	98	259	99
rect	258	99	259	100
rect	258	100	259	101
rect	258	101	259	102
rect	258	102	259	103
rect	258	103	259	104
rect	258	104	259	105
rect	258	105	259	106
rect	258	106	259	107
rect	258	107	259	108
rect	258	108	259	109
rect	258	109	259	110
rect	258	110	259	111
rect	258	111	259	112
rect	258	112	259	113
rect	258	113	259	114
rect	258	114	259	115
rect	258	115	259	116
rect	258	116	259	117
rect	258	117	259	118
rect	258	118	259	119
rect	258	119	259	120
rect	258	120	259	121
rect	258	121	259	122
rect	258	122	259	123
rect	258	123	259	124
rect	258	124	259	125
rect	258	125	259	126
rect	258	126	259	127
rect	258	127	259	128
rect	258	128	259	129
rect	258	129	259	130
rect	258	130	259	131
rect	258	131	259	132
rect	258	132	259	133
rect	258	133	259	134
rect	258	134	259	135
rect	258	135	259	136
rect	258	136	259	137
rect	258	137	259	138
rect	258	138	259	139
rect	258	139	259	140
rect	258	140	259	141
rect	258	141	259	142
rect	258	142	259	143
rect	258	143	259	144
rect	258	144	259	145
rect	258	145	259	146
rect	258	146	259	147
rect	258	147	259	148
rect	258	148	259	149
rect	258	149	259	150
rect	258	150	259	151
rect	258	151	259	152
rect	258	152	259	153
rect	258	153	259	154
rect	258	154	259	155
rect	258	155	259	156
rect	258	156	259	157
rect	258	157	259	158
rect	258	158	259	159
rect	258	159	259	160
rect	258	160	259	161
rect	258	161	259	162
rect	258	162	259	163
rect	258	163	259	164
rect	258	164	259	165
rect	258	165	259	166
rect	258	166	259	167
rect	258	167	259	168
rect	258	168	259	169
rect	258	169	259	170
rect	258	170	259	171
rect	258	171	259	172
rect	258	172	259	173
rect	258	173	259	174
rect	258	174	259	175
rect	258	175	259	176
rect	258	176	259	177
rect	258	177	259	178
rect	258	178	259	179
rect	258	179	259	180
rect	258	180	259	181
rect	258	181	259	182
rect	258	182	259	183
rect	258	183	259	184
rect	258	184	259	185
rect	258	185	259	186
rect	258	186	259	187
rect	258	187	259	188
rect	258	188	259	189
rect	258	189	259	190
rect	258	190	259	191
rect	258	191	259	192
rect	258	192	259	193
rect	258	193	259	194
rect	258	194	259	195
rect	258	195	259	196
rect	258	196	259	197
rect	258	197	259	198
rect	258	198	259	199
rect	258	199	259	200
rect	258	200	259	201
rect	258	201	259	202
rect	258	202	259	203
rect	258	203	259	204
rect	258	204	259	205
rect	258	205	259	206
rect	258	206	259	207
rect	258	207	259	208
rect	258	208	259	209
rect	258	209	259	210
rect	258	210	259	211
rect	258	211	259	212
rect	258	212	259	213
rect	258	213	259	214
rect	258	214	259	215
rect	258	215	259	216
rect	258	216	259	217
rect	258	217	259	218
rect	258	218	259	219
rect	258	219	259	220
rect	258	220	259	221
rect	258	221	259	222
rect	258	222	259	223
rect	258	223	259	224
rect	258	224	259	225
rect	258	225	259	226
rect	258	226	259	227
rect	258	227	259	228
rect	258	228	259	229
rect	258	229	259	230
rect	258	230	259	231
rect	258	231	259	232
rect	258	232	259	233
rect	258	233	259	234
rect	258	234	259	235
rect	258	235	259	236
rect	258	236	259	237
rect	258	237	259	238
rect	258	238	259	239
rect	258	239	259	240
rect	258	240	259	241
rect	258	241	259	242
rect	258	242	259	243
rect	258	243	259	244
rect	258	244	259	245
rect	258	245	259	246
rect	258	246	259	247
rect	258	247	259	248
rect	258	248	259	249
rect	258	249	259	250
rect	258	250	259	251
rect	258	251	259	252
rect	258	252	259	253
rect	258	253	259	254
rect	258	254	259	255
rect	258	255	259	256
rect	258	256	259	257
rect	258	257	259	258
rect	258	258	259	259
rect	258	259	259	260
rect	258	260	259	261
rect	258	261	259	262
rect	258	262	259	263
rect	258	263	259	264
rect	258	264	259	265
rect	258	265	259	266
rect	258	266	259	267
rect	258	267	259	268
rect	258	268	259	269
rect	258	269	259	270
rect	258	270	259	271
rect	258	271	259	272
rect	258	272	259	273
rect	258	273	259	274
rect	258	274	259	275
rect	258	275	259	276
rect	258	276	259	277
rect	258	277	259	278
rect	258	278	259	279
rect	258	279	259	280
rect	258	280	259	281
rect	258	281	259	282
rect	258	282	259	283
rect	258	283	259	284
rect	258	284	259	285
rect	258	285	259	286
rect	258	286	259	287
rect	258	287	259	288
rect	258	288	259	289
rect	258	289	259	290
rect	258	290	259	291
rect	258	291	259	292
rect	258	292	259	293
rect	258	293	259	294
rect	258	294	259	295
rect	258	295	259	296
rect	258	296	259	297
rect	258	297	259	298
rect	258	298	259	299
rect	258	299	259	300
rect	258	300	259	301
rect	258	301	259	302
rect	258	302	259	303
rect	258	303	259	304
rect	258	304	259	305
rect	258	305	259	306
rect	258	306	259	307
rect	258	307	259	308
rect	258	308	259	309
rect	258	309	259	310
rect	258	310	259	311
rect	258	311	259	312
rect	258	312	259	313
rect	258	313	259	314
rect	258	314	259	315
rect	258	315	259	316
rect	258	316	259	317
rect	258	317	259	318
rect	258	318	259	319
rect	258	319	259	320
rect	258	320	259	321
rect	258	321	259	322
rect	258	322	259	323
rect	258	323	259	324
rect	258	324	259	325
rect	258	325	259	326
rect	258	326	259	327
rect	258	327	259	328
rect	258	328	259	329
rect	258	329	259	330
rect	258	330	259	331
rect	258	331	259	332
rect	258	332	259	333
rect	258	333	259	334
rect	258	334	259	335
rect	258	335	259	336
rect	258	336	259	337
rect	258	337	259	338
rect	258	338	259	339
rect	258	339	259	340
rect	258	340	259	341
rect	258	341	259	342
rect	258	342	259	343
rect	258	343	259	344
rect	258	344	259	345
rect	258	345	259	346
rect	258	346	259	347
rect	258	347	259	348
rect	258	348	259	349
rect	258	349	259	350
rect	258	350	259	351
rect	258	351	259	352
rect	258	352	259	353
rect	258	353	259	354
rect	258	354	259	355
rect	258	355	259	356
rect	258	356	259	357
rect	258	357	259	358
rect	258	358	259	359
rect	258	359	259	360
rect	258	360	259	361
rect	258	361	259	362
rect	258	362	259	363
rect	258	363	259	364
rect	258	364	259	365
rect	258	365	259	366
rect	294	0	295	1
rect	294	1	295	2
rect	294	2	295	3
rect	294	3	295	4
rect	294	4	295	5
rect	294	5	295	6
rect	294	6	295	7
rect	294	7	295	8
rect	294	8	295	9
rect	294	9	295	10
rect	294	10	295	11
rect	294	11	295	12
rect	294	12	295	13
rect	294	13	295	14
rect	294	14	295	15
rect	294	15	295	16
rect	294	16	295	17
rect	294	17	295	18
rect	294	18	295	19
rect	294	19	295	20
rect	294	20	295	21
rect	294	21	295	22
rect	294	22	295	23
rect	294	23	295	24
rect	294	24	295	25
rect	294	25	295	26
rect	294	26	295	27
rect	294	27	295	28
rect	294	28	295	29
rect	294	29	295	30
rect	294	30	295	31
rect	294	31	295	32
rect	294	32	295	33
rect	294	33	295	34
rect	294	34	295	35
rect	294	35	295	36
rect	294	36	295	37
rect	294	37	295	38
rect	294	38	295	39
rect	294	39	295	40
rect	294	40	295	41
rect	294	41	295	42
rect	294	42	295	43
rect	294	43	295	44
rect	294	44	295	45
rect	294	45	295	46
rect	294	46	295	47
rect	294	47	295	48
rect	294	48	295	49
rect	294	49	295	50
rect	294	50	295	51
rect	294	51	295	52
rect	294	52	295	53
rect	294	53	295	54
rect	294	54	295	55
rect	294	55	295	56
rect	294	56	295	57
rect	294	57	295	58
rect	294	58	295	59
rect	294	59	295	60
rect	294	60	295	61
rect	294	61	295	62
rect	294	62	295	63
rect	294	63	295	64
rect	294	64	295	65
rect	294	65	295	66
rect	294	66	295	67
rect	294	67	295	68
rect	294	68	295	69
rect	294	69	295	70
rect	294	70	295	71
rect	294	71	295	72
rect	294	72	295	73
rect	294	73	295	74
rect	294	74	295	75
rect	294	75	295	76
rect	294	76	295	77
rect	294	77	295	78
rect	294	78	295	79
rect	294	79	295	80
rect	294	80	295	81
rect	294	81	295	82
rect	294	82	295	83
rect	294	83	295	84
rect	294	84	295	85
rect	294	85	295	86
rect	294	86	295	87
rect	294	87	295	88
rect	294	88	295	89
rect	294	89	295	90
rect	294	90	295	91
rect	294	91	295	92
rect	294	92	295	93
rect	294	93	295	94
rect	294	94	295	95
rect	294	95	295	96
rect	294	96	295	97
rect	294	97	295	98
rect	294	98	295	99
rect	294	99	295	100
rect	294	100	295	101
rect	294	101	295	102
rect	294	102	295	103
rect	294	103	295	104
rect	294	104	295	105
rect	294	105	295	106
rect	294	106	295	107
rect	294	107	295	108
rect	294	108	295	109
rect	294	109	295	110
rect	294	110	295	111
rect	294	111	295	112
rect	294	112	295	113
rect	294	113	295	114
rect	294	114	295	115
rect	294	115	295	116
rect	294	116	295	117
rect	294	117	295	118
rect	294	118	295	119
rect	294	119	295	120
rect	294	120	295	121
rect	294	121	295	122
rect	294	122	295	123
rect	294	123	295	124
rect	294	124	295	125
rect	294	125	295	126
rect	294	126	295	127
rect	294	127	295	128
rect	294	128	295	129
rect	294	129	295	130
rect	294	130	295	131
rect	294	131	295	132
rect	294	132	295	133
rect	294	133	295	134
rect	294	134	295	135
rect	294	135	295	136
rect	294	136	295	137
rect	294	137	295	138
rect	294	138	295	139
rect	294	139	295	140
rect	294	140	295	141
rect	294	141	295	142
rect	294	142	295	143
rect	294	143	295	144
rect	294	144	295	145
rect	294	145	295	146
rect	294	146	295	147
rect	294	147	295	148
rect	294	148	295	149
rect	294	149	295	150
rect	294	150	295	151
rect	294	151	295	152
rect	294	152	295	153
rect	294	153	295	154
rect	294	154	295	155
rect	294	155	295	156
rect	294	156	295	157
rect	294	157	295	158
rect	294	158	295	159
rect	294	159	295	160
rect	294	160	295	161
rect	294	161	295	162
rect	294	162	295	163
rect	294	163	295	164
rect	294	164	295	165
rect	294	165	295	166
rect	294	166	295	167
rect	294	167	295	168
rect	294	168	295	169
rect	294	169	295	170
rect	294	170	295	171
rect	294	171	295	172
rect	294	172	295	173
rect	294	173	295	174
rect	294	174	295	175
rect	294	175	295	176
rect	294	176	295	177
rect	294	177	295	178
rect	294	178	295	179
rect	294	179	295	180
rect	294	180	295	181
rect	294	181	295	182
rect	294	182	295	183
rect	294	183	295	184
rect	294	184	295	185
rect	294	185	295	186
rect	294	186	295	187
rect	294	187	295	188
rect	294	188	295	189
rect	294	189	295	190
rect	294	190	295	191
rect	294	191	295	192
rect	294	192	295	193
rect	294	193	295	194
rect	294	194	295	195
rect	294	195	295	196
rect	294	196	295	197
rect	294	197	295	198
rect	294	198	295	199
rect	294	199	295	200
rect	294	200	295	201
rect	294	201	295	202
rect	294	202	295	203
rect	294	203	295	204
rect	294	204	295	205
rect	294	205	295	206
rect	294	206	295	207
rect	294	207	295	208
rect	294	208	295	209
rect	294	209	295	210
rect	294	210	295	211
rect	294	211	295	212
rect	294	212	295	213
rect	294	213	295	214
rect	294	214	295	215
rect	294	215	295	216
rect	294	216	295	217
rect	294	217	295	218
rect	294	218	295	219
rect	294	219	295	220
rect	294	220	295	221
rect	294	221	295	222
rect	294	222	295	223
rect	294	223	295	224
rect	294	224	295	225
rect	294	225	295	226
rect	294	226	295	227
rect	294	227	295	228
rect	294	228	295	229
rect	294	229	295	230
rect	294	230	295	231
rect	294	231	295	232
rect	294	232	295	233
rect	294	233	295	234
rect	294	234	295	235
rect	294	235	295	236
rect	294	236	295	237
rect	294	237	295	238
rect	294	238	295	239
rect	294	239	295	240
rect	294	240	295	241
rect	294	241	295	242
rect	294	242	295	243
rect	294	243	295	244
rect	294	244	295	245
rect	294	245	295	246
rect	294	246	295	247
rect	294	247	295	248
rect	294	248	295	249
rect	294	249	295	250
rect	294	250	295	251
rect	294	251	295	252
rect	294	252	295	253
rect	294	253	295	254
rect	294	254	295	255
rect	294	255	295	256
rect	294	256	295	257
rect	294	257	295	258
rect	294	258	295	259
rect	294	259	295	260
rect	294	260	295	261
rect	294	261	295	262
rect	294	262	295	263
rect	294	263	295	264
rect	294	264	295	265
rect	294	265	295	266
rect	294	266	295	267
rect	294	267	295	268
rect	294	268	295	269
rect	294	269	295	270
rect	294	270	295	271
rect	294	271	295	272
rect	294	272	295	273
rect	294	273	295	274
rect	294	274	295	275
rect	294	275	295	276
rect	294	276	295	277
rect	294	277	295	278
rect	294	278	295	279
rect	294	279	295	280
rect	294	280	295	281
rect	294	281	295	282
rect	294	282	295	283
rect	294	283	295	284
rect	294	284	295	285
rect	294	285	295	286
rect	294	286	295	287
rect	294	287	295	288
rect	294	288	295	289
rect	294	289	295	290
rect	294	290	295	291
rect	294	291	295	292
rect	294	292	295	293
rect	294	293	295	294
rect	294	294	295	295
rect	294	295	295	296
rect	294	296	295	297
rect	294	297	295	298
rect	294	298	295	299
rect	294	299	295	300
rect	294	300	295	301
rect	294	301	295	302
rect	294	302	295	303
rect	294	303	295	304
rect	294	304	295	305
rect	294	305	295	306
rect	294	306	295	307
rect	294	307	295	308
rect	294	308	295	309
rect	294	309	295	310
rect	294	310	295	311
rect	294	311	295	312
rect	294	312	295	313
rect	294	313	295	314
rect	294	314	295	315
rect	294	315	295	316
rect	294	316	295	317
rect	294	317	295	318
rect	294	318	295	319
rect	294	319	295	320
rect	294	320	295	321
rect	294	321	295	322
rect	294	322	295	323
rect	294	323	295	324
rect	294	324	295	325
rect	294	325	295	326
rect	294	326	295	327
rect	294	327	295	328
rect	294	328	295	329
rect	294	329	295	330
rect	294	330	295	331
rect	294	331	295	332
rect	294	332	295	333
rect	294	333	295	334
rect	294	334	295	335
rect	294	335	295	336
rect	294	336	295	337
rect	294	337	295	338
rect	294	338	295	339
rect	294	339	295	340
rect	294	340	295	341
rect	294	341	295	342
rect	294	342	295	343
rect	294	343	295	344
rect	294	344	295	345
rect	294	345	295	346
rect	294	346	295	347
rect	294	347	295	348
rect	294	348	295	349
rect	294	349	295	350
rect	294	350	295	351
rect	294	351	295	352
rect	294	352	295	353
rect	294	353	295	354
rect	294	354	295	355
rect	294	355	295	356
rect	294	356	295	357
rect	294	357	295	358
rect	294	358	295	359
rect	294	359	295	360
rect	294	360	295	361
rect	294	361	295	362
rect	294	362	295	363
rect	294	363	295	364
rect	294	364	295	365
rect	294	365	295	366
rect	295	0	296	1
rect	295	1	296	2
rect	295	2	296	3
rect	295	3	296	4
rect	295	4	296	5
rect	295	5	296	6
rect	295	6	296	7
rect	295	7	296	8
rect	295	8	296	9
rect	295	9	296	10
rect	295	10	296	11
rect	295	11	296	12
rect	295	12	296	13
rect	295	13	296	14
rect	295	14	296	15
rect	295	15	296	16
rect	295	16	296	17
rect	295	17	296	18
rect	295	18	296	19
rect	295	19	296	20
rect	295	20	296	21
rect	295	21	296	22
rect	295	22	296	23
rect	295	23	296	24
rect	295	24	296	25
rect	295	25	296	26
rect	295	26	296	27
rect	295	27	296	28
rect	295	28	296	29
rect	295	29	296	30
rect	295	30	296	31
rect	295	31	296	32
rect	295	32	296	33
rect	295	33	296	34
rect	295	34	296	35
rect	295	35	296	36
rect	295	36	296	37
rect	295	37	296	38
rect	295	38	296	39
rect	295	39	296	40
rect	295	40	296	41
rect	295	41	296	42
rect	295	42	296	43
rect	295	43	296	44
rect	295	44	296	45
rect	295	45	296	46
rect	295	46	296	47
rect	295	47	296	48
rect	295	48	296	49
rect	295	49	296	50
rect	295	50	296	51
rect	295	51	296	52
rect	295	52	296	53
rect	295	53	296	54
rect	295	54	296	55
rect	295	55	296	56
rect	295	56	296	57
rect	295	57	296	58
rect	295	58	296	59
rect	295	59	296	60
rect	295	60	296	61
rect	295	61	296	62
rect	295	62	296	63
rect	295	63	296	64
rect	295	64	296	65
rect	295	65	296	66
rect	295	66	296	67
rect	295	67	296	68
rect	295	68	296	69
rect	295	69	296	70
rect	295	70	296	71
rect	295	71	296	72
rect	295	72	296	73
rect	295	73	296	74
rect	295	74	296	75
rect	295	75	296	76
rect	295	76	296	77
rect	295	77	296	78
rect	295	78	296	79
rect	295	79	296	80
rect	295	80	296	81
rect	295	81	296	82
rect	295	82	296	83
rect	295	83	296	84
rect	295	84	296	85
rect	295	85	296	86
rect	295	86	296	87
rect	295	87	296	88
rect	295	88	296	89
rect	295	89	296	90
rect	295	90	296	91
rect	295	91	296	92
rect	295	92	296	93
rect	295	93	296	94
rect	295	94	296	95
rect	295	95	296	96
rect	295	96	296	97
rect	295	97	296	98
rect	295	98	296	99
rect	295	99	296	100
rect	295	100	296	101
rect	295	101	296	102
rect	295	102	296	103
rect	295	103	296	104
rect	295	104	296	105
rect	295	105	296	106
rect	295	106	296	107
rect	295	107	296	108
rect	295	108	296	109
rect	295	109	296	110
rect	295	110	296	111
rect	295	111	296	112
rect	295	112	296	113
rect	295	113	296	114
rect	295	114	296	115
rect	295	115	296	116
rect	295	116	296	117
rect	295	117	296	118
rect	295	118	296	119
rect	295	119	296	120
rect	295	120	296	121
rect	295	121	296	122
rect	295	122	296	123
rect	295	123	296	124
rect	295	124	296	125
rect	295	125	296	126
rect	295	126	296	127
rect	295	127	296	128
rect	295	128	296	129
rect	295	129	296	130
rect	295	130	296	131
rect	295	131	296	132
rect	295	132	296	133
rect	295	133	296	134
rect	295	134	296	135
rect	295	135	296	136
rect	295	136	296	137
rect	295	137	296	138
rect	295	138	296	139
rect	295	139	296	140
rect	295	140	296	141
rect	295	141	296	142
rect	295	142	296	143
rect	295	143	296	144
rect	295	144	296	145
rect	295	145	296	146
rect	295	146	296	147
rect	295	147	296	148
rect	295	148	296	149
rect	295	149	296	150
rect	295	150	296	151
rect	295	151	296	152
rect	295	152	296	153
rect	295	153	296	154
rect	295	154	296	155
rect	295	155	296	156
rect	295	156	296	157
rect	295	157	296	158
rect	295	158	296	159
rect	295	159	296	160
rect	295	160	296	161
rect	295	161	296	162
rect	295	162	296	163
rect	295	163	296	164
rect	295	164	296	165
rect	295	165	296	166
rect	295	166	296	167
rect	295	167	296	168
rect	295	168	296	169
rect	295	169	296	170
rect	295	170	296	171
rect	295	171	296	172
rect	295	172	296	173
rect	295	173	296	174
rect	295	174	296	175
rect	295	175	296	176
rect	295	176	296	177
rect	295	177	296	178
rect	295	178	296	179
rect	295	179	296	180
rect	295	180	296	181
rect	295	181	296	182
rect	295	182	296	183
rect	295	183	296	184
rect	295	184	296	185
rect	295	185	296	186
rect	295	186	296	187
rect	295	187	296	188
rect	295	188	296	189
rect	295	189	296	190
rect	295	190	296	191
rect	295	191	296	192
rect	295	192	296	193
rect	295	193	296	194
rect	295	194	296	195
rect	295	195	296	196
rect	295	196	296	197
rect	295	197	296	198
rect	295	198	296	199
rect	295	199	296	200
rect	295	200	296	201
rect	295	201	296	202
rect	295	202	296	203
rect	295	203	296	204
rect	295	204	296	205
rect	295	205	296	206
rect	295	206	296	207
rect	295	207	296	208
rect	295	208	296	209
rect	295	209	296	210
rect	295	210	296	211
rect	295	211	296	212
rect	295	212	296	213
rect	295	213	296	214
rect	295	214	296	215
rect	295	215	296	216
rect	295	216	296	217
rect	295	217	296	218
rect	295	218	296	219
rect	295	219	296	220
rect	295	220	296	221
rect	295	221	296	222
rect	295	222	296	223
rect	295	223	296	224
rect	295	224	296	225
rect	295	225	296	226
rect	295	226	296	227
rect	295	227	296	228
rect	295	228	296	229
rect	295	229	296	230
rect	295	230	296	231
rect	295	231	296	232
rect	295	232	296	233
rect	295	233	296	234
rect	295	234	296	235
rect	295	235	296	236
rect	295	236	296	237
rect	295	237	296	238
rect	295	238	296	239
rect	295	239	296	240
rect	295	240	296	241
rect	295	241	296	242
rect	295	242	296	243
rect	295	243	296	244
rect	295	244	296	245
rect	295	245	296	246
rect	295	246	296	247
rect	295	247	296	248
rect	295	248	296	249
rect	295	249	296	250
rect	295	250	296	251
rect	295	251	296	252
rect	295	252	296	253
rect	295	253	296	254
rect	295	254	296	255
rect	295	255	296	256
rect	295	256	296	257
rect	295	257	296	258
rect	295	258	296	259
rect	295	259	296	260
rect	295	260	296	261
rect	295	261	296	262
rect	295	262	296	263
rect	295	263	296	264
rect	295	264	296	265
rect	295	265	296	266
rect	295	266	296	267
rect	295	267	296	268
rect	295	268	296	269
rect	295	269	296	270
rect	295	270	296	271
rect	295	271	296	272
rect	295	272	296	273
rect	295	273	296	274
rect	295	274	296	275
rect	295	275	296	276
rect	295	276	296	277
rect	295	277	296	278
rect	295	278	296	279
rect	295	279	296	280
rect	295	280	296	281
rect	295	281	296	282
rect	295	282	296	283
rect	295	283	296	284
rect	295	284	296	285
rect	295	285	296	286
rect	295	286	296	287
rect	295	287	296	288
rect	295	288	296	289
rect	295	289	296	290
rect	295	290	296	291
rect	295	291	296	292
rect	295	292	296	293
rect	295	293	296	294
rect	295	294	296	295
rect	295	295	296	296
rect	295	296	296	297
rect	295	297	296	298
rect	295	298	296	299
rect	295	299	296	300
rect	295	300	296	301
rect	295	301	296	302
rect	295	302	296	303
rect	295	303	296	304
rect	295	304	296	305
rect	295	305	296	306
rect	295	306	296	307
rect	295	307	296	308
rect	295	308	296	309
rect	295	309	296	310
rect	295	310	296	311
rect	295	311	296	312
rect	295	312	296	313
rect	295	313	296	314
rect	295	314	296	315
rect	295	315	296	316
rect	295	316	296	317
rect	295	317	296	318
rect	295	318	296	319
rect	295	319	296	320
rect	295	320	296	321
rect	295	321	296	322
rect	295	322	296	323
rect	295	323	296	324
rect	295	324	296	325
rect	295	325	296	326
rect	295	326	296	327
rect	295	327	296	328
rect	295	328	296	329
rect	295	329	296	330
rect	295	330	296	331
rect	295	331	296	332
rect	295	332	296	333
rect	295	333	296	334
rect	295	334	296	335
rect	295	335	296	336
rect	295	336	296	337
rect	295	337	296	338
rect	295	338	296	339
rect	295	339	296	340
rect	295	340	296	341
rect	295	341	296	342
rect	295	342	296	343
rect	295	343	296	344
rect	295	344	296	345
rect	295	345	296	346
rect	295	346	296	347
rect	295	347	296	348
rect	295	348	296	349
rect	295	349	296	350
rect	295	350	296	351
rect	295	351	296	352
rect	295	352	296	353
rect	295	353	296	354
rect	295	354	296	355
rect	295	355	296	356
rect	295	356	296	357
rect	295	357	296	358
rect	295	358	296	359
rect	295	359	296	360
rect	295	360	296	361
rect	295	361	296	362
rect	295	362	296	363
rect	295	363	296	364
rect	295	364	296	365
rect	295	365	296	366
rect	296	0	297	1
rect	296	1	297	2
rect	296	2	297	3
rect	296	3	297	4
rect	296	4	297	5
rect	296	5	297	6
rect	296	6	297	7
rect	296	7	297	8
rect	296	8	297	9
rect	296	9	297	10
rect	296	10	297	11
rect	296	11	297	12
rect	296	12	297	13
rect	296	13	297	14
rect	296	14	297	15
rect	296	15	297	16
rect	296	16	297	17
rect	296	17	297	18
rect	296	18	297	19
rect	296	19	297	20
rect	296	20	297	21
rect	296	21	297	22
rect	296	22	297	23
rect	296	23	297	24
rect	296	24	297	25
rect	296	25	297	26
rect	296	26	297	27
rect	296	27	297	28
rect	296	28	297	29
rect	296	29	297	30
rect	296	30	297	31
rect	296	31	297	32
rect	296	32	297	33
rect	296	33	297	34
rect	296	34	297	35
rect	296	35	297	36
rect	296	36	297	37
rect	296	37	297	38
rect	296	38	297	39
rect	296	39	297	40
rect	296	40	297	41
rect	296	41	297	42
rect	296	42	297	43
rect	296	43	297	44
rect	296	44	297	45
rect	296	45	297	46
rect	296	46	297	47
rect	296	47	297	48
rect	296	48	297	49
rect	296	49	297	50
rect	296	50	297	51
rect	296	51	297	52
rect	296	52	297	53
rect	296	53	297	54
rect	296	54	297	55
rect	296	55	297	56
rect	296	56	297	57
rect	296	57	297	58
rect	296	58	297	59
rect	296	59	297	60
rect	296	60	297	61
rect	296	61	297	62
rect	296	62	297	63
rect	296	63	297	64
rect	296	64	297	65
rect	296	65	297	66
rect	296	66	297	67
rect	296	67	297	68
rect	296	68	297	69
rect	296	69	297	70
rect	296	70	297	71
rect	296	71	297	72
rect	296	72	297	73
rect	296	73	297	74
rect	296	74	297	75
rect	296	75	297	76
rect	296	76	297	77
rect	296	77	297	78
rect	296	78	297	79
rect	296	79	297	80
rect	296	80	297	81
rect	296	81	297	82
rect	296	82	297	83
rect	296	83	297	84
rect	296	84	297	85
rect	296	85	297	86
rect	296	86	297	87
rect	296	87	297	88
rect	296	88	297	89
rect	296	89	297	90
rect	296	90	297	91
rect	296	91	297	92
rect	296	92	297	93
rect	296	93	297	94
rect	296	94	297	95
rect	296	95	297	96
rect	296	96	297	97
rect	296	97	297	98
rect	296	98	297	99
rect	296	99	297	100
rect	296	100	297	101
rect	296	101	297	102
rect	296	102	297	103
rect	296	103	297	104
rect	296	104	297	105
rect	296	105	297	106
rect	296	106	297	107
rect	296	107	297	108
rect	296	108	297	109
rect	296	109	297	110
rect	296	110	297	111
rect	296	111	297	112
rect	296	112	297	113
rect	296	113	297	114
rect	296	114	297	115
rect	296	115	297	116
rect	296	116	297	117
rect	296	117	297	118
rect	296	118	297	119
rect	296	119	297	120
rect	296	120	297	121
rect	296	121	297	122
rect	296	122	297	123
rect	296	123	297	124
rect	296	124	297	125
rect	296	125	297	126
rect	296	126	297	127
rect	296	127	297	128
rect	296	128	297	129
rect	296	129	297	130
rect	296	130	297	131
rect	296	131	297	132
rect	296	132	297	133
rect	296	133	297	134
rect	296	134	297	135
rect	296	135	297	136
rect	296	136	297	137
rect	296	137	297	138
rect	296	138	297	139
rect	296	139	297	140
rect	296	140	297	141
rect	296	141	297	142
rect	296	142	297	143
rect	296	143	297	144
rect	296	144	297	145
rect	296	145	297	146
rect	296	146	297	147
rect	296	147	297	148
rect	296	148	297	149
rect	296	149	297	150
rect	296	150	297	151
rect	296	151	297	152
rect	296	152	297	153
rect	296	153	297	154
rect	296	154	297	155
rect	296	155	297	156
rect	296	156	297	157
rect	296	157	297	158
rect	296	158	297	159
rect	296	159	297	160
rect	296	160	297	161
rect	296	161	297	162
rect	296	162	297	163
rect	296	163	297	164
rect	296	164	297	165
rect	296	165	297	166
rect	296	166	297	167
rect	296	167	297	168
rect	296	168	297	169
rect	296	169	297	170
rect	296	170	297	171
rect	296	171	297	172
rect	296	172	297	173
rect	296	173	297	174
rect	296	174	297	175
rect	296	175	297	176
rect	296	176	297	177
rect	296	177	297	178
rect	296	178	297	179
rect	296	179	297	180
rect	296	180	297	181
rect	296	181	297	182
rect	296	182	297	183
rect	296	183	297	184
rect	296	184	297	185
rect	296	185	297	186
rect	296	186	297	187
rect	296	187	297	188
rect	296	188	297	189
rect	296	189	297	190
rect	296	190	297	191
rect	296	191	297	192
rect	296	192	297	193
rect	296	193	297	194
rect	296	194	297	195
rect	296	195	297	196
rect	296	196	297	197
rect	296	197	297	198
rect	296	198	297	199
rect	296	199	297	200
rect	296	200	297	201
rect	296	201	297	202
rect	296	202	297	203
rect	296	203	297	204
rect	296	204	297	205
rect	296	205	297	206
rect	296	206	297	207
rect	296	207	297	208
rect	296	208	297	209
rect	296	209	297	210
rect	296	210	297	211
rect	296	211	297	212
rect	296	212	297	213
rect	296	213	297	214
rect	296	214	297	215
rect	296	215	297	216
rect	296	216	297	217
rect	296	217	297	218
rect	296	218	297	219
rect	296	219	297	220
rect	296	220	297	221
rect	296	221	297	222
rect	296	222	297	223
rect	296	223	297	224
rect	296	224	297	225
rect	296	225	297	226
rect	296	226	297	227
rect	296	227	297	228
rect	296	228	297	229
rect	296	229	297	230
rect	296	230	297	231
rect	296	231	297	232
rect	296	232	297	233
rect	296	233	297	234
rect	296	234	297	235
rect	296	235	297	236
rect	296	236	297	237
rect	296	237	297	238
rect	296	238	297	239
rect	296	239	297	240
rect	296	240	297	241
rect	296	241	297	242
rect	296	242	297	243
rect	296	243	297	244
rect	296	244	297	245
rect	296	245	297	246
rect	296	246	297	247
rect	296	247	297	248
rect	296	248	297	249
rect	296	249	297	250
rect	296	250	297	251
rect	296	251	297	252
rect	296	252	297	253
rect	296	253	297	254
rect	296	254	297	255
rect	296	255	297	256
rect	296	256	297	257
rect	296	257	297	258
rect	296	258	297	259
rect	296	259	297	260
rect	296	260	297	261
rect	296	261	297	262
rect	296	262	297	263
rect	296	263	297	264
rect	296	264	297	265
rect	296	265	297	266
rect	296	266	297	267
rect	296	267	297	268
rect	296	268	297	269
rect	296	269	297	270
rect	296	270	297	271
rect	296	271	297	272
rect	296	272	297	273
rect	296	273	297	274
rect	296	274	297	275
rect	296	275	297	276
rect	296	276	297	277
rect	296	277	297	278
rect	296	278	297	279
rect	296	279	297	280
rect	296	280	297	281
rect	296	281	297	282
rect	296	282	297	283
rect	296	283	297	284
rect	296	284	297	285
rect	296	285	297	286
rect	296	286	297	287
rect	296	287	297	288
rect	296	288	297	289
rect	296	289	297	290
rect	296	290	297	291
rect	296	291	297	292
rect	296	292	297	293
rect	296	293	297	294
rect	296	294	297	295
rect	296	295	297	296
rect	296	296	297	297
rect	296	297	297	298
rect	296	298	297	299
rect	296	299	297	300
rect	296	300	297	301
rect	296	301	297	302
rect	296	302	297	303
rect	296	303	297	304
rect	296	304	297	305
rect	296	305	297	306
rect	296	306	297	307
rect	296	307	297	308
rect	296	308	297	309
rect	296	309	297	310
rect	296	310	297	311
rect	296	311	297	312
rect	296	312	297	313
rect	296	313	297	314
rect	296	314	297	315
rect	296	315	297	316
rect	296	316	297	317
rect	296	317	297	318
rect	296	318	297	319
rect	296	319	297	320
rect	296	320	297	321
rect	296	321	297	322
rect	296	322	297	323
rect	296	323	297	324
rect	296	324	297	325
rect	296	325	297	326
rect	296	326	297	327
rect	296	327	297	328
rect	296	328	297	329
rect	296	329	297	330
rect	296	330	297	331
rect	296	331	297	332
rect	296	332	297	333
rect	296	333	297	334
rect	296	334	297	335
rect	296	335	297	336
rect	296	336	297	337
rect	296	337	297	338
rect	296	338	297	339
rect	296	339	297	340
rect	296	340	297	341
rect	296	341	297	342
rect	296	342	297	343
rect	296	343	297	344
rect	296	344	297	345
rect	296	345	297	346
rect	296	346	297	347
rect	296	347	297	348
rect	296	348	297	349
rect	296	349	297	350
rect	296	350	297	351
rect	296	351	297	352
rect	296	352	297	353
rect	296	353	297	354
rect	296	354	297	355
rect	296	355	297	356
rect	296	356	297	357
rect	296	357	297	358
rect	296	358	297	359
rect	296	359	297	360
rect	296	360	297	361
rect	296	361	297	362
rect	296	362	297	363
rect	296	363	297	364
rect	296	364	297	365
rect	296	365	297	366
rect	297	0	298	1
rect	297	1	298	2
rect	297	2	298	3
rect	297	3	298	4
rect	297	4	298	5
rect	297	5	298	6
rect	297	6	298	7
rect	297	7	298	8
rect	297	8	298	9
rect	297	9	298	10
rect	297	10	298	11
rect	297	11	298	12
rect	297	12	298	13
rect	297	13	298	14
rect	297	14	298	15
rect	297	15	298	16
rect	297	16	298	17
rect	297	17	298	18
rect	297	18	298	19
rect	297	19	298	20
rect	297	20	298	21
rect	297	21	298	22
rect	297	22	298	23
rect	297	23	298	24
rect	297	24	298	25
rect	297	25	298	26
rect	297	26	298	27
rect	297	27	298	28
rect	297	28	298	29
rect	297	29	298	30
rect	297	30	298	31
rect	297	31	298	32
rect	297	32	298	33
rect	297	33	298	34
rect	297	34	298	35
rect	297	35	298	36
rect	297	36	298	37
rect	297	37	298	38
rect	297	38	298	39
rect	297	39	298	40
rect	297	40	298	41
rect	297	41	298	42
rect	297	42	298	43
rect	297	43	298	44
rect	297	44	298	45
rect	297	45	298	46
rect	297	46	298	47
rect	297	47	298	48
rect	297	48	298	49
rect	297	49	298	50
rect	297	50	298	51
rect	297	51	298	52
rect	297	52	298	53
rect	297	53	298	54
rect	297	54	298	55
rect	297	55	298	56
rect	297	56	298	57
rect	297	57	298	58
rect	297	58	298	59
rect	297	59	298	60
rect	297	60	298	61
rect	297	61	298	62
rect	297	62	298	63
rect	297	63	298	64
rect	297	64	298	65
rect	297	65	298	66
rect	297	66	298	67
rect	297	67	298	68
rect	297	68	298	69
rect	297	69	298	70
rect	297	70	298	71
rect	297	71	298	72
rect	297	72	298	73
rect	297	73	298	74
rect	297	74	298	75
rect	297	75	298	76
rect	297	76	298	77
rect	297	77	298	78
rect	297	78	298	79
rect	297	79	298	80
rect	297	80	298	81
rect	297	81	298	82
rect	297	82	298	83
rect	297	83	298	84
rect	297	84	298	85
rect	297	85	298	86
rect	297	86	298	87
rect	297	87	298	88
rect	297	88	298	89
rect	297	89	298	90
rect	297	90	298	91
rect	297	91	298	92
rect	297	92	298	93
rect	297	93	298	94
rect	297	94	298	95
rect	297	95	298	96
rect	297	96	298	97
rect	297	97	298	98
rect	297	98	298	99
rect	297	99	298	100
rect	297	100	298	101
rect	297	101	298	102
rect	297	102	298	103
rect	297	103	298	104
rect	297	104	298	105
rect	297	105	298	106
rect	297	106	298	107
rect	297	107	298	108
rect	297	108	298	109
rect	297	109	298	110
rect	297	110	298	111
rect	297	111	298	112
rect	297	112	298	113
rect	297	113	298	114
rect	297	114	298	115
rect	297	115	298	116
rect	297	116	298	117
rect	297	117	298	118
rect	297	118	298	119
rect	297	119	298	120
rect	297	120	298	121
rect	297	121	298	122
rect	297	122	298	123
rect	297	123	298	124
rect	297	124	298	125
rect	297	125	298	126
rect	297	126	298	127
rect	297	127	298	128
rect	297	128	298	129
rect	297	129	298	130
rect	297	130	298	131
rect	297	131	298	132
rect	297	132	298	133
rect	297	133	298	134
rect	297	134	298	135
rect	297	135	298	136
rect	297	136	298	137
rect	297	137	298	138
rect	297	138	298	139
rect	297	139	298	140
rect	297	140	298	141
rect	297	141	298	142
rect	297	142	298	143
rect	297	143	298	144
rect	297	144	298	145
rect	297	145	298	146
rect	297	146	298	147
rect	297	147	298	148
rect	297	148	298	149
rect	297	149	298	150
rect	297	150	298	151
rect	297	151	298	152
rect	297	152	298	153
rect	297	153	298	154
rect	297	154	298	155
rect	297	155	298	156
rect	297	156	298	157
rect	297	157	298	158
rect	297	158	298	159
rect	297	159	298	160
rect	297	160	298	161
rect	297	161	298	162
rect	297	162	298	163
rect	297	163	298	164
rect	297	164	298	165
rect	297	165	298	166
rect	297	166	298	167
rect	297	167	298	168
rect	297	168	298	169
rect	297	169	298	170
rect	297	170	298	171
rect	297	171	298	172
rect	297	172	298	173
rect	297	173	298	174
rect	297	174	298	175
rect	297	175	298	176
rect	297	176	298	177
rect	297	177	298	178
rect	297	178	298	179
rect	297	179	298	180
rect	297	180	298	181
rect	297	181	298	182
rect	297	182	298	183
rect	297	183	298	184
rect	297	184	298	185
rect	297	185	298	186
rect	297	186	298	187
rect	297	187	298	188
rect	297	188	298	189
rect	297	189	298	190
rect	297	190	298	191
rect	297	191	298	192
rect	297	192	298	193
rect	297	193	298	194
rect	297	194	298	195
rect	297	195	298	196
rect	297	196	298	197
rect	297	197	298	198
rect	297	198	298	199
rect	297	199	298	200
rect	297	200	298	201
rect	297	201	298	202
rect	297	202	298	203
rect	297	203	298	204
rect	297	204	298	205
rect	297	205	298	206
rect	297	206	298	207
rect	297	207	298	208
rect	297	208	298	209
rect	297	209	298	210
rect	297	210	298	211
rect	297	211	298	212
rect	297	212	298	213
rect	297	213	298	214
rect	297	214	298	215
rect	297	215	298	216
rect	297	216	298	217
rect	297	217	298	218
rect	297	218	298	219
rect	297	219	298	220
rect	297	220	298	221
rect	297	221	298	222
rect	297	222	298	223
rect	297	223	298	224
rect	297	224	298	225
rect	297	225	298	226
rect	297	226	298	227
rect	297	227	298	228
rect	297	228	298	229
rect	297	229	298	230
rect	297	230	298	231
rect	297	231	298	232
rect	297	232	298	233
rect	297	233	298	234
rect	297	234	298	235
rect	297	235	298	236
rect	297	236	298	237
rect	297	237	298	238
rect	297	238	298	239
rect	297	239	298	240
rect	297	240	298	241
rect	297	241	298	242
rect	297	242	298	243
rect	297	243	298	244
rect	297	244	298	245
rect	297	245	298	246
rect	297	246	298	247
rect	297	247	298	248
rect	297	248	298	249
rect	297	249	298	250
rect	297	250	298	251
rect	297	251	298	252
rect	297	252	298	253
rect	297	253	298	254
rect	297	254	298	255
rect	297	255	298	256
rect	297	256	298	257
rect	297	257	298	258
rect	297	258	298	259
rect	297	259	298	260
rect	297	260	298	261
rect	297	261	298	262
rect	297	262	298	263
rect	297	263	298	264
rect	297	264	298	265
rect	297	265	298	266
rect	297	266	298	267
rect	297	267	298	268
rect	297	268	298	269
rect	297	269	298	270
rect	297	270	298	271
rect	297	271	298	272
rect	297	272	298	273
rect	297	273	298	274
rect	297	274	298	275
rect	297	275	298	276
rect	297	276	298	277
rect	297	277	298	278
rect	297	278	298	279
rect	297	279	298	280
rect	297	280	298	281
rect	297	281	298	282
rect	297	282	298	283
rect	297	283	298	284
rect	297	284	298	285
rect	297	285	298	286
rect	297	286	298	287
rect	297	287	298	288
rect	297	288	298	289
rect	297	289	298	290
rect	297	290	298	291
rect	297	291	298	292
rect	297	292	298	293
rect	297	293	298	294
rect	297	294	298	295
rect	297	295	298	296
rect	297	296	298	297
rect	297	297	298	298
rect	297	298	298	299
rect	297	299	298	300
rect	297	300	298	301
rect	297	301	298	302
rect	297	302	298	303
rect	297	303	298	304
rect	297	304	298	305
rect	297	305	298	306
rect	297	306	298	307
rect	297	307	298	308
rect	297	308	298	309
rect	297	309	298	310
rect	297	310	298	311
rect	297	311	298	312
rect	297	312	298	313
rect	297	313	298	314
rect	297	314	298	315
rect	297	315	298	316
rect	297	316	298	317
rect	297	317	298	318
rect	297	318	298	319
rect	297	319	298	320
rect	297	320	298	321
rect	297	321	298	322
rect	297	322	298	323
rect	297	323	298	324
rect	297	324	298	325
rect	297	325	298	326
rect	297	326	298	327
rect	297	327	298	328
rect	297	328	298	329
rect	297	329	298	330
rect	297	330	298	331
rect	297	331	298	332
rect	297	332	298	333
rect	297	333	298	334
rect	297	334	298	335
rect	297	335	298	336
rect	297	336	298	337
rect	297	337	298	338
rect	297	338	298	339
rect	297	339	298	340
rect	297	340	298	341
rect	297	341	298	342
rect	297	342	298	343
rect	297	343	298	344
rect	297	344	298	345
rect	297	345	298	346
rect	297	346	298	347
rect	297	347	298	348
rect	297	348	298	349
rect	297	349	298	350
rect	297	350	298	351
rect	297	351	298	352
rect	297	352	298	353
rect	297	353	298	354
rect	297	354	298	355
rect	297	355	298	356
rect	297	356	298	357
rect	297	357	298	358
rect	297	358	298	359
rect	297	359	298	360
rect	297	360	298	361
rect	297	361	298	362
rect	297	362	298	363
rect	297	363	298	364
rect	297	364	298	365
rect	297	365	298	366
rect	298	0	299	1
rect	298	1	299	2
rect	298	2	299	3
rect	298	3	299	4
rect	298	4	299	5
rect	298	5	299	6
rect	298	6	299	7
rect	298	7	299	8
rect	298	8	299	9
rect	298	9	299	10
rect	298	10	299	11
rect	298	11	299	12
rect	298	12	299	13
rect	298	13	299	14
rect	298	14	299	15
rect	298	15	299	16
rect	298	16	299	17
rect	298	17	299	18
rect	298	18	299	19
rect	298	19	299	20
rect	298	20	299	21
rect	298	21	299	22
rect	298	22	299	23
rect	298	23	299	24
rect	298	24	299	25
rect	298	25	299	26
rect	298	26	299	27
rect	298	27	299	28
rect	298	28	299	29
rect	298	29	299	30
rect	298	30	299	31
rect	298	31	299	32
rect	298	32	299	33
rect	298	33	299	34
rect	298	34	299	35
rect	298	35	299	36
rect	298	36	299	37
rect	298	37	299	38
rect	298	38	299	39
rect	298	39	299	40
rect	298	40	299	41
rect	298	41	299	42
rect	298	42	299	43
rect	298	43	299	44
rect	298	44	299	45
rect	298	45	299	46
rect	298	46	299	47
rect	298	47	299	48
rect	298	48	299	49
rect	298	49	299	50
rect	298	50	299	51
rect	298	51	299	52
rect	298	52	299	53
rect	298	53	299	54
rect	298	54	299	55
rect	298	55	299	56
rect	298	56	299	57
rect	298	57	299	58
rect	298	58	299	59
rect	298	59	299	60
rect	298	60	299	61
rect	298	61	299	62
rect	298	62	299	63
rect	298	63	299	64
rect	298	64	299	65
rect	298	65	299	66
rect	298	66	299	67
rect	298	67	299	68
rect	298	68	299	69
rect	298	69	299	70
rect	298	70	299	71
rect	298	71	299	72
rect	298	72	299	73
rect	298	73	299	74
rect	298	74	299	75
rect	298	75	299	76
rect	298	76	299	77
rect	298	77	299	78
rect	298	78	299	79
rect	298	79	299	80
rect	298	80	299	81
rect	298	81	299	82
rect	298	82	299	83
rect	298	83	299	84
rect	298	84	299	85
rect	298	85	299	86
rect	298	86	299	87
rect	298	87	299	88
rect	298	88	299	89
rect	298	89	299	90
rect	298	90	299	91
rect	298	91	299	92
rect	298	92	299	93
rect	298	93	299	94
rect	298	94	299	95
rect	298	95	299	96
rect	298	96	299	97
rect	298	97	299	98
rect	298	98	299	99
rect	298	99	299	100
rect	298	100	299	101
rect	298	101	299	102
rect	298	102	299	103
rect	298	103	299	104
rect	298	104	299	105
rect	298	105	299	106
rect	298	106	299	107
rect	298	107	299	108
rect	298	108	299	109
rect	298	109	299	110
rect	298	110	299	111
rect	298	111	299	112
rect	298	112	299	113
rect	298	113	299	114
rect	298	114	299	115
rect	298	115	299	116
rect	298	116	299	117
rect	298	117	299	118
rect	298	118	299	119
rect	298	119	299	120
rect	298	120	299	121
rect	298	121	299	122
rect	298	122	299	123
rect	298	123	299	124
rect	298	124	299	125
rect	298	125	299	126
rect	298	126	299	127
rect	298	127	299	128
rect	298	128	299	129
rect	298	129	299	130
rect	298	130	299	131
rect	298	131	299	132
rect	298	132	299	133
rect	298	133	299	134
rect	298	134	299	135
rect	298	135	299	136
rect	298	136	299	137
rect	298	137	299	138
rect	298	138	299	139
rect	298	139	299	140
rect	298	140	299	141
rect	298	141	299	142
rect	298	142	299	143
rect	298	143	299	144
rect	298	144	299	145
rect	298	145	299	146
rect	298	146	299	147
rect	298	147	299	148
rect	298	148	299	149
rect	298	149	299	150
rect	298	150	299	151
rect	298	151	299	152
rect	298	152	299	153
rect	298	153	299	154
rect	298	154	299	155
rect	298	155	299	156
rect	298	156	299	157
rect	298	157	299	158
rect	298	158	299	159
rect	298	159	299	160
rect	298	160	299	161
rect	298	161	299	162
rect	298	162	299	163
rect	298	163	299	164
rect	298	164	299	165
rect	298	165	299	166
rect	298	166	299	167
rect	298	167	299	168
rect	298	168	299	169
rect	298	169	299	170
rect	298	170	299	171
rect	298	171	299	172
rect	298	172	299	173
rect	298	173	299	174
rect	298	174	299	175
rect	298	175	299	176
rect	298	176	299	177
rect	298	177	299	178
rect	298	178	299	179
rect	298	179	299	180
rect	298	180	299	181
rect	298	181	299	182
rect	298	182	299	183
rect	298	183	299	184
rect	298	184	299	185
rect	298	185	299	186
rect	298	186	299	187
rect	298	187	299	188
rect	298	188	299	189
rect	298	189	299	190
rect	298	190	299	191
rect	298	191	299	192
rect	298	192	299	193
rect	298	193	299	194
rect	298	194	299	195
rect	298	195	299	196
rect	298	196	299	197
rect	298	197	299	198
rect	298	198	299	199
rect	298	199	299	200
rect	298	200	299	201
rect	298	201	299	202
rect	298	202	299	203
rect	298	203	299	204
rect	298	204	299	205
rect	298	205	299	206
rect	298	206	299	207
rect	298	207	299	208
rect	298	208	299	209
rect	298	209	299	210
rect	298	210	299	211
rect	298	211	299	212
rect	298	212	299	213
rect	298	213	299	214
rect	298	214	299	215
rect	298	215	299	216
rect	298	216	299	217
rect	298	217	299	218
rect	298	218	299	219
rect	298	219	299	220
rect	298	220	299	221
rect	298	221	299	222
rect	298	222	299	223
rect	298	223	299	224
rect	298	224	299	225
rect	298	225	299	226
rect	298	226	299	227
rect	298	227	299	228
rect	298	228	299	229
rect	298	229	299	230
rect	298	230	299	231
rect	298	231	299	232
rect	298	232	299	233
rect	298	233	299	234
rect	298	234	299	235
rect	298	235	299	236
rect	298	236	299	237
rect	298	237	299	238
rect	298	238	299	239
rect	298	239	299	240
rect	298	240	299	241
rect	298	241	299	242
rect	298	242	299	243
rect	298	243	299	244
rect	298	244	299	245
rect	298	245	299	246
rect	298	246	299	247
rect	298	247	299	248
rect	298	248	299	249
rect	298	249	299	250
rect	298	250	299	251
rect	298	251	299	252
rect	298	252	299	253
rect	298	253	299	254
rect	298	254	299	255
rect	298	255	299	256
rect	298	256	299	257
rect	298	257	299	258
rect	298	258	299	259
rect	298	259	299	260
rect	298	260	299	261
rect	298	261	299	262
rect	298	262	299	263
rect	298	263	299	264
rect	298	264	299	265
rect	298	265	299	266
rect	298	266	299	267
rect	298	267	299	268
rect	298	268	299	269
rect	298	269	299	270
rect	298	270	299	271
rect	298	271	299	272
rect	298	272	299	273
rect	298	273	299	274
rect	298	274	299	275
rect	298	275	299	276
rect	298	276	299	277
rect	298	277	299	278
rect	298	278	299	279
rect	298	279	299	280
rect	298	280	299	281
rect	298	281	299	282
rect	298	282	299	283
rect	298	283	299	284
rect	298	284	299	285
rect	298	285	299	286
rect	298	286	299	287
rect	298	287	299	288
rect	298	288	299	289
rect	298	289	299	290
rect	298	290	299	291
rect	298	291	299	292
rect	298	292	299	293
rect	298	293	299	294
rect	298	294	299	295
rect	298	295	299	296
rect	298	296	299	297
rect	298	297	299	298
rect	298	298	299	299
rect	298	299	299	300
rect	298	300	299	301
rect	298	301	299	302
rect	298	302	299	303
rect	298	303	299	304
rect	298	304	299	305
rect	298	305	299	306
rect	298	306	299	307
rect	298	307	299	308
rect	298	308	299	309
rect	298	309	299	310
rect	298	310	299	311
rect	298	311	299	312
rect	298	312	299	313
rect	298	313	299	314
rect	298	314	299	315
rect	298	315	299	316
rect	298	316	299	317
rect	298	317	299	318
rect	298	318	299	319
rect	298	319	299	320
rect	298	320	299	321
rect	298	321	299	322
rect	298	322	299	323
rect	298	323	299	324
rect	298	324	299	325
rect	298	325	299	326
rect	298	326	299	327
rect	298	327	299	328
rect	298	328	299	329
rect	298	329	299	330
rect	298	330	299	331
rect	298	331	299	332
rect	298	332	299	333
rect	298	333	299	334
rect	298	334	299	335
rect	298	335	299	336
rect	298	336	299	337
rect	298	337	299	338
rect	298	338	299	339
rect	298	339	299	340
rect	298	340	299	341
rect	298	341	299	342
rect	298	342	299	343
rect	298	343	299	344
rect	298	344	299	345
rect	298	345	299	346
rect	298	346	299	347
rect	298	347	299	348
rect	298	348	299	349
rect	298	349	299	350
rect	298	350	299	351
rect	298	351	299	352
rect	298	352	299	353
rect	298	353	299	354
rect	298	354	299	355
rect	298	355	299	356
rect	298	356	299	357
rect	298	357	299	358
rect	298	358	299	359
rect	298	359	299	360
rect	298	360	299	361
rect	298	361	299	362
rect	298	362	299	363
rect	298	363	299	364
rect	298	364	299	365
rect	298	365	299	366
rect	299	0	300	1
rect	299	1	300	2
rect	299	2	300	3
rect	299	3	300	4
rect	299	4	300	5
rect	299	5	300	6
rect	299	6	300	7
rect	299	7	300	8
rect	299	8	300	9
rect	299	9	300	10
rect	299	10	300	11
rect	299	11	300	12
rect	299	12	300	13
rect	299	13	300	14
rect	299	14	300	15
rect	299	15	300	16
rect	299	16	300	17
rect	299	17	300	18
rect	299	18	300	19
rect	299	19	300	20
rect	299	20	300	21
rect	299	21	300	22
rect	299	22	300	23
rect	299	23	300	24
rect	299	24	300	25
rect	299	25	300	26
rect	299	26	300	27
rect	299	27	300	28
rect	299	28	300	29
rect	299	29	300	30
rect	299	30	300	31
rect	299	31	300	32
rect	299	32	300	33
rect	299	33	300	34
rect	299	34	300	35
rect	299	35	300	36
rect	299	36	300	37
rect	299	37	300	38
rect	299	38	300	39
rect	299	39	300	40
rect	299	40	300	41
rect	299	41	300	42
rect	299	42	300	43
rect	299	43	300	44
rect	299	44	300	45
rect	299	45	300	46
rect	299	46	300	47
rect	299	47	300	48
rect	299	48	300	49
rect	299	49	300	50
rect	299	50	300	51
rect	299	51	300	52
rect	299	52	300	53
rect	299	53	300	54
rect	299	54	300	55
rect	299	55	300	56
rect	299	56	300	57
rect	299	57	300	58
rect	299	58	300	59
rect	299	59	300	60
rect	299	60	300	61
rect	299	61	300	62
rect	299	62	300	63
rect	299	63	300	64
rect	299	64	300	65
rect	299	65	300	66
rect	299	66	300	67
rect	299	67	300	68
rect	299	68	300	69
rect	299	69	300	70
rect	299	70	300	71
rect	299	71	300	72
rect	299	72	300	73
rect	299	73	300	74
rect	299	74	300	75
rect	299	75	300	76
rect	299	76	300	77
rect	299	77	300	78
rect	299	78	300	79
rect	299	79	300	80
rect	299	80	300	81
rect	299	81	300	82
rect	299	82	300	83
rect	299	83	300	84
rect	299	84	300	85
rect	299	85	300	86
rect	299	86	300	87
rect	299	87	300	88
rect	299	88	300	89
rect	299	89	300	90
rect	299	90	300	91
rect	299	91	300	92
rect	299	92	300	93
rect	299	93	300	94
rect	299	94	300	95
rect	299	95	300	96
rect	299	96	300	97
rect	299	97	300	98
rect	299	98	300	99
rect	299	99	300	100
rect	299	100	300	101
rect	299	101	300	102
rect	299	102	300	103
rect	299	103	300	104
rect	299	104	300	105
rect	299	105	300	106
rect	299	106	300	107
rect	299	107	300	108
rect	299	108	300	109
rect	299	109	300	110
rect	299	110	300	111
rect	299	111	300	112
rect	299	112	300	113
rect	299	113	300	114
rect	299	114	300	115
rect	299	115	300	116
rect	299	116	300	117
rect	299	117	300	118
rect	299	118	300	119
rect	299	119	300	120
rect	299	120	300	121
rect	299	121	300	122
rect	299	122	300	123
rect	299	123	300	124
rect	299	124	300	125
rect	299	125	300	126
rect	299	126	300	127
rect	299	127	300	128
rect	299	128	300	129
rect	299	129	300	130
rect	299	130	300	131
rect	299	131	300	132
rect	299	132	300	133
rect	299	133	300	134
rect	299	134	300	135
rect	299	135	300	136
rect	299	136	300	137
rect	299	137	300	138
rect	299	138	300	139
rect	299	139	300	140
rect	299	140	300	141
rect	299	141	300	142
rect	299	142	300	143
rect	299	143	300	144
rect	299	144	300	145
rect	299	145	300	146
rect	299	146	300	147
rect	299	147	300	148
rect	299	148	300	149
rect	299	149	300	150
rect	299	150	300	151
rect	299	151	300	152
rect	299	152	300	153
rect	299	153	300	154
rect	299	154	300	155
rect	299	155	300	156
rect	299	156	300	157
rect	299	157	300	158
rect	299	158	300	159
rect	299	159	300	160
rect	299	160	300	161
rect	299	161	300	162
rect	299	162	300	163
rect	299	163	300	164
rect	299	164	300	165
rect	299	165	300	166
rect	299	166	300	167
rect	299	167	300	168
rect	299	168	300	169
rect	299	169	300	170
rect	299	170	300	171
rect	299	171	300	172
rect	299	172	300	173
rect	299	173	300	174
rect	299	174	300	175
rect	299	175	300	176
rect	299	176	300	177
rect	299	177	300	178
rect	299	178	300	179
rect	299	179	300	180
rect	299	180	300	181
rect	299	181	300	182
rect	299	182	300	183
rect	299	183	300	184
rect	299	184	300	185
rect	299	185	300	186
rect	299	186	300	187
rect	299	187	300	188
rect	299	188	300	189
rect	299	189	300	190
rect	299	190	300	191
rect	299	191	300	192
rect	299	192	300	193
rect	299	193	300	194
rect	299	194	300	195
rect	299	195	300	196
rect	299	196	300	197
rect	299	197	300	198
rect	299	198	300	199
rect	299	199	300	200
rect	299	200	300	201
rect	299	201	300	202
rect	299	202	300	203
rect	299	203	300	204
rect	299	204	300	205
rect	299	205	300	206
rect	299	206	300	207
rect	299	207	300	208
rect	299	208	300	209
rect	299	209	300	210
rect	299	210	300	211
rect	299	211	300	212
rect	299	212	300	213
rect	299	213	300	214
rect	299	214	300	215
rect	299	215	300	216
rect	299	216	300	217
rect	299	217	300	218
rect	299	218	300	219
rect	299	219	300	220
rect	299	220	300	221
rect	299	221	300	222
rect	299	222	300	223
rect	299	223	300	224
rect	299	224	300	225
rect	299	225	300	226
rect	299	226	300	227
rect	299	227	300	228
rect	299	228	300	229
rect	299	229	300	230
rect	299	230	300	231
rect	299	231	300	232
rect	299	232	300	233
rect	299	233	300	234
rect	299	234	300	235
rect	299	235	300	236
rect	299	236	300	237
rect	299	237	300	238
rect	299	238	300	239
rect	299	239	300	240
rect	299	240	300	241
rect	299	241	300	242
rect	299	242	300	243
rect	299	243	300	244
rect	299	244	300	245
rect	299	245	300	246
rect	299	246	300	247
rect	299	247	300	248
rect	299	248	300	249
rect	299	249	300	250
rect	299	250	300	251
rect	299	251	300	252
rect	299	252	300	253
rect	299	253	300	254
rect	299	254	300	255
rect	299	255	300	256
rect	299	256	300	257
rect	299	257	300	258
rect	299	258	300	259
rect	299	259	300	260
rect	299	260	300	261
rect	299	261	300	262
rect	299	262	300	263
rect	299	263	300	264
rect	299	264	300	265
rect	299	265	300	266
rect	299	266	300	267
rect	299	267	300	268
rect	299	268	300	269
rect	299	269	300	270
rect	299	270	300	271
rect	299	271	300	272
rect	299	272	300	273
rect	299	273	300	274
rect	299	274	300	275
rect	299	275	300	276
rect	299	276	300	277
rect	299	277	300	278
rect	299	278	300	279
rect	299	279	300	280
rect	299	280	300	281
rect	299	281	300	282
rect	299	282	300	283
rect	299	283	300	284
rect	299	284	300	285
rect	299	285	300	286
rect	299	286	300	287
rect	299	287	300	288
rect	299	288	300	289
rect	299	289	300	290
rect	299	290	300	291
rect	299	291	300	292
rect	299	292	300	293
rect	299	293	300	294
rect	299	294	300	295
rect	299	295	300	296
rect	299	296	300	297
rect	299	297	300	298
rect	299	298	300	299
rect	299	299	300	300
rect	299	300	300	301
rect	299	301	300	302
rect	299	302	300	303
rect	299	303	300	304
rect	299	304	300	305
rect	299	305	300	306
rect	299	306	300	307
rect	299	307	300	308
rect	299	308	300	309
rect	299	309	300	310
rect	299	310	300	311
rect	299	311	300	312
rect	299	312	300	313
rect	299	313	300	314
rect	299	314	300	315
rect	299	315	300	316
rect	299	316	300	317
rect	299	317	300	318
rect	299	318	300	319
rect	299	319	300	320
rect	299	320	300	321
rect	299	321	300	322
rect	299	322	300	323
rect	299	323	300	324
rect	299	324	300	325
rect	299	325	300	326
rect	299	326	300	327
rect	299	327	300	328
rect	299	328	300	329
rect	299	329	300	330
rect	299	330	300	331
rect	299	331	300	332
rect	299	332	300	333
rect	299	333	300	334
rect	299	334	300	335
rect	299	335	300	336
rect	299	336	300	337
rect	299	337	300	338
rect	299	338	300	339
rect	299	339	300	340
rect	299	340	300	341
rect	299	341	300	342
rect	299	342	300	343
rect	299	343	300	344
rect	299	344	300	345
rect	299	345	300	346
rect	299	346	300	347
rect	299	347	300	348
rect	299	348	300	349
rect	299	349	300	350
rect	299	350	300	351
rect	299	351	300	352
rect	299	352	300	353
rect	299	353	300	354
rect	299	354	300	355
rect	299	355	300	356
rect	299	356	300	357
rect	299	357	300	358
rect	299	358	300	359
rect	299	359	300	360
rect	299	360	300	361
rect	299	361	300	362
rect	299	362	300	363
rect	299	363	300	364
rect	299	364	300	365
rect	299	365	300	366
rect	337	0	338	1
rect	337	1	338	2
rect	337	2	338	3
rect	337	3	338	4
rect	337	4	338	5
rect	337	5	338	6
rect	337	6	338	7
rect	337	7	338	8
rect	337	8	338	9
rect	337	9	338	10
rect	337	10	338	11
rect	337	11	338	12
rect	337	12	338	13
rect	337	13	338	14
rect	337	14	338	15
rect	337	15	338	16
rect	337	16	338	17
rect	337	17	338	18
rect	337	18	338	19
rect	337	19	338	20
rect	337	20	338	21
rect	337	21	338	22
rect	337	22	338	23
rect	337	23	338	24
rect	337	24	338	25
rect	337	25	338	26
rect	337	26	338	27
rect	337	27	338	28
rect	337	28	338	29
rect	337	29	338	30
rect	337	30	338	31
rect	337	31	338	32
rect	337	32	338	33
rect	337	33	338	34
rect	337	34	338	35
rect	337	35	338	36
rect	337	36	338	37
rect	337	37	338	38
rect	337	38	338	39
rect	337	39	338	40
rect	337	40	338	41
rect	337	41	338	42
rect	337	42	338	43
rect	337	43	338	44
rect	337	44	338	45
rect	337	45	338	46
rect	337	46	338	47
rect	337	47	338	48
rect	337	48	338	49
rect	337	49	338	50
rect	337	50	338	51
rect	337	51	338	52
rect	337	52	338	53
rect	337	53	338	54
rect	337	54	338	55
rect	337	55	338	56
rect	337	56	338	57
rect	337	57	338	58
rect	337	58	338	59
rect	337	59	338	60
rect	337	60	338	61
rect	337	61	338	62
rect	337	62	338	63
rect	337	63	338	64
rect	337	64	338	65
rect	337	65	338	66
rect	337	66	338	67
rect	337	67	338	68
rect	337	68	338	69
rect	337	69	338	70
rect	337	70	338	71
rect	337	71	338	72
rect	337	72	338	73
rect	337	73	338	74
rect	337	74	338	75
rect	337	75	338	76
rect	337	76	338	77
rect	337	77	338	78
rect	337	78	338	79
rect	337	79	338	80
rect	337	80	338	81
rect	337	81	338	82
rect	337	82	338	83
rect	337	83	338	84
rect	337	84	338	85
rect	337	85	338	86
rect	337	86	338	87
rect	337	87	338	88
rect	337	88	338	89
rect	337	89	338	90
rect	337	90	338	91
rect	337	91	338	92
rect	337	92	338	93
rect	337	93	338	94
rect	337	94	338	95
rect	337	95	338	96
rect	337	96	338	97
rect	337	97	338	98
rect	337	98	338	99
rect	337	99	338	100
rect	337	100	338	101
rect	337	101	338	102
rect	337	102	338	103
rect	337	103	338	104
rect	337	104	338	105
rect	337	105	338	106
rect	337	106	338	107
rect	337	107	338	108
rect	337	108	338	109
rect	337	109	338	110
rect	337	110	338	111
rect	337	111	338	112
rect	337	112	338	113
rect	337	113	338	114
rect	337	114	338	115
rect	337	115	338	116
rect	337	116	338	117
rect	337	117	338	118
rect	337	118	338	119
rect	337	119	338	120
rect	337	120	338	121
rect	337	121	338	122
rect	337	122	338	123
rect	337	123	338	124
rect	337	124	338	125
rect	337	125	338	126
rect	337	126	338	127
rect	337	127	338	128
rect	337	128	338	129
rect	337	129	338	130
rect	337	130	338	131
rect	337	131	338	132
rect	337	132	338	133
rect	337	133	338	134
rect	337	134	338	135
rect	337	135	338	136
rect	337	136	338	137
rect	337	137	338	138
rect	337	138	338	139
rect	337	139	338	140
rect	337	140	338	141
rect	337	141	338	142
rect	337	142	338	143
rect	337	143	338	144
rect	337	144	338	145
rect	337	145	338	146
rect	337	146	338	147
rect	337	147	338	148
rect	337	148	338	149
rect	337	149	338	150
rect	337	150	338	151
rect	337	151	338	152
rect	337	152	338	153
rect	337	153	338	154
rect	337	154	338	155
rect	337	155	338	156
rect	337	156	338	157
rect	337	157	338	158
rect	337	158	338	159
rect	337	159	338	160
rect	337	160	338	161
rect	337	161	338	162
rect	337	162	338	163
rect	337	163	338	164
rect	337	164	338	165
rect	337	165	338	166
rect	337	166	338	167
rect	337	167	338	168
rect	337	168	338	169
rect	337	169	338	170
rect	337	170	338	171
rect	337	171	338	172
rect	337	172	338	173
rect	337	173	338	174
rect	337	174	338	175
rect	337	175	338	176
rect	337	176	338	177
rect	337	177	338	178
rect	337	178	338	179
rect	337	179	338	180
rect	337	180	338	181
rect	337	181	338	182
rect	337	182	338	183
rect	337	183	338	184
rect	337	184	338	185
rect	337	185	338	186
rect	337	186	338	187
rect	337	187	338	188
rect	337	188	338	189
rect	337	189	338	190
rect	337	190	338	191
rect	337	191	338	192
rect	337	192	338	193
rect	337	193	338	194
rect	337	194	338	195
rect	337	195	338	196
rect	337	196	338	197
rect	337	197	338	198
rect	337	198	338	199
rect	337	199	338	200
rect	337	200	338	201
rect	337	201	338	202
rect	337	202	338	203
rect	337	203	338	204
rect	337	204	338	205
rect	337	205	338	206
rect	337	206	338	207
rect	337	207	338	208
rect	337	208	338	209
rect	337	209	338	210
rect	337	210	338	211
rect	337	211	338	212
rect	337	212	338	213
rect	337	213	338	214
rect	337	214	338	215
rect	337	215	338	216
rect	337	216	338	217
rect	337	217	338	218
rect	337	218	338	219
rect	337	219	338	220
rect	337	220	338	221
rect	337	221	338	222
rect	337	222	338	223
rect	337	223	338	224
rect	337	224	338	225
rect	337	225	338	226
rect	337	226	338	227
rect	337	227	338	228
rect	337	228	338	229
rect	337	229	338	230
rect	337	230	338	231
rect	337	231	338	232
rect	337	232	338	233
rect	337	233	338	234
rect	337	234	338	235
rect	337	235	338	236
rect	337	236	338	237
rect	337	237	338	238
rect	337	238	338	239
rect	337	239	338	240
rect	337	240	338	241
rect	337	241	338	242
rect	337	242	338	243
rect	337	243	338	244
rect	337	244	338	245
rect	337	245	338	246
rect	337	246	338	247
rect	337	247	338	248
rect	337	248	338	249
rect	337	249	338	250
rect	337	250	338	251
rect	337	251	338	252
rect	337	252	338	253
rect	337	253	338	254
rect	337	254	338	255
rect	337	255	338	256
rect	337	256	338	257
rect	337	257	338	258
rect	337	258	338	259
rect	337	259	338	260
rect	337	260	338	261
rect	337	261	338	262
rect	337	262	338	263
rect	337	263	338	264
rect	337	264	338	265
rect	337	265	338	266
rect	337	266	338	267
rect	337	267	338	268
rect	337	268	338	269
rect	337	269	338	270
rect	337	270	338	271
rect	337	271	338	272
rect	337	272	338	273
rect	337	273	338	274
rect	337	274	338	275
rect	337	275	338	276
rect	337	276	338	277
rect	337	277	338	278
rect	337	278	338	279
rect	337	279	338	280
rect	337	280	338	281
rect	337	281	338	282
rect	337	282	338	283
rect	337	283	338	284
rect	337	284	338	285
rect	337	285	338	286
rect	337	286	338	287
rect	337	287	338	288
rect	337	288	338	289
rect	337	289	338	290
rect	337	290	338	291
rect	337	291	338	292
rect	337	292	338	293
rect	337	293	338	294
rect	337	294	338	295
rect	337	295	338	296
rect	337	296	338	297
rect	337	297	338	298
rect	337	298	338	299
rect	337	299	338	300
rect	337	300	338	301
rect	337	301	338	302
rect	337	302	338	303
rect	337	303	338	304
rect	337	304	338	305
rect	337	305	338	306
rect	337	306	338	307
rect	337	307	338	308
rect	337	308	338	309
rect	337	309	338	310
rect	337	310	338	311
rect	337	311	338	312
rect	337	312	338	313
rect	337	313	338	314
rect	337	314	338	315
rect	337	315	338	316
rect	337	316	338	317
rect	337	317	338	318
rect	337	318	338	319
rect	337	319	338	320
rect	337	320	338	321
rect	337	321	338	322
rect	337	322	338	323
rect	337	323	338	324
rect	337	324	338	325
rect	337	325	338	326
rect	337	326	338	327
rect	337	327	338	328
rect	337	328	338	329
rect	337	329	338	330
rect	337	330	338	331
rect	337	331	338	332
rect	337	332	338	333
rect	337	333	338	334
rect	337	334	338	335
rect	337	335	338	336
rect	337	336	338	337
rect	337	337	338	338
rect	337	338	338	339
rect	337	339	338	340
rect	337	340	338	341
rect	337	341	338	342
rect	337	342	338	343
rect	337	343	338	344
rect	337	344	338	345
rect	337	345	338	346
rect	337	346	338	347
rect	337	347	338	348
rect	337	348	338	349
rect	337	349	338	350
rect	337	350	338	351
rect	337	351	338	352
rect	337	352	338	353
rect	337	353	338	354
rect	337	354	338	355
rect	337	355	338	356
rect	337	356	338	357
rect	337	357	338	358
rect	337	358	338	359
rect	337	359	338	360
rect	337	360	338	361
rect	337	361	338	362
rect	337	362	338	363
rect	337	363	338	364
rect	337	364	338	365
rect	337	365	338	366
rect	337	366	338	367
rect	337	367	338	368
rect	337	368	338	369
rect	337	369	338	370
rect	337	370	338	371
rect	337	371	338	372
rect	337	372	338	373
rect	337	373	338	374
rect	337	374	338	375
rect	337	375	338	376
rect	337	376	338	377
rect	337	377	338	378
rect	337	378	338	379
rect	337	379	338	380
rect	337	380	338	381
rect	337	381	338	382
rect	337	382	338	383
rect	337	383	338	384
rect	337	384	338	385
rect	337	385	338	386
rect	337	386	338	387
rect	338	0	339	1
rect	338	1	339	2
rect	338	2	339	3
rect	338	3	339	4
rect	338	4	339	5
rect	338	5	339	6
rect	338	6	339	7
rect	338	7	339	8
rect	338	8	339	9
rect	338	9	339	10
rect	338	10	339	11
rect	338	11	339	12
rect	338	12	339	13
rect	338	13	339	14
rect	338	14	339	15
rect	338	15	339	16
rect	338	16	339	17
rect	338	17	339	18
rect	338	18	339	19
rect	338	19	339	20
rect	338	20	339	21
rect	338	21	339	22
rect	338	22	339	23
rect	338	23	339	24
rect	338	24	339	25
rect	338	25	339	26
rect	338	26	339	27
rect	338	27	339	28
rect	338	28	339	29
rect	338	29	339	30
rect	338	30	339	31
rect	338	31	339	32
rect	338	32	339	33
rect	338	33	339	34
rect	338	34	339	35
rect	338	35	339	36
rect	338	36	339	37
rect	338	37	339	38
rect	338	38	339	39
rect	338	39	339	40
rect	338	40	339	41
rect	338	41	339	42
rect	338	42	339	43
rect	338	43	339	44
rect	338	44	339	45
rect	338	45	339	46
rect	338	46	339	47
rect	338	47	339	48
rect	338	48	339	49
rect	338	49	339	50
rect	338	50	339	51
rect	338	51	339	52
rect	338	52	339	53
rect	338	53	339	54
rect	338	54	339	55
rect	338	55	339	56
rect	338	56	339	57
rect	338	57	339	58
rect	338	58	339	59
rect	338	59	339	60
rect	338	60	339	61
rect	338	61	339	62
rect	338	62	339	63
rect	338	63	339	64
rect	338	64	339	65
rect	338	65	339	66
rect	338	66	339	67
rect	338	67	339	68
rect	338	68	339	69
rect	338	69	339	70
rect	338	70	339	71
rect	338	71	339	72
rect	338	72	339	73
rect	338	73	339	74
rect	338	74	339	75
rect	338	75	339	76
rect	338	76	339	77
rect	338	77	339	78
rect	338	78	339	79
rect	338	79	339	80
rect	338	80	339	81
rect	338	81	339	82
rect	338	82	339	83
rect	338	83	339	84
rect	338	84	339	85
rect	338	85	339	86
rect	338	86	339	87
rect	338	87	339	88
rect	338	88	339	89
rect	338	89	339	90
rect	338	90	339	91
rect	338	91	339	92
rect	338	92	339	93
rect	338	93	339	94
rect	338	94	339	95
rect	338	95	339	96
rect	338	96	339	97
rect	338	97	339	98
rect	338	98	339	99
rect	338	99	339	100
rect	338	100	339	101
rect	338	101	339	102
rect	338	102	339	103
rect	338	103	339	104
rect	338	104	339	105
rect	338	105	339	106
rect	338	106	339	107
rect	338	107	339	108
rect	338	108	339	109
rect	338	109	339	110
rect	338	110	339	111
rect	338	111	339	112
rect	338	112	339	113
rect	338	113	339	114
rect	338	114	339	115
rect	338	115	339	116
rect	338	116	339	117
rect	338	117	339	118
rect	338	118	339	119
rect	338	119	339	120
rect	338	120	339	121
rect	338	121	339	122
rect	338	122	339	123
rect	338	123	339	124
rect	338	124	339	125
rect	338	125	339	126
rect	338	126	339	127
rect	338	127	339	128
rect	338	128	339	129
rect	338	129	339	130
rect	338	130	339	131
rect	338	131	339	132
rect	338	132	339	133
rect	338	133	339	134
rect	338	134	339	135
rect	338	135	339	136
rect	338	136	339	137
rect	338	137	339	138
rect	338	138	339	139
rect	338	139	339	140
rect	338	140	339	141
rect	338	141	339	142
rect	338	142	339	143
rect	338	143	339	144
rect	338	144	339	145
rect	338	145	339	146
rect	338	146	339	147
rect	338	147	339	148
rect	338	148	339	149
rect	338	149	339	150
rect	338	150	339	151
rect	338	151	339	152
rect	338	152	339	153
rect	338	153	339	154
rect	338	154	339	155
rect	338	155	339	156
rect	338	156	339	157
rect	338	157	339	158
rect	338	158	339	159
rect	338	159	339	160
rect	338	160	339	161
rect	338	161	339	162
rect	338	162	339	163
rect	338	163	339	164
rect	338	164	339	165
rect	338	165	339	166
rect	338	166	339	167
rect	338	167	339	168
rect	338	168	339	169
rect	338	169	339	170
rect	338	170	339	171
rect	338	171	339	172
rect	338	172	339	173
rect	338	173	339	174
rect	338	174	339	175
rect	338	175	339	176
rect	338	176	339	177
rect	338	177	339	178
rect	338	178	339	179
rect	338	179	339	180
rect	338	180	339	181
rect	338	181	339	182
rect	338	182	339	183
rect	338	183	339	184
rect	338	184	339	185
rect	338	185	339	186
rect	338	186	339	187
rect	338	187	339	188
rect	338	188	339	189
rect	338	189	339	190
rect	338	190	339	191
rect	338	191	339	192
rect	338	192	339	193
rect	338	193	339	194
rect	338	194	339	195
rect	338	195	339	196
rect	338	196	339	197
rect	338	197	339	198
rect	338	198	339	199
rect	338	199	339	200
rect	338	200	339	201
rect	338	201	339	202
rect	338	202	339	203
rect	338	203	339	204
rect	338	204	339	205
rect	338	205	339	206
rect	338	206	339	207
rect	338	207	339	208
rect	338	208	339	209
rect	338	209	339	210
rect	338	210	339	211
rect	338	211	339	212
rect	338	212	339	213
rect	338	213	339	214
rect	338	214	339	215
rect	338	215	339	216
rect	338	216	339	217
rect	338	217	339	218
rect	338	218	339	219
rect	338	219	339	220
rect	338	220	339	221
rect	338	221	339	222
rect	338	222	339	223
rect	338	223	339	224
rect	338	224	339	225
rect	338	225	339	226
rect	338	226	339	227
rect	338	227	339	228
rect	338	228	339	229
rect	338	229	339	230
rect	338	230	339	231
rect	338	231	339	232
rect	338	232	339	233
rect	338	233	339	234
rect	338	234	339	235
rect	338	235	339	236
rect	338	236	339	237
rect	338	237	339	238
rect	338	238	339	239
rect	338	239	339	240
rect	338	240	339	241
rect	338	241	339	242
rect	338	242	339	243
rect	338	243	339	244
rect	338	244	339	245
rect	338	245	339	246
rect	338	246	339	247
rect	338	247	339	248
rect	338	248	339	249
rect	338	249	339	250
rect	338	250	339	251
rect	338	251	339	252
rect	338	252	339	253
rect	338	253	339	254
rect	338	254	339	255
rect	338	255	339	256
rect	338	256	339	257
rect	338	257	339	258
rect	338	258	339	259
rect	338	259	339	260
rect	338	260	339	261
rect	338	261	339	262
rect	338	262	339	263
rect	338	263	339	264
rect	338	264	339	265
rect	338	265	339	266
rect	338	266	339	267
rect	338	267	339	268
rect	338	268	339	269
rect	338	269	339	270
rect	338	270	339	271
rect	338	271	339	272
rect	338	272	339	273
rect	338	273	339	274
rect	338	274	339	275
rect	338	275	339	276
rect	338	276	339	277
rect	338	277	339	278
rect	338	278	339	279
rect	338	279	339	280
rect	338	280	339	281
rect	338	281	339	282
rect	338	282	339	283
rect	338	283	339	284
rect	338	284	339	285
rect	338	285	339	286
rect	338	286	339	287
rect	338	287	339	288
rect	338	288	339	289
rect	338	289	339	290
rect	338	290	339	291
rect	338	291	339	292
rect	338	292	339	293
rect	338	293	339	294
rect	338	294	339	295
rect	338	295	339	296
rect	338	296	339	297
rect	338	297	339	298
rect	338	298	339	299
rect	338	299	339	300
rect	338	300	339	301
rect	338	301	339	302
rect	338	302	339	303
rect	338	303	339	304
rect	338	304	339	305
rect	338	305	339	306
rect	338	306	339	307
rect	338	307	339	308
rect	338	308	339	309
rect	338	309	339	310
rect	338	310	339	311
rect	338	311	339	312
rect	338	312	339	313
rect	338	313	339	314
rect	338	314	339	315
rect	338	315	339	316
rect	338	316	339	317
rect	338	317	339	318
rect	338	318	339	319
rect	338	319	339	320
rect	338	320	339	321
rect	338	321	339	322
rect	338	322	339	323
rect	338	323	339	324
rect	338	324	339	325
rect	338	325	339	326
rect	338	326	339	327
rect	338	327	339	328
rect	338	328	339	329
rect	338	329	339	330
rect	338	330	339	331
rect	338	331	339	332
rect	338	332	339	333
rect	338	333	339	334
rect	338	334	339	335
rect	338	335	339	336
rect	338	336	339	337
rect	338	337	339	338
rect	338	338	339	339
rect	338	339	339	340
rect	338	340	339	341
rect	338	341	339	342
rect	338	342	339	343
rect	338	343	339	344
rect	338	344	339	345
rect	338	345	339	346
rect	338	346	339	347
rect	338	347	339	348
rect	338	348	339	349
rect	338	349	339	350
rect	338	350	339	351
rect	338	351	339	352
rect	338	352	339	353
rect	338	353	339	354
rect	338	354	339	355
rect	338	355	339	356
rect	338	356	339	357
rect	338	357	339	358
rect	338	358	339	359
rect	338	359	339	360
rect	338	360	339	361
rect	338	361	339	362
rect	338	362	339	363
rect	338	363	339	364
rect	338	364	339	365
rect	338	365	339	366
rect	338	366	339	367
rect	338	367	339	368
rect	338	368	339	369
rect	338	369	339	370
rect	338	370	339	371
rect	338	371	339	372
rect	338	372	339	373
rect	338	373	339	374
rect	338	374	339	375
rect	338	375	339	376
rect	338	376	339	377
rect	338	377	339	378
rect	338	378	339	379
rect	338	379	339	380
rect	338	380	339	381
rect	338	381	339	382
rect	338	382	339	383
rect	338	383	339	384
rect	338	384	339	385
rect	338	385	339	386
rect	338	386	339	387
rect	339	0	340	1
rect	339	1	340	2
rect	339	2	340	3
rect	339	3	340	4
rect	339	4	340	5
rect	339	5	340	6
rect	339	6	340	7
rect	339	7	340	8
rect	339	8	340	9
rect	339	9	340	10
rect	339	10	340	11
rect	339	11	340	12
rect	339	12	340	13
rect	339	13	340	14
rect	339	14	340	15
rect	339	15	340	16
rect	339	16	340	17
rect	339	17	340	18
rect	339	18	340	19
rect	339	19	340	20
rect	339	20	340	21
rect	339	21	340	22
rect	339	22	340	23
rect	339	23	340	24
rect	339	24	340	25
rect	339	25	340	26
rect	339	26	340	27
rect	339	27	340	28
rect	339	28	340	29
rect	339	29	340	30
rect	339	30	340	31
rect	339	31	340	32
rect	339	32	340	33
rect	339	33	340	34
rect	339	34	340	35
rect	339	35	340	36
rect	339	36	340	37
rect	339	37	340	38
rect	339	38	340	39
rect	339	39	340	40
rect	339	40	340	41
rect	339	41	340	42
rect	339	42	340	43
rect	339	43	340	44
rect	339	44	340	45
rect	339	45	340	46
rect	339	46	340	47
rect	339	47	340	48
rect	339	48	340	49
rect	339	49	340	50
rect	339	50	340	51
rect	339	51	340	52
rect	339	52	340	53
rect	339	53	340	54
rect	339	54	340	55
rect	339	55	340	56
rect	339	56	340	57
rect	339	57	340	58
rect	339	58	340	59
rect	339	59	340	60
rect	339	60	340	61
rect	339	61	340	62
rect	339	62	340	63
rect	339	63	340	64
rect	339	64	340	65
rect	339	65	340	66
rect	339	66	340	67
rect	339	67	340	68
rect	339	68	340	69
rect	339	69	340	70
rect	339	70	340	71
rect	339	71	340	72
rect	339	72	340	73
rect	339	73	340	74
rect	339	74	340	75
rect	339	75	340	76
rect	339	76	340	77
rect	339	77	340	78
rect	339	78	340	79
rect	339	79	340	80
rect	339	80	340	81
rect	339	81	340	82
rect	339	82	340	83
rect	339	83	340	84
rect	339	84	340	85
rect	339	85	340	86
rect	339	86	340	87
rect	339	87	340	88
rect	339	88	340	89
rect	339	89	340	90
rect	339	90	340	91
rect	339	91	340	92
rect	339	92	340	93
rect	339	93	340	94
rect	339	94	340	95
rect	339	95	340	96
rect	339	96	340	97
rect	339	97	340	98
rect	339	98	340	99
rect	339	99	340	100
rect	339	100	340	101
rect	339	101	340	102
rect	339	102	340	103
rect	339	103	340	104
rect	339	104	340	105
rect	339	105	340	106
rect	339	106	340	107
rect	339	107	340	108
rect	339	108	340	109
rect	339	109	340	110
rect	339	110	340	111
rect	339	111	340	112
rect	339	112	340	113
rect	339	113	340	114
rect	339	114	340	115
rect	339	115	340	116
rect	339	116	340	117
rect	339	117	340	118
rect	339	118	340	119
rect	339	119	340	120
rect	339	120	340	121
rect	339	121	340	122
rect	339	122	340	123
rect	339	123	340	124
rect	339	124	340	125
rect	339	125	340	126
rect	339	126	340	127
rect	339	127	340	128
rect	339	128	340	129
rect	339	129	340	130
rect	339	130	340	131
rect	339	131	340	132
rect	339	132	340	133
rect	339	133	340	134
rect	339	134	340	135
rect	339	135	340	136
rect	339	136	340	137
rect	339	137	340	138
rect	339	138	340	139
rect	339	139	340	140
rect	339	140	340	141
rect	339	141	340	142
rect	339	142	340	143
rect	339	143	340	144
rect	339	144	340	145
rect	339	145	340	146
rect	339	146	340	147
rect	339	147	340	148
rect	339	148	340	149
rect	339	149	340	150
rect	339	150	340	151
rect	339	151	340	152
rect	339	152	340	153
rect	339	153	340	154
rect	339	154	340	155
rect	339	155	340	156
rect	339	156	340	157
rect	339	157	340	158
rect	339	158	340	159
rect	339	159	340	160
rect	339	160	340	161
rect	339	161	340	162
rect	339	162	340	163
rect	339	163	340	164
rect	339	164	340	165
rect	339	165	340	166
rect	339	166	340	167
rect	339	167	340	168
rect	339	168	340	169
rect	339	169	340	170
rect	339	170	340	171
rect	339	171	340	172
rect	339	172	340	173
rect	339	173	340	174
rect	339	174	340	175
rect	339	175	340	176
rect	339	176	340	177
rect	339	177	340	178
rect	339	178	340	179
rect	339	179	340	180
rect	339	180	340	181
rect	339	181	340	182
rect	339	182	340	183
rect	339	183	340	184
rect	339	184	340	185
rect	339	185	340	186
rect	339	186	340	187
rect	339	187	340	188
rect	339	188	340	189
rect	339	189	340	190
rect	339	190	340	191
rect	339	191	340	192
rect	339	192	340	193
rect	339	193	340	194
rect	339	194	340	195
rect	339	195	340	196
rect	339	196	340	197
rect	339	197	340	198
rect	339	198	340	199
rect	339	199	340	200
rect	339	200	340	201
rect	339	201	340	202
rect	339	202	340	203
rect	339	203	340	204
rect	339	204	340	205
rect	339	205	340	206
rect	339	206	340	207
rect	339	207	340	208
rect	339	208	340	209
rect	339	209	340	210
rect	339	210	340	211
rect	339	211	340	212
rect	339	212	340	213
rect	339	213	340	214
rect	339	214	340	215
rect	339	215	340	216
rect	339	216	340	217
rect	339	217	340	218
rect	339	218	340	219
rect	339	219	340	220
rect	339	220	340	221
rect	339	221	340	222
rect	339	222	340	223
rect	339	223	340	224
rect	339	224	340	225
rect	339	225	340	226
rect	339	226	340	227
rect	339	227	340	228
rect	339	228	340	229
rect	339	229	340	230
rect	339	230	340	231
rect	339	231	340	232
rect	339	232	340	233
rect	339	233	340	234
rect	339	234	340	235
rect	339	235	340	236
rect	339	236	340	237
rect	339	237	340	238
rect	339	238	340	239
rect	339	239	340	240
rect	339	240	340	241
rect	339	241	340	242
rect	339	242	340	243
rect	339	243	340	244
rect	339	244	340	245
rect	339	245	340	246
rect	339	246	340	247
rect	339	247	340	248
rect	339	248	340	249
rect	339	249	340	250
rect	339	250	340	251
rect	339	251	340	252
rect	339	252	340	253
rect	339	253	340	254
rect	339	254	340	255
rect	339	255	340	256
rect	339	256	340	257
rect	339	257	340	258
rect	339	258	340	259
rect	339	259	340	260
rect	339	260	340	261
rect	339	261	340	262
rect	339	262	340	263
rect	339	263	340	264
rect	339	264	340	265
rect	339	265	340	266
rect	339	266	340	267
rect	339	267	340	268
rect	339	268	340	269
rect	339	269	340	270
rect	339	270	340	271
rect	339	271	340	272
rect	339	272	340	273
rect	339	273	340	274
rect	339	274	340	275
rect	339	275	340	276
rect	339	276	340	277
rect	339	277	340	278
rect	339	278	340	279
rect	339	279	340	280
rect	339	280	340	281
rect	339	281	340	282
rect	339	282	340	283
rect	339	283	340	284
rect	339	284	340	285
rect	339	285	340	286
rect	339	286	340	287
rect	339	287	340	288
rect	339	288	340	289
rect	339	289	340	290
rect	339	290	340	291
rect	339	291	340	292
rect	339	292	340	293
rect	339	293	340	294
rect	339	294	340	295
rect	339	295	340	296
rect	339	296	340	297
rect	339	297	340	298
rect	339	298	340	299
rect	339	299	340	300
rect	339	300	340	301
rect	339	301	340	302
rect	339	302	340	303
rect	339	303	340	304
rect	339	304	340	305
rect	339	305	340	306
rect	339	306	340	307
rect	339	307	340	308
rect	339	308	340	309
rect	339	309	340	310
rect	339	310	340	311
rect	339	311	340	312
rect	339	312	340	313
rect	339	313	340	314
rect	339	314	340	315
rect	339	315	340	316
rect	339	316	340	317
rect	339	317	340	318
rect	339	318	340	319
rect	339	319	340	320
rect	339	320	340	321
rect	339	321	340	322
rect	339	322	340	323
rect	339	323	340	324
rect	339	324	340	325
rect	339	325	340	326
rect	339	326	340	327
rect	339	327	340	328
rect	339	328	340	329
rect	339	329	340	330
rect	339	330	340	331
rect	339	331	340	332
rect	339	332	340	333
rect	339	333	340	334
rect	339	334	340	335
rect	339	335	340	336
rect	339	336	340	337
rect	339	337	340	338
rect	339	338	340	339
rect	339	339	340	340
rect	339	340	340	341
rect	339	341	340	342
rect	339	342	340	343
rect	339	343	340	344
rect	339	344	340	345
rect	339	345	340	346
rect	339	346	340	347
rect	339	347	340	348
rect	339	348	340	349
rect	339	349	340	350
rect	339	350	340	351
rect	339	351	340	352
rect	339	352	340	353
rect	339	353	340	354
rect	339	354	340	355
rect	339	355	340	356
rect	339	356	340	357
rect	339	357	340	358
rect	339	358	340	359
rect	339	359	340	360
rect	339	360	340	361
rect	339	361	340	362
rect	339	362	340	363
rect	339	363	340	364
rect	339	364	340	365
rect	339	365	340	366
rect	339	366	340	367
rect	339	367	340	368
rect	339	368	340	369
rect	339	369	340	370
rect	339	370	340	371
rect	339	371	340	372
rect	339	372	340	373
rect	339	373	340	374
rect	339	374	340	375
rect	339	375	340	376
rect	339	376	340	377
rect	339	377	340	378
rect	339	378	340	379
rect	339	379	340	380
rect	339	380	340	381
rect	339	381	340	382
rect	339	382	340	383
rect	339	383	340	384
rect	339	384	340	385
rect	339	385	340	386
rect	339	386	340	387
rect	340	0	341	1
rect	340	1	341	2
rect	340	2	341	3
rect	340	3	341	4
rect	340	4	341	5
rect	340	5	341	6
rect	340	6	341	7
rect	340	7	341	8
rect	340	8	341	9
rect	340	9	341	10
rect	340	10	341	11
rect	340	11	341	12
rect	340	12	341	13
rect	340	13	341	14
rect	340	14	341	15
rect	340	15	341	16
rect	340	16	341	17
rect	340	17	341	18
rect	340	18	341	19
rect	340	19	341	20
rect	340	20	341	21
rect	340	21	341	22
rect	340	22	341	23
rect	340	23	341	24
rect	340	24	341	25
rect	340	25	341	26
rect	340	26	341	27
rect	340	27	341	28
rect	340	28	341	29
rect	340	29	341	30
rect	340	30	341	31
rect	340	31	341	32
rect	340	32	341	33
rect	340	33	341	34
rect	340	34	341	35
rect	340	35	341	36
rect	340	36	341	37
rect	340	37	341	38
rect	340	38	341	39
rect	340	39	341	40
rect	340	40	341	41
rect	340	41	341	42
rect	340	42	341	43
rect	340	43	341	44
rect	340	44	341	45
rect	340	45	341	46
rect	340	46	341	47
rect	340	47	341	48
rect	340	48	341	49
rect	340	49	341	50
rect	340	50	341	51
rect	340	51	341	52
rect	340	52	341	53
rect	340	53	341	54
rect	340	54	341	55
rect	340	55	341	56
rect	340	56	341	57
rect	340	57	341	58
rect	340	58	341	59
rect	340	59	341	60
rect	340	60	341	61
rect	340	61	341	62
rect	340	62	341	63
rect	340	63	341	64
rect	340	64	341	65
rect	340	65	341	66
rect	340	66	341	67
rect	340	67	341	68
rect	340	68	341	69
rect	340	69	341	70
rect	340	70	341	71
rect	340	71	341	72
rect	340	72	341	73
rect	340	73	341	74
rect	340	74	341	75
rect	340	75	341	76
rect	340	76	341	77
rect	340	77	341	78
rect	340	78	341	79
rect	340	79	341	80
rect	340	80	341	81
rect	340	81	341	82
rect	340	82	341	83
rect	340	83	341	84
rect	340	84	341	85
rect	340	85	341	86
rect	340	86	341	87
rect	340	87	341	88
rect	340	88	341	89
rect	340	89	341	90
rect	340	90	341	91
rect	340	91	341	92
rect	340	92	341	93
rect	340	93	341	94
rect	340	94	341	95
rect	340	95	341	96
rect	340	96	341	97
rect	340	97	341	98
rect	340	98	341	99
rect	340	99	341	100
rect	340	100	341	101
rect	340	101	341	102
rect	340	102	341	103
rect	340	103	341	104
rect	340	104	341	105
rect	340	105	341	106
rect	340	106	341	107
rect	340	107	341	108
rect	340	108	341	109
rect	340	109	341	110
rect	340	110	341	111
rect	340	111	341	112
rect	340	112	341	113
rect	340	113	341	114
rect	340	114	341	115
rect	340	115	341	116
rect	340	116	341	117
rect	340	117	341	118
rect	340	118	341	119
rect	340	119	341	120
rect	340	120	341	121
rect	340	121	341	122
rect	340	122	341	123
rect	340	123	341	124
rect	340	124	341	125
rect	340	125	341	126
rect	340	126	341	127
rect	340	127	341	128
rect	340	128	341	129
rect	340	129	341	130
rect	340	130	341	131
rect	340	131	341	132
rect	340	132	341	133
rect	340	133	341	134
rect	340	134	341	135
rect	340	135	341	136
rect	340	136	341	137
rect	340	137	341	138
rect	340	138	341	139
rect	340	139	341	140
rect	340	140	341	141
rect	340	141	341	142
rect	340	142	341	143
rect	340	143	341	144
rect	340	144	341	145
rect	340	145	341	146
rect	340	146	341	147
rect	340	147	341	148
rect	340	148	341	149
rect	340	149	341	150
rect	340	150	341	151
rect	340	151	341	152
rect	340	152	341	153
rect	340	153	341	154
rect	340	154	341	155
rect	340	155	341	156
rect	340	156	341	157
rect	340	157	341	158
rect	340	158	341	159
rect	340	159	341	160
rect	340	160	341	161
rect	340	161	341	162
rect	340	162	341	163
rect	340	163	341	164
rect	340	164	341	165
rect	340	165	341	166
rect	340	166	341	167
rect	340	167	341	168
rect	340	168	341	169
rect	340	169	341	170
rect	340	170	341	171
rect	340	171	341	172
rect	340	172	341	173
rect	340	173	341	174
rect	340	174	341	175
rect	340	175	341	176
rect	340	176	341	177
rect	340	177	341	178
rect	340	178	341	179
rect	340	179	341	180
rect	340	180	341	181
rect	340	181	341	182
rect	340	182	341	183
rect	340	183	341	184
rect	340	184	341	185
rect	340	185	341	186
rect	340	186	341	187
rect	340	187	341	188
rect	340	188	341	189
rect	340	189	341	190
rect	340	190	341	191
rect	340	191	341	192
rect	340	192	341	193
rect	340	193	341	194
rect	340	194	341	195
rect	340	195	341	196
rect	340	196	341	197
rect	340	197	341	198
rect	340	198	341	199
rect	340	199	341	200
rect	340	200	341	201
rect	340	201	341	202
rect	340	202	341	203
rect	340	203	341	204
rect	340	204	341	205
rect	340	205	341	206
rect	340	206	341	207
rect	340	207	341	208
rect	340	208	341	209
rect	340	209	341	210
rect	340	210	341	211
rect	340	211	341	212
rect	340	212	341	213
rect	340	213	341	214
rect	340	214	341	215
rect	340	215	341	216
rect	340	216	341	217
rect	340	217	341	218
rect	340	218	341	219
rect	340	219	341	220
rect	340	220	341	221
rect	340	221	341	222
rect	340	222	341	223
rect	340	223	341	224
rect	340	224	341	225
rect	340	225	341	226
rect	340	226	341	227
rect	340	227	341	228
rect	340	228	341	229
rect	340	229	341	230
rect	340	230	341	231
rect	340	231	341	232
rect	340	232	341	233
rect	340	233	341	234
rect	340	234	341	235
rect	340	235	341	236
rect	340	236	341	237
rect	340	237	341	238
rect	340	238	341	239
rect	340	239	341	240
rect	340	240	341	241
rect	340	241	341	242
rect	340	242	341	243
rect	340	243	341	244
rect	340	244	341	245
rect	340	245	341	246
rect	340	246	341	247
rect	340	247	341	248
rect	340	248	341	249
rect	340	249	341	250
rect	340	250	341	251
rect	340	251	341	252
rect	340	252	341	253
rect	340	253	341	254
rect	340	254	341	255
rect	340	255	341	256
rect	340	256	341	257
rect	340	257	341	258
rect	340	258	341	259
rect	340	259	341	260
rect	340	260	341	261
rect	340	261	341	262
rect	340	262	341	263
rect	340	263	341	264
rect	340	264	341	265
rect	340	265	341	266
rect	340	266	341	267
rect	340	267	341	268
rect	340	268	341	269
rect	340	269	341	270
rect	340	270	341	271
rect	340	271	341	272
rect	340	272	341	273
rect	340	273	341	274
rect	340	274	341	275
rect	340	275	341	276
rect	340	276	341	277
rect	340	277	341	278
rect	340	278	341	279
rect	340	279	341	280
rect	340	280	341	281
rect	340	281	341	282
rect	340	282	341	283
rect	340	283	341	284
rect	340	284	341	285
rect	340	285	341	286
rect	340	286	341	287
rect	340	287	341	288
rect	340	288	341	289
rect	340	289	341	290
rect	340	290	341	291
rect	340	291	341	292
rect	340	292	341	293
rect	340	293	341	294
rect	340	294	341	295
rect	340	295	341	296
rect	340	296	341	297
rect	340	297	341	298
rect	340	298	341	299
rect	340	299	341	300
rect	340	300	341	301
rect	340	301	341	302
rect	340	302	341	303
rect	340	303	341	304
rect	340	304	341	305
rect	340	305	341	306
rect	340	306	341	307
rect	340	307	341	308
rect	340	308	341	309
rect	340	309	341	310
rect	340	310	341	311
rect	340	311	341	312
rect	340	312	341	313
rect	340	313	341	314
rect	340	314	341	315
rect	340	315	341	316
rect	340	316	341	317
rect	340	317	341	318
rect	340	318	341	319
rect	340	319	341	320
rect	340	320	341	321
rect	340	321	341	322
rect	340	322	341	323
rect	340	323	341	324
rect	340	324	341	325
rect	340	325	341	326
rect	340	326	341	327
rect	340	327	341	328
rect	340	328	341	329
rect	340	329	341	330
rect	340	330	341	331
rect	340	331	341	332
rect	340	332	341	333
rect	340	333	341	334
rect	340	334	341	335
rect	340	335	341	336
rect	340	336	341	337
rect	340	337	341	338
rect	340	338	341	339
rect	340	339	341	340
rect	340	340	341	341
rect	340	341	341	342
rect	340	342	341	343
rect	340	343	341	344
rect	340	344	341	345
rect	340	345	341	346
rect	340	346	341	347
rect	340	347	341	348
rect	340	348	341	349
rect	340	349	341	350
rect	340	350	341	351
rect	340	351	341	352
rect	340	352	341	353
rect	340	353	341	354
rect	340	354	341	355
rect	340	355	341	356
rect	340	356	341	357
rect	340	357	341	358
rect	340	358	341	359
rect	340	359	341	360
rect	340	360	341	361
rect	340	361	341	362
rect	340	362	341	363
rect	340	363	341	364
rect	340	364	341	365
rect	340	365	341	366
rect	340	366	341	367
rect	340	367	341	368
rect	340	368	341	369
rect	340	369	341	370
rect	340	370	341	371
rect	340	371	341	372
rect	340	372	341	373
rect	340	373	341	374
rect	340	374	341	375
rect	340	375	341	376
rect	340	376	341	377
rect	340	377	341	378
rect	340	378	341	379
rect	340	379	341	380
rect	340	380	341	381
rect	340	381	341	382
rect	340	382	341	383
rect	340	383	341	384
rect	340	384	341	385
rect	340	385	341	386
rect	340	386	341	387
rect	341	0	342	1
rect	341	1	342	2
rect	341	2	342	3
rect	341	3	342	4
rect	341	4	342	5
rect	341	5	342	6
rect	341	6	342	7
rect	341	7	342	8
rect	341	8	342	9
rect	341	9	342	10
rect	341	10	342	11
rect	341	11	342	12
rect	341	12	342	13
rect	341	13	342	14
rect	341	14	342	15
rect	341	15	342	16
rect	341	16	342	17
rect	341	17	342	18
rect	341	18	342	19
rect	341	19	342	20
rect	341	20	342	21
rect	341	21	342	22
rect	341	22	342	23
rect	341	23	342	24
rect	341	24	342	25
rect	341	25	342	26
rect	341	26	342	27
rect	341	27	342	28
rect	341	28	342	29
rect	341	29	342	30
rect	341	30	342	31
rect	341	31	342	32
rect	341	32	342	33
rect	341	33	342	34
rect	341	34	342	35
rect	341	35	342	36
rect	341	36	342	37
rect	341	37	342	38
rect	341	38	342	39
rect	341	39	342	40
rect	341	40	342	41
rect	341	41	342	42
rect	341	42	342	43
rect	341	43	342	44
rect	341	44	342	45
rect	341	45	342	46
rect	341	46	342	47
rect	341	47	342	48
rect	341	48	342	49
rect	341	49	342	50
rect	341	50	342	51
rect	341	51	342	52
rect	341	52	342	53
rect	341	53	342	54
rect	341	54	342	55
rect	341	55	342	56
rect	341	56	342	57
rect	341	57	342	58
rect	341	58	342	59
rect	341	59	342	60
rect	341	60	342	61
rect	341	61	342	62
rect	341	62	342	63
rect	341	63	342	64
rect	341	64	342	65
rect	341	65	342	66
rect	341	66	342	67
rect	341	67	342	68
rect	341	68	342	69
rect	341	69	342	70
rect	341	70	342	71
rect	341	71	342	72
rect	341	72	342	73
rect	341	73	342	74
rect	341	74	342	75
rect	341	75	342	76
rect	341	76	342	77
rect	341	77	342	78
rect	341	78	342	79
rect	341	79	342	80
rect	341	80	342	81
rect	341	81	342	82
rect	341	82	342	83
rect	341	83	342	84
rect	341	84	342	85
rect	341	85	342	86
rect	341	86	342	87
rect	341	87	342	88
rect	341	88	342	89
rect	341	89	342	90
rect	341	90	342	91
rect	341	91	342	92
rect	341	92	342	93
rect	341	93	342	94
rect	341	94	342	95
rect	341	95	342	96
rect	341	96	342	97
rect	341	97	342	98
rect	341	98	342	99
rect	341	99	342	100
rect	341	100	342	101
rect	341	101	342	102
rect	341	102	342	103
rect	341	103	342	104
rect	341	104	342	105
rect	341	105	342	106
rect	341	106	342	107
rect	341	107	342	108
rect	341	108	342	109
rect	341	109	342	110
rect	341	110	342	111
rect	341	111	342	112
rect	341	112	342	113
rect	341	113	342	114
rect	341	114	342	115
rect	341	115	342	116
rect	341	116	342	117
rect	341	117	342	118
rect	341	118	342	119
rect	341	119	342	120
rect	341	120	342	121
rect	341	121	342	122
rect	341	122	342	123
rect	341	123	342	124
rect	341	124	342	125
rect	341	125	342	126
rect	341	126	342	127
rect	341	127	342	128
rect	341	128	342	129
rect	341	129	342	130
rect	341	130	342	131
rect	341	131	342	132
rect	341	132	342	133
rect	341	133	342	134
rect	341	134	342	135
rect	341	135	342	136
rect	341	136	342	137
rect	341	137	342	138
rect	341	138	342	139
rect	341	139	342	140
rect	341	140	342	141
rect	341	141	342	142
rect	341	142	342	143
rect	341	143	342	144
rect	341	144	342	145
rect	341	145	342	146
rect	341	146	342	147
rect	341	147	342	148
rect	341	148	342	149
rect	341	149	342	150
rect	341	150	342	151
rect	341	151	342	152
rect	341	152	342	153
rect	341	153	342	154
rect	341	154	342	155
rect	341	155	342	156
rect	341	156	342	157
rect	341	157	342	158
rect	341	158	342	159
rect	341	159	342	160
rect	341	160	342	161
rect	341	161	342	162
rect	341	162	342	163
rect	341	163	342	164
rect	341	164	342	165
rect	341	165	342	166
rect	341	166	342	167
rect	341	167	342	168
rect	341	168	342	169
rect	341	169	342	170
rect	341	170	342	171
rect	341	171	342	172
rect	341	172	342	173
rect	341	173	342	174
rect	341	174	342	175
rect	341	175	342	176
rect	341	176	342	177
rect	341	177	342	178
rect	341	178	342	179
rect	341	179	342	180
rect	341	180	342	181
rect	341	181	342	182
rect	341	182	342	183
rect	341	183	342	184
rect	341	184	342	185
rect	341	185	342	186
rect	341	186	342	187
rect	341	187	342	188
rect	341	188	342	189
rect	341	189	342	190
rect	341	190	342	191
rect	341	191	342	192
rect	341	192	342	193
rect	341	193	342	194
rect	341	194	342	195
rect	341	195	342	196
rect	341	196	342	197
rect	341	197	342	198
rect	341	198	342	199
rect	341	199	342	200
rect	341	200	342	201
rect	341	201	342	202
rect	341	202	342	203
rect	341	203	342	204
rect	341	204	342	205
rect	341	205	342	206
rect	341	206	342	207
rect	341	207	342	208
rect	341	208	342	209
rect	341	209	342	210
rect	341	210	342	211
rect	341	211	342	212
rect	341	212	342	213
rect	341	213	342	214
rect	341	214	342	215
rect	341	215	342	216
rect	341	216	342	217
rect	341	217	342	218
rect	341	218	342	219
rect	341	219	342	220
rect	341	220	342	221
rect	341	221	342	222
rect	341	222	342	223
rect	341	223	342	224
rect	341	224	342	225
rect	341	225	342	226
rect	341	226	342	227
rect	341	227	342	228
rect	341	228	342	229
rect	341	229	342	230
rect	341	230	342	231
rect	341	231	342	232
rect	341	232	342	233
rect	341	233	342	234
rect	341	234	342	235
rect	341	235	342	236
rect	341	236	342	237
rect	341	237	342	238
rect	341	238	342	239
rect	341	239	342	240
rect	341	240	342	241
rect	341	241	342	242
rect	341	242	342	243
rect	341	243	342	244
rect	341	244	342	245
rect	341	245	342	246
rect	341	246	342	247
rect	341	247	342	248
rect	341	248	342	249
rect	341	249	342	250
rect	341	250	342	251
rect	341	251	342	252
rect	341	252	342	253
rect	341	253	342	254
rect	341	254	342	255
rect	341	255	342	256
rect	341	256	342	257
rect	341	257	342	258
rect	341	258	342	259
rect	341	259	342	260
rect	341	260	342	261
rect	341	261	342	262
rect	341	262	342	263
rect	341	263	342	264
rect	341	264	342	265
rect	341	265	342	266
rect	341	266	342	267
rect	341	267	342	268
rect	341	268	342	269
rect	341	269	342	270
rect	341	270	342	271
rect	341	271	342	272
rect	341	272	342	273
rect	341	273	342	274
rect	341	274	342	275
rect	341	275	342	276
rect	341	276	342	277
rect	341	277	342	278
rect	341	278	342	279
rect	341	279	342	280
rect	341	280	342	281
rect	341	281	342	282
rect	341	282	342	283
rect	341	283	342	284
rect	341	284	342	285
rect	341	285	342	286
rect	341	286	342	287
rect	341	287	342	288
rect	341	288	342	289
rect	341	289	342	290
rect	341	290	342	291
rect	341	291	342	292
rect	341	292	342	293
rect	341	293	342	294
rect	341	294	342	295
rect	341	295	342	296
rect	341	296	342	297
rect	341	297	342	298
rect	341	298	342	299
rect	341	299	342	300
rect	341	300	342	301
rect	341	301	342	302
rect	341	302	342	303
rect	341	303	342	304
rect	341	304	342	305
rect	341	305	342	306
rect	341	306	342	307
rect	341	307	342	308
rect	341	308	342	309
rect	341	309	342	310
rect	341	310	342	311
rect	341	311	342	312
rect	341	312	342	313
rect	341	313	342	314
rect	341	314	342	315
rect	341	315	342	316
rect	341	316	342	317
rect	341	317	342	318
rect	341	318	342	319
rect	341	319	342	320
rect	341	320	342	321
rect	341	321	342	322
rect	341	322	342	323
rect	341	323	342	324
rect	341	324	342	325
rect	341	325	342	326
rect	341	326	342	327
rect	341	327	342	328
rect	341	328	342	329
rect	341	329	342	330
rect	341	330	342	331
rect	341	331	342	332
rect	341	332	342	333
rect	341	333	342	334
rect	341	334	342	335
rect	341	335	342	336
rect	341	336	342	337
rect	341	337	342	338
rect	341	338	342	339
rect	341	339	342	340
rect	341	340	342	341
rect	341	341	342	342
rect	341	342	342	343
rect	341	343	342	344
rect	341	344	342	345
rect	341	345	342	346
rect	341	346	342	347
rect	341	347	342	348
rect	341	348	342	349
rect	341	349	342	350
rect	341	350	342	351
rect	341	351	342	352
rect	341	352	342	353
rect	341	353	342	354
rect	341	354	342	355
rect	341	355	342	356
rect	341	356	342	357
rect	341	357	342	358
rect	341	358	342	359
rect	341	359	342	360
rect	341	360	342	361
rect	341	361	342	362
rect	341	362	342	363
rect	341	363	342	364
rect	341	364	342	365
rect	341	365	342	366
rect	341	366	342	367
rect	341	367	342	368
rect	341	368	342	369
rect	341	369	342	370
rect	341	370	342	371
rect	341	371	342	372
rect	341	372	342	373
rect	341	373	342	374
rect	341	374	342	375
rect	341	375	342	376
rect	341	376	342	377
rect	341	377	342	378
rect	341	378	342	379
rect	341	379	342	380
rect	341	380	342	381
rect	341	381	342	382
rect	341	382	342	383
rect	341	383	342	384
rect	341	384	342	385
rect	341	385	342	386
rect	341	386	342	387
rect	342	0	343	1
rect	342	1	343	2
rect	342	2	343	3
rect	342	3	343	4
rect	342	4	343	5
rect	342	5	343	6
rect	342	6	343	7
rect	342	7	343	8
rect	342	8	343	9
rect	342	9	343	10
rect	342	10	343	11
rect	342	11	343	12
rect	342	12	343	13
rect	342	13	343	14
rect	342	14	343	15
rect	342	15	343	16
rect	342	16	343	17
rect	342	17	343	18
rect	342	18	343	19
rect	342	19	343	20
rect	342	20	343	21
rect	342	21	343	22
rect	342	22	343	23
rect	342	23	343	24
rect	342	24	343	25
rect	342	25	343	26
rect	342	26	343	27
rect	342	27	343	28
rect	342	28	343	29
rect	342	29	343	30
rect	342	30	343	31
rect	342	31	343	32
rect	342	32	343	33
rect	342	33	343	34
rect	342	34	343	35
rect	342	35	343	36
rect	342	36	343	37
rect	342	37	343	38
rect	342	38	343	39
rect	342	39	343	40
rect	342	40	343	41
rect	342	41	343	42
rect	342	42	343	43
rect	342	43	343	44
rect	342	44	343	45
rect	342	45	343	46
rect	342	46	343	47
rect	342	47	343	48
rect	342	48	343	49
rect	342	49	343	50
rect	342	50	343	51
rect	342	51	343	52
rect	342	52	343	53
rect	342	53	343	54
rect	342	54	343	55
rect	342	55	343	56
rect	342	56	343	57
rect	342	57	343	58
rect	342	58	343	59
rect	342	59	343	60
rect	342	60	343	61
rect	342	61	343	62
rect	342	62	343	63
rect	342	63	343	64
rect	342	64	343	65
rect	342	65	343	66
rect	342	66	343	67
rect	342	67	343	68
rect	342	68	343	69
rect	342	69	343	70
rect	342	70	343	71
rect	342	71	343	72
rect	342	72	343	73
rect	342	73	343	74
rect	342	74	343	75
rect	342	75	343	76
rect	342	76	343	77
rect	342	77	343	78
rect	342	78	343	79
rect	342	79	343	80
rect	342	80	343	81
rect	342	81	343	82
rect	342	82	343	83
rect	342	83	343	84
rect	342	84	343	85
rect	342	85	343	86
rect	342	86	343	87
rect	342	87	343	88
rect	342	88	343	89
rect	342	89	343	90
rect	342	90	343	91
rect	342	91	343	92
rect	342	92	343	93
rect	342	93	343	94
rect	342	94	343	95
rect	342	95	343	96
rect	342	96	343	97
rect	342	97	343	98
rect	342	98	343	99
rect	342	99	343	100
rect	342	100	343	101
rect	342	101	343	102
rect	342	102	343	103
rect	342	103	343	104
rect	342	104	343	105
rect	342	105	343	106
rect	342	106	343	107
rect	342	107	343	108
rect	342	108	343	109
rect	342	109	343	110
rect	342	110	343	111
rect	342	111	343	112
rect	342	112	343	113
rect	342	113	343	114
rect	342	114	343	115
rect	342	115	343	116
rect	342	116	343	117
rect	342	117	343	118
rect	342	118	343	119
rect	342	119	343	120
rect	342	120	343	121
rect	342	121	343	122
rect	342	122	343	123
rect	342	123	343	124
rect	342	124	343	125
rect	342	125	343	126
rect	342	126	343	127
rect	342	127	343	128
rect	342	128	343	129
rect	342	129	343	130
rect	342	130	343	131
rect	342	131	343	132
rect	342	132	343	133
rect	342	133	343	134
rect	342	134	343	135
rect	342	135	343	136
rect	342	136	343	137
rect	342	137	343	138
rect	342	138	343	139
rect	342	139	343	140
rect	342	140	343	141
rect	342	141	343	142
rect	342	142	343	143
rect	342	143	343	144
rect	342	144	343	145
rect	342	145	343	146
rect	342	146	343	147
rect	342	147	343	148
rect	342	148	343	149
rect	342	149	343	150
rect	342	150	343	151
rect	342	151	343	152
rect	342	152	343	153
rect	342	153	343	154
rect	342	154	343	155
rect	342	155	343	156
rect	342	156	343	157
rect	342	157	343	158
rect	342	158	343	159
rect	342	159	343	160
rect	342	160	343	161
rect	342	161	343	162
rect	342	162	343	163
rect	342	163	343	164
rect	342	164	343	165
rect	342	165	343	166
rect	342	166	343	167
rect	342	167	343	168
rect	342	168	343	169
rect	342	169	343	170
rect	342	170	343	171
rect	342	171	343	172
rect	342	172	343	173
rect	342	173	343	174
rect	342	174	343	175
rect	342	175	343	176
rect	342	176	343	177
rect	342	177	343	178
rect	342	178	343	179
rect	342	179	343	180
rect	342	180	343	181
rect	342	181	343	182
rect	342	182	343	183
rect	342	183	343	184
rect	342	184	343	185
rect	342	185	343	186
rect	342	186	343	187
rect	342	187	343	188
rect	342	188	343	189
rect	342	189	343	190
rect	342	190	343	191
rect	342	191	343	192
rect	342	192	343	193
rect	342	193	343	194
rect	342	194	343	195
rect	342	195	343	196
rect	342	196	343	197
rect	342	197	343	198
rect	342	198	343	199
rect	342	199	343	200
rect	342	200	343	201
rect	342	201	343	202
rect	342	202	343	203
rect	342	203	343	204
rect	342	204	343	205
rect	342	205	343	206
rect	342	206	343	207
rect	342	207	343	208
rect	342	208	343	209
rect	342	209	343	210
rect	342	210	343	211
rect	342	211	343	212
rect	342	212	343	213
rect	342	213	343	214
rect	342	214	343	215
rect	342	215	343	216
rect	342	216	343	217
rect	342	217	343	218
rect	342	218	343	219
rect	342	219	343	220
rect	342	220	343	221
rect	342	221	343	222
rect	342	222	343	223
rect	342	223	343	224
rect	342	224	343	225
rect	342	225	343	226
rect	342	226	343	227
rect	342	227	343	228
rect	342	228	343	229
rect	342	229	343	230
rect	342	230	343	231
rect	342	231	343	232
rect	342	232	343	233
rect	342	233	343	234
rect	342	234	343	235
rect	342	235	343	236
rect	342	236	343	237
rect	342	237	343	238
rect	342	238	343	239
rect	342	239	343	240
rect	342	240	343	241
rect	342	241	343	242
rect	342	242	343	243
rect	342	243	343	244
rect	342	244	343	245
rect	342	245	343	246
rect	342	246	343	247
rect	342	247	343	248
rect	342	248	343	249
rect	342	249	343	250
rect	342	250	343	251
rect	342	251	343	252
rect	342	252	343	253
rect	342	253	343	254
rect	342	254	343	255
rect	342	255	343	256
rect	342	256	343	257
rect	342	257	343	258
rect	342	258	343	259
rect	342	259	343	260
rect	342	260	343	261
rect	342	261	343	262
rect	342	262	343	263
rect	342	263	343	264
rect	342	264	343	265
rect	342	265	343	266
rect	342	266	343	267
rect	342	267	343	268
rect	342	268	343	269
rect	342	269	343	270
rect	342	270	343	271
rect	342	271	343	272
rect	342	272	343	273
rect	342	273	343	274
rect	342	274	343	275
rect	342	275	343	276
rect	342	276	343	277
rect	342	277	343	278
rect	342	278	343	279
rect	342	279	343	280
rect	342	280	343	281
rect	342	281	343	282
rect	342	282	343	283
rect	342	283	343	284
rect	342	284	343	285
rect	342	285	343	286
rect	342	286	343	287
rect	342	287	343	288
rect	342	288	343	289
rect	342	289	343	290
rect	342	290	343	291
rect	342	291	343	292
rect	342	292	343	293
rect	342	293	343	294
rect	342	294	343	295
rect	342	295	343	296
rect	342	296	343	297
rect	342	297	343	298
rect	342	298	343	299
rect	342	299	343	300
rect	342	300	343	301
rect	342	301	343	302
rect	342	302	343	303
rect	342	303	343	304
rect	342	304	343	305
rect	342	305	343	306
rect	342	306	343	307
rect	342	307	343	308
rect	342	308	343	309
rect	342	309	343	310
rect	342	310	343	311
rect	342	311	343	312
rect	342	312	343	313
rect	342	313	343	314
rect	342	314	343	315
rect	342	315	343	316
rect	342	316	343	317
rect	342	317	343	318
rect	342	318	343	319
rect	342	319	343	320
rect	342	320	343	321
rect	342	321	343	322
rect	342	322	343	323
rect	342	323	343	324
rect	342	324	343	325
rect	342	325	343	326
rect	342	326	343	327
rect	342	327	343	328
rect	342	328	343	329
rect	342	329	343	330
rect	342	330	343	331
rect	342	331	343	332
rect	342	332	343	333
rect	342	333	343	334
rect	342	334	343	335
rect	342	335	343	336
rect	342	336	343	337
rect	342	337	343	338
rect	342	338	343	339
rect	342	339	343	340
rect	342	340	343	341
rect	342	341	343	342
rect	342	342	343	343
rect	342	343	343	344
rect	342	344	343	345
rect	342	345	343	346
rect	342	346	343	347
rect	342	347	343	348
rect	342	348	343	349
rect	342	349	343	350
rect	342	350	343	351
rect	342	351	343	352
rect	342	352	343	353
rect	342	353	343	354
rect	342	354	343	355
rect	342	355	343	356
rect	342	356	343	357
rect	342	357	343	358
rect	342	358	343	359
rect	342	359	343	360
rect	342	360	343	361
rect	342	361	343	362
rect	342	362	343	363
rect	342	363	343	364
rect	342	364	343	365
rect	342	365	343	366
rect	342	366	343	367
rect	342	367	343	368
rect	342	368	343	369
rect	342	369	343	370
rect	342	370	343	371
rect	342	371	343	372
rect	342	372	343	373
rect	342	373	343	374
rect	342	374	343	375
rect	342	375	343	376
rect	342	376	343	377
rect	342	377	343	378
rect	342	378	343	379
rect	342	379	343	380
rect	342	380	343	381
rect	342	381	343	382
rect	342	382	343	383
rect	342	383	343	384
rect	342	384	343	385
rect	342	385	343	386
rect	342	386	343	387
rect	370	0	371	1
rect	370	1	371	2
rect	370	2	371	3
rect	370	3	371	4
rect	370	4	371	5
rect	370	5	371	6
rect	370	6	371	7
rect	370	7	371	8
rect	370	8	371	9
rect	370	9	371	10
rect	370	10	371	11
rect	370	11	371	12
rect	370	12	371	13
rect	370	13	371	14
rect	370	14	371	15
rect	370	15	371	16
rect	370	16	371	17
rect	370	17	371	18
rect	370	18	371	19
rect	370	19	371	20
rect	370	20	371	21
rect	370	21	371	22
rect	370	22	371	23
rect	370	23	371	24
rect	370	24	371	25
rect	370	25	371	26
rect	370	26	371	27
rect	370	27	371	28
rect	370	28	371	29
rect	370	29	371	30
rect	370	30	371	31
rect	370	31	371	32
rect	370	32	371	33
rect	370	33	371	34
rect	370	34	371	35
rect	370	35	371	36
rect	370	36	371	37
rect	370	37	371	38
rect	370	38	371	39
rect	370	39	371	40
rect	370	40	371	41
rect	370	41	371	42
rect	370	42	371	43
rect	370	43	371	44
rect	370	44	371	45
rect	370	45	371	46
rect	370	46	371	47
rect	370	47	371	48
rect	370	48	371	49
rect	370	49	371	50
rect	370	50	371	51
rect	370	51	371	52
rect	370	52	371	53
rect	370	53	371	54
rect	370	54	371	55
rect	370	55	371	56
rect	370	56	371	57
rect	370	57	371	58
rect	370	58	371	59
rect	370	59	371	60
rect	370	60	371	61
rect	370	61	371	62
rect	370	62	371	63
rect	370	63	371	64
rect	370	64	371	65
rect	370	65	371	66
rect	370	66	371	67
rect	370	67	371	68
rect	370	68	371	69
rect	370	69	371	70
rect	370	70	371	71
rect	370	71	371	72
rect	370	72	371	73
rect	370	73	371	74
rect	370	74	371	75
rect	370	75	371	76
rect	370	76	371	77
rect	370	77	371	78
rect	370	78	371	79
rect	370	79	371	80
rect	370	80	371	81
rect	370	81	371	82
rect	370	82	371	83
rect	370	83	371	84
rect	370	84	371	85
rect	370	85	371	86
rect	370	86	371	87
rect	370	87	371	88
rect	370	88	371	89
rect	370	89	371	90
rect	370	90	371	91
rect	370	91	371	92
rect	370	92	371	93
rect	370	93	371	94
rect	370	94	371	95
rect	370	95	371	96
rect	370	96	371	97
rect	370	97	371	98
rect	370	98	371	99
rect	370	99	371	100
rect	370	100	371	101
rect	370	101	371	102
rect	370	102	371	103
rect	370	103	371	104
rect	370	104	371	105
rect	370	105	371	106
rect	370	106	371	107
rect	370	107	371	108
rect	370	108	371	109
rect	370	109	371	110
rect	370	110	371	111
rect	370	111	371	112
rect	370	112	371	113
rect	370	113	371	114
rect	370	114	371	115
rect	370	115	371	116
rect	370	116	371	117
rect	370	117	371	118
rect	370	118	371	119
rect	370	119	371	120
rect	370	120	371	121
rect	370	121	371	122
rect	370	122	371	123
rect	370	123	371	124
rect	370	124	371	125
rect	370	125	371	126
rect	370	126	371	127
rect	370	127	371	128
rect	370	128	371	129
rect	370	129	371	130
rect	370	130	371	131
rect	370	131	371	132
rect	370	132	371	133
rect	370	133	371	134
rect	370	134	371	135
rect	370	135	371	136
rect	370	136	371	137
rect	370	137	371	138
rect	370	138	371	139
rect	370	139	371	140
rect	370	140	371	141
rect	370	141	371	142
rect	370	142	371	143
rect	370	143	371	144
rect	370	144	371	145
rect	370	145	371	146
rect	370	146	371	147
rect	370	147	371	148
rect	370	148	371	149
rect	370	149	371	150
rect	370	150	371	151
rect	370	151	371	152
rect	370	152	371	153
rect	370	153	371	154
rect	370	154	371	155
rect	370	155	371	156
rect	370	156	371	157
rect	370	157	371	158
rect	370	158	371	159
rect	370	159	371	160
rect	370	160	371	161
rect	370	161	371	162
rect	370	162	371	163
rect	370	163	371	164
rect	370	164	371	165
rect	370	165	371	166
rect	370	166	371	167
rect	370	167	371	168
rect	370	168	371	169
rect	370	169	371	170
rect	370	170	371	171
rect	370	171	371	172
rect	370	172	371	173
rect	370	173	371	174
rect	370	174	371	175
rect	370	175	371	176
rect	370	176	371	177
rect	370	177	371	178
rect	370	178	371	179
rect	370	179	371	180
rect	370	180	371	181
rect	370	181	371	182
rect	370	182	371	183
rect	370	183	371	184
rect	370	184	371	185
rect	370	185	371	186
rect	370	186	371	187
rect	370	187	371	188
rect	370	188	371	189
rect	370	189	371	190
rect	370	190	371	191
rect	370	191	371	192
rect	370	192	371	193
rect	370	193	371	194
rect	370	194	371	195
rect	370	195	371	196
rect	370	196	371	197
rect	370	197	371	198
rect	370	198	371	199
rect	370	199	371	200
rect	370	200	371	201
rect	370	201	371	202
rect	370	202	371	203
rect	370	203	371	204
rect	370	204	371	205
rect	370	205	371	206
rect	370	206	371	207
rect	370	207	371	208
rect	370	208	371	209
rect	370	209	371	210
rect	370	210	371	211
rect	370	211	371	212
rect	370	212	371	213
rect	370	213	371	214
rect	370	214	371	215
rect	370	215	371	216
rect	370	216	371	217
rect	370	217	371	218
rect	370	218	371	219
rect	370	219	371	220
rect	370	220	371	221
rect	370	221	371	222
rect	370	222	371	223
rect	370	223	371	224
rect	370	224	371	225
rect	370	225	371	226
rect	370	226	371	227
rect	370	227	371	228
rect	370	228	371	229
rect	370	229	371	230
rect	370	230	371	231
rect	370	231	371	232
rect	370	232	371	233
rect	370	233	371	234
rect	370	234	371	235
rect	370	235	371	236
rect	370	236	371	237
rect	370	237	371	238
rect	370	238	371	239
rect	370	239	371	240
rect	370	240	371	241
rect	370	241	371	242
rect	370	242	371	243
rect	370	243	371	244
rect	370	244	371	245
rect	370	245	371	246
rect	370	246	371	247
rect	370	247	371	248
rect	370	248	371	249
rect	370	249	371	250
rect	370	250	371	251
rect	370	251	371	252
rect	370	252	371	253
rect	370	253	371	254
rect	370	254	371	255
rect	370	255	371	256
rect	370	256	371	257
rect	370	257	371	258
rect	370	258	371	259
rect	370	259	371	260
rect	370	260	371	261
rect	370	261	371	262
rect	370	262	371	263
rect	370	263	371	264
rect	370	264	371	265
rect	370	265	371	266
rect	370	266	371	267
rect	370	267	371	268
rect	370	268	371	269
rect	370	269	371	270
rect	370	270	371	271
rect	370	271	371	272
rect	370	272	371	273
rect	370	273	371	274
rect	370	274	371	275
rect	370	275	371	276
rect	370	276	371	277
rect	370	277	371	278
rect	370	278	371	279
rect	370	279	371	280
rect	370	280	371	281
rect	370	281	371	282
rect	370	282	371	283
rect	370	283	371	284
rect	370	284	371	285
rect	370	285	371	286
rect	370	286	371	287
rect	370	287	371	288
rect	370	288	371	289
rect	370	289	371	290
rect	370	290	371	291
rect	370	291	371	292
rect	370	292	371	293
rect	370	293	371	294
rect	370	294	371	295
rect	370	295	371	296
rect	370	296	371	297
rect	370	297	371	298
rect	370	298	371	299
rect	370	299	371	300
rect	370	300	371	301
rect	370	301	371	302
rect	370	302	371	303
rect	370	303	371	304
rect	370	304	371	305
rect	370	305	371	306
rect	370	306	371	307
rect	370	307	371	308
rect	370	308	371	309
rect	370	309	371	310
rect	370	310	371	311
rect	370	311	371	312
rect	370	312	371	313
rect	370	313	371	314
rect	370	314	371	315
rect	370	315	371	316
rect	370	316	371	317
rect	370	317	371	318
rect	370	318	371	319
rect	370	319	371	320
rect	370	320	371	321
rect	370	321	371	322
rect	370	322	371	323
rect	370	323	371	324
rect	370	324	371	325
rect	370	325	371	326
rect	370	326	371	327
rect	370	327	371	328
rect	370	328	371	329
rect	370	329	371	330
rect	370	330	371	331
rect	370	331	371	332
rect	370	332	371	333
rect	370	333	371	334
rect	370	334	371	335
rect	370	335	371	336
rect	370	336	371	337
rect	370	337	371	338
rect	370	338	371	339
rect	370	339	371	340
rect	370	340	371	341
rect	370	341	371	342
rect	370	342	371	343
rect	370	343	371	344
rect	370	344	371	345
rect	370	345	371	346
rect	370	346	371	347
rect	370	347	371	348
rect	370	348	371	349
rect	370	349	371	350
rect	370	350	371	351
rect	370	351	371	352
rect	370	352	371	353
rect	370	353	371	354
rect	370	354	371	355
rect	370	355	371	356
rect	370	356	371	357
rect	370	357	371	358
rect	370	358	371	359
rect	370	359	371	360
rect	370	360	371	361
rect	370	361	371	362
rect	370	362	371	363
rect	370	363	371	364
rect	370	364	371	365
rect	370	365	371	366
rect	370	366	371	367
rect	370	367	371	368
rect	370	368	371	369
rect	371	0	372	1
rect	371	1	372	2
rect	371	2	372	3
rect	371	3	372	4
rect	371	4	372	5
rect	371	5	372	6
rect	371	6	372	7
rect	371	7	372	8
rect	371	8	372	9
rect	371	9	372	10
rect	371	10	372	11
rect	371	11	372	12
rect	371	12	372	13
rect	371	13	372	14
rect	371	14	372	15
rect	371	15	372	16
rect	371	16	372	17
rect	371	17	372	18
rect	371	18	372	19
rect	371	19	372	20
rect	371	20	372	21
rect	371	21	372	22
rect	371	22	372	23
rect	371	23	372	24
rect	371	24	372	25
rect	371	25	372	26
rect	371	26	372	27
rect	371	27	372	28
rect	371	28	372	29
rect	371	29	372	30
rect	371	30	372	31
rect	371	31	372	32
rect	371	32	372	33
rect	371	33	372	34
rect	371	34	372	35
rect	371	35	372	36
rect	371	36	372	37
rect	371	37	372	38
rect	371	38	372	39
rect	371	39	372	40
rect	371	40	372	41
rect	371	41	372	42
rect	371	42	372	43
rect	371	43	372	44
rect	371	44	372	45
rect	371	45	372	46
rect	371	46	372	47
rect	371	47	372	48
rect	371	48	372	49
rect	371	49	372	50
rect	371	50	372	51
rect	371	51	372	52
rect	371	52	372	53
rect	371	53	372	54
rect	371	54	372	55
rect	371	55	372	56
rect	371	56	372	57
rect	371	57	372	58
rect	371	58	372	59
rect	371	59	372	60
rect	371	60	372	61
rect	371	61	372	62
rect	371	62	372	63
rect	371	63	372	64
rect	371	64	372	65
rect	371	65	372	66
rect	371	66	372	67
rect	371	67	372	68
rect	371	68	372	69
rect	371	69	372	70
rect	371	70	372	71
rect	371	71	372	72
rect	371	72	372	73
rect	371	73	372	74
rect	371	74	372	75
rect	371	75	372	76
rect	371	76	372	77
rect	371	77	372	78
rect	371	78	372	79
rect	371	79	372	80
rect	371	80	372	81
rect	371	81	372	82
rect	371	82	372	83
rect	371	83	372	84
rect	371	84	372	85
rect	371	85	372	86
rect	371	86	372	87
rect	371	87	372	88
rect	371	88	372	89
rect	371	89	372	90
rect	371	90	372	91
rect	371	91	372	92
rect	371	92	372	93
rect	371	93	372	94
rect	371	94	372	95
rect	371	95	372	96
rect	371	96	372	97
rect	371	97	372	98
rect	371	98	372	99
rect	371	99	372	100
rect	371	100	372	101
rect	371	101	372	102
rect	371	102	372	103
rect	371	103	372	104
rect	371	104	372	105
rect	371	105	372	106
rect	371	106	372	107
rect	371	107	372	108
rect	371	108	372	109
rect	371	109	372	110
rect	371	110	372	111
rect	371	111	372	112
rect	371	112	372	113
rect	371	113	372	114
rect	371	114	372	115
rect	371	115	372	116
rect	371	116	372	117
rect	371	117	372	118
rect	371	118	372	119
rect	371	119	372	120
rect	371	120	372	121
rect	371	121	372	122
rect	371	122	372	123
rect	371	123	372	124
rect	371	124	372	125
rect	371	125	372	126
rect	371	126	372	127
rect	371	127	372	128
rect	371	128	372	129
rect	371	129	372	130
rect	371	130	372	131
rect	371	131	372	132
rect	371	132	372	133
rect	371	133	372	134
rect	371	134	372	135
rect	371	135	372	136
rect	371	136	372	137
rect	371	137	372	138
rect	371	138	372	139
rect	371	139	372	140
rect	371	140	372	141
rect	371	141	372	142
rect	371	142	372	143
rect	371	143	372	144
rect	371	144	372	145
rect	371	145	372	146
rect	371	146	372	147
rect	371	147	372	148
rect	371	148	372	149
rect	371	149	372	150
rect	371	150	372	151
rect	371	151	372	152
rect	371	152	372	153
rect	371	153	372	154
rect	371	154	372	155
rect	371	155	372	156
rect	371	156	372	157
rect	371	157	372	158
rect	371	158	372	159
rect	371	159	372	160
rect	371	160	372	161
rect	371	161	372	162
rect	371	162	372	163
rect	371	163	372	164
rect	371	164	372	165
rect	371	165	372	166
rect	371	166	372	167
rect	371	167	372	168
rect	371	168	372	169
rect	371	169	372	170
rect	371	170	372	171
rect	371	171	372	172
rect	371	172	372	173
rect	371	173	372	174
rect	371	174	372	175
rect	371	175	372	176
rect	371	176	372	177
rect	371	177	372	178
rect	371	178	372	179
rect	371	179	372	180
rect	371	180	372	181
rect	371	181	372	182
rect	371	182	372	183
rect	371	183	372	184
rect	371	184	372	185
rect	371	185	372	186
rect	371	186	372	187
rect	371	187	372	188
rect	371	188	372	189
rect	371	189	372	190
rect	371	190	372	191
rect	371	191	372	192
rect	371	192	372	193
rect	371	193	372	194
rect	371	194	372	195
rect	371	195	372	196
rect	371	196	372	197
rect	371	197	372	198
rect	371	198	372	199
rect	371	199	372	200
rect	371	200	372	201
rect	371	201	372	202
rect	371	202	372	203
rect	371	203	372	204
rect	371	204	372	205
rect	371	205	372	206
rect	371	206	372	207
rect	371	207	372	208
rect	371	208	372	209
rect	371	209	372	210
rect	371	210	372	211
rect	371	211	372	212
rect	371	212	372	213
rect	371	213	372	214
rect	371	214	372	215
rect	371	215	372	216
rect	371	216	372	217
rect	371	217	372	218
rect	371	218	372	219
rect	371	219	372	220
rect	371	220	372	221
rect	371	221	372	222
rect	371	222	372	223
rect	371	223	372	224
rect	371	224	372	225
rect	371	225	372	226
rect	371	226	372	227
rect	371	227	372	228
rect	371	228	372	229
rect	371	229	372	230
rect	371	230	372	231
rect	371	231	372	232
rect	371	232	372	233
rect	371	233	372	234
rect	371	234	372	235
rect	371	235	372	236
rect	371	236	372	237
rect	371	237	372	238
rect	371	238	372	239
rect	371	239	372	240
rect	371	240	372	241
rect	371	241	372	242
rect	371	242	372	243
rect	371	243	372	244
rect	371	244	372	245
rect	371	245	372	246
rect	371	246	372	247
rect	371	247	372	248
rect	371	248	372	249
rect	371	249	372	250
rect	371	250	372	251
rect	371	251	372	252
rect	371	252	372	253
rect	371	253	372	254
rect	371	254	372	255
rect	371	255	372	256
rect	371	256	372	257
rect	371	257	372	258
rect	371	258	372	259
rect	371	259	372	260
rect	371	260	372	261
rect	371	261	372	262
rect	371	262	372	263
rect	371	263	372	264
rect	371	264	372	265
rect	371	265	372	266
rect	371	266	372	267
rect	371	267	372	268
rect	371	268	372	269
rect	371	269	372	270
rect	371	270	372	271
rect	371	271	372	272
rect	371	272	372	273
rect	371	273	372	274
rect	371	274	372	275
rect	371	275	372	276
rect	371	276	372	277
rect	371	277	372	278
rect	371	278	372	279
rect	371	279	372	280
rect	371	280	372	281
rect	371	281	372	282
rect	371	282	372	283
rect	371	283	372	284
rect	371	284	372	285
rect	371	285	372	286
rect	371	286	372	287
rect	371	287	372	288
rect	371	288	372	289
rect	371	289	372	290
rect	371	290	372	291
rect	371	291	372	292
rect	371	292	372	293
rect	371	293	372	294
rect	371	294	372	295
rect	371	295	372	296
rect	371	296	372	297
rect	371	297	372	298
rect	371	298	372	299
rect	371	299	372	300
rect	371	300	372	301
rect	371	301	372	302
rect	371	302	372	303
rect	371	303	372	304
rect	371	304	372	305
rect	371	305	372	306
rect	371	306	372	307
rect	371	307	372	308
rect	371	308	372	309
rect	371	309	372	310
rect	371	310	372	311
rect	371	311	372	312
rect	371	312	372	313
rect	371	313	372	314
rect	371	314	372	315
rect	371	315	372	316
rect	371	316	372	317
rect	371	317	372	318
rect	371	318	372	319
rect	371	319	372	320
rect	371	320	372	321
rect	371	321	372	322
rect	371	322	372	323
rect	371	323	372	324
rect	371	324	372	325
rect	371	325	372	326
rect	371	326	372	327
rect	371	327	372	328
rect	371	328	372	329
rect	371	329	372	330
rect	371	330	372	331
rect	371	331	372	332
rect	371	332	372	333
rect	371	333	372	334
rect	371	334	372	335
rect	371	335	372	336
rect	371	336	372	337
rect	371	337	372	338
rect	371	338	372	339
rect	371	339	372	340
rect	371	340	372	341
rect	371	341	372	342
rect	371	342	372	343
rect	371	343	372	344
rect	371	344	372	345
rect	371	345	372	346
rect	371	346	372	347
rect	371	347	372	348
rect	371	348	372	349
rect	371	349	372	350
rect	371	350	372	351
rect	371	351	372	352
rect	371	352	372	353
rect	371	353	372	354
rect	371	354	372	355
rect	371	355	372	356
rect	371	356	372	357
rect	371	357	372	358
rect	371	358	372	359
rect	371	359	372	360
rect	371	360	372	361
rect	371	361	372	362
rect	371	362	372	363
rect	371	363	372	364
rect	371	364	372	365
rect	371	365	372	366
rect	371	366	372	367
rect	371	367	372	368
rect	371	368	372	369
rect	372	0	373	1
rect	372	1	373	2
rect	372	2	373	3
rect	372	3	373	4
rect	372	4	373	5
rect	372	5	373	6
rect	372	6	373	7
rect	372	7	373	8
rect	372	8	373	9
rect	372	9	373	10
rect	372	10	373	11
rect	372	11	373	12
rect	372	12	373	13
rect	372	13	373	14
rect	372	14	373	15
rect	372	15	373	16
rect	372	16	373	17
rect	372	17	373	18
rect	372	18	373	19
rect	372	19	373	20
rect	372	20	373	21
rect	372	21	373	22
rect	372	22	373	23
rect	372	23	373	24
rect	372	24	373	25
rect	372	25	373	26
rect	372	26	373	27
rect	372	27	373	28
rect	372	28	373	29
rect	372	29	373	30
rect	372	30	373	31
rect	372	31	373	32
rect	372	32	373	33
rect	372	33	373	34
rect	372	34	373	35
rect	372	35	373	36
rect	372	36	373	37
rect	372	37	373	38
rect	372	38	373	39
rect	372	39	373	40
rect	372	40	373	41
rect	372	41	373	42
rect	372	42	373	43
rect	372	43	373	44
rect	372	44	373	45
rect	372	45	373	46
rect	372	46	373	47
rect	372	47	373	48
rect	372	48	373	49
rect	372	49	373	50
rect	372	50	373	51
rect	372	51	373	52
rect	372	52	373	53
rect	372	53	373	54
rect	372	54	373	55
rect	372	55	373	56
rect	372	56	373	57
rect	372	57	373	58
rect	372	58	373	59
rect	372	59	373	60
rect	372	60	373	61
rect	372	61	373	62
rect	372	62	373	63
rect	372	63	373	64
rect	372	64	373	65
rect	372	65	373	66
rect	372	66	373	67
rect	372	67	373	68
rect	372	68	373	69
rect	372	69	373	70
rect	372	70	373	71
rect	372	71	373	72
rect	372	72	373	73
rect	372	73	373	74
rect	372	74	373	75
rect	372	75	373	76
rect	372	76	373	77
rect	372	77	373	78
rect	372	78	373	79
rect	372	79	373	80
rect	372	80	373	81
rect	372	81	373	82
rect	372	82	373	83
rect	372	83	373	84
rect	372	84	373	85
rect	372	85	373	86
rect	372	86	373	87
rect	372	87	373	88
rect	372	88	373	89
rect	372	89	373	90
rect	372	90	373	91
rect	372	91	373	92
rect	372	92	373	93
rect	372	93	373	94
rect	372	94	373	95
rect	372	95	373	96
rect	372	96	373	97
rect	372	97	373	98
rect	372	98	373	99
rect	372	99	373	100
rect	372	100	373	101
rect	372	101	373	102
rect	372	102	373	103
rect	372	103	373	104
rect	372	104	373	105
rect	372	105	373	106
rect	372	106	373	107
rect	372	107	373	108
rect	372	108	373	109
rect	372	109	373	110
rect	372	110	373	111
rect	372	111	373	112
rect	372	112	373	113
rect	372	113	373	114
rect	372	114	373	115
rect	372	115	373	116
rect	372	116	373	117
rect	372	117	373	118
rect	372	118	373	119
rect	372	119	373	120
rect	372	120	373	121
rect	372	121	373	122
rect	372	122	373	123
rect	372	123	373	124
rect	372	124	373	125
rect	372	125	373	126
rect	372	126	373	127
rect	372	127	373	128
rect	372	128	373	129
rect	372	129	373	130
rect	372	130	373	131
rect	372	131	373	132
rect	372	132	373	133
rect	372	133	373	134
rect	372	134	373	135
rect	372	135	373	136
rect	372	136	373	137
rect	372	137	373	138
rect	372	138	373	139
rect	372	139	373	140
rect	372	140	373	141
rect	372	141	373	142
rect	372	142	373	143
rect	372	143	373	144
rect	372	144	373	145
rect	372	145	373	146
rect	372	146	373	147
rect	372	147	373	148
rect	372	148	373	149
rect	372	149	373	150
rect	372	150	373	151
rect	372	151	373	152
rect	372	152	373	153
rect	372	153	373	154
rect	372	154	373	155
rect	372	155	373	156
rect	372	156	373	157
rect	372	157	373	158
rect	372	158	373	159
rect	372	159	373	160
rect	372	160	373	161
rect	372	161	373	162
rect	372	162	373	163
rect	372	163	373	164
rect	372	164	373	165
rect	372	165	373	166
rect	372	166	373	167
rect	372	167	373	168
rect	372	168	373	169
rect	372	169	373	170
rect	372	170	373	171
rect	372	171	373	172
rect	372	172	373	173
rect	372	173	373	174
rect	372	174	373	175
rect	372	175	373	176
rect	372	176	373	177
rect	372	177	373	178
rect	372	178	373	179
rect	372	179	373	180
rect	372	180	373	181
rect	372	181	373	182
rect	372	182	373	183
rect	372	183	373	184
rect	372	184	373	185
rect	372	185	373	186
rect	372	186	373	187
rect	372	187	373	188
rect	372	188	373	189
rect	372	189	373	190
rect	372	190	373	191
rect	372	191	373	192
rect	372	192	373	193
rect	372	193	373	194
rect	372	194	373	195
rect	372	195	373	196
rect	372	196	373	197
rect	372	197	373	198
rect	372	198	373	199
rect	372	199	373	200
rect	372	200	373	201
rect	372	201	373	202
rect	372	202	373	203
rect	372	203	373	204
rect	372	204	373	205
rect	372	205	373	206
rect	372	206	373	207
rect	372	207	373	208
rect	372	208	373	209
rect	372	209	373	210
rect	372	210	373	211
rect	372	211	373	212
rect	372	212	373	213
rect	372	213	373	214
rect	372	214	373	215
rect	372	215	373	216
rect	372	216	373	217
rect	372	217	373	218
rect	372	218	373	219
rect	372	219	373	220
rect	372	220	373	221
rect	372	221	373	222
rect	372	222	373	223
rect	372	223	373	224
rect	372	224	373	225
rect	372	225	373	226
rect	372	226	373	227
rect	372	227	373	228
rect	372	228	373	229
rect	372	229	373	230
rect	372	230	373	231
rect	372	231	373	232
rect	372	232	373	233
rect	372	233	373	234
rect	372	234	373	235
rect	372	235	373	236
rect	372	236	373	237
rect	372	237	373	238
rect	372	238	373	239
rect	372	239	373	240
rect	372	240	373	241
rect	372	241	373	242
rect	372	242	373	243
rect	372	243	373	244
rect	372	244	373	245
rect	372	245	373	246
rect	372	246	373	247
rect	372	247	373	248
rect	372	248	373	249
rect	372	249	373	250
rect	372	250	373	251
rect	372	251	373	252
rect	372	252	373	253
rect	372	253	373	254
rect	372	254	373	255
rect	372	255	373	256
rect	372	256	373	257
rect	372	257	373	258
rect	372	258	373	259
rect	372	259	373	260
rect	372	260	373	261
rect	372	261	373	262
rect	372	262	373	263
rect	372	263	373	264
rect	372	264	373	265
rect	372	265	373	266
rect	372	266	373	267
rect	372	267	373	268
rect	372	268	373	269
rect	372	269	373	270
rect	372	270	373	271
rect	372	271	373	272
rect	372	272	373	273
rect	372	273	373	274
rect	372	274	373	275
rect	372	275	373	276
rect	372	276	373	277
rect	372	277	373	278
rect	372	278	373	279
rect	372	279	373	280
rect	372	280	373	281
rect	372	281	373	282
rect	372	282	373	283
rect	372	283	373	284
rect	372	284	373	285
rect	372	285	373	286
rect	372	286	373	287
rect	372	287	373	288
rect	372	288	373	289
rect	372	289	373	290
rect	372	290	373	291
rect	372	291	373	292
rect	372	292	373	293
rect	372	293	373	294
rect	372	294	373	295
rect	372	295	373	296
rect	372	296	373	297
rect	372	297	373	298
rect	372	298	373	299
rect	372	299	373	300
rect	372	300	373	301
rect	372	301	373	302
rect	372	302	373	303
rect	372	303	373	304
rect	372	304	373	305
rect	372	305	373	306
rect	372	306	373	307
rect	372	307	373	308
rect	372	308	373	309
rect	372	309	373	310
rect	372	310	373	311
rect	372	311	373	312
rect	372	312	373	313
rect	372	313	373	314
rect	372	314	373	315
rect	372	315	373	316
rect	372	316	373	317
rect	372	317	373	318
rect	372	318	373	319
rect	372	319	373	320
rect	372	320	373	321
rect	372	321	373	322
rect	372	322	373	323
rect	372	323	373	324
rect	372	324	373	325
rect	372	325	373	326
rect	372	326	373	327
rect	372	327	373	328
rect	372	328	373	329
rect	372	329	373	330
rect	372	330	373	331
rect	372	331	373	332
rect	372	332	373	333
rect	372	333	373	334
rect	372	334	373	335
rect	372	335	373	336
rect	372	336	373	337
rect	372	337	373	338
rect	372	338	373	339
rect	372	339	373	340
rect	372	340	373	341
rect	372	341	373	342
rect	372	342	373	343
rect	372	343	373	344
rect	372	344	373	345
rect	372	345	373	346
rect	372	346	373	347
rect	372	347	373	348
rect	372	348	373	349
rect	372	349	373	350
rect	372	350	373	351
rect	372	351	373	352
rect	372	352	373	353
rect	372	353	373	354
rect	372	354	373	355
rect	372	355	373	356
rect	372	356	373	357
rect	372	357	373	358
rect	372	358	373	359
rect	372	359	373	360
rect	372	360	373	361
rect	372	361	373	362
rect	372	362	373	363
rect	372	363	373	364
rect	372	364	373	365
rect	372	365	373	366
rect	372	366	373	367
rect	372	367	373	368
rect	372	368	373	369
rect	373	0	374	1
rect	373	1	374	2
rect	373	2	374	3
rect	373	3	374	4
rect	373	4	374	5
rect	373	5	374	6
rect	373	6	374	7
rect	373	7	374	8
rect	373	8	374	9
rect	373	9	374	10
rect	373	10	374	11
rect	373	11	374	12
rect	373	12	374	13
rect	373	13	374	14
rect	373	14	374	15
rect	373	15	374	16
rect	373	16	374	17
rect	373	17	374	18
rect	373	18	374	19
rect	373	19	374	20
rect	373	20	374	21
rect	373	21	374	22
rect	373	22	374	23
rect	373	23	374	24
rect	373	24	374	25
rect	373	25	374	26
rect	373	26	374	27
rect	373	27	374	28
rect	373	28	374	29
rect	373	29	374	30
rect	373	30	374	31
rect	373	31	374	32
rect	373	32	374	33
rect	373	33	374	34
rect	373	34	374	35
rect	373	35	374	36
rect	373	36	374	37
rect	373	37	374	38
rect	373	38	374	39
rect	373	39	374	40
rect	373	40	374	41
rect	373	41	374	42
rect	373	42	374	43
rect	373	43	374	44
rect	373	44	374	45
rect	373	45	374	46
rect	373	46	374	47
rect	373	47	374	48
rect	373	48	374	49
rect	373	49	374	50
rect	373	50	374	51
rect	373	51	374	52
rect	373	52	374	53
rect	373	53	374	54
rect	373	54	374	55
rect	373	55	374	56
rect	373	56	374	57
rect	373	57	374	58
rect	373	58	374	59
rect	373	59	374	60
rect	373	60	374	61
rect	373	61	374	62
rect	373	62	374	63
rect	373	63	374	64
rect	373	64	374	65
rect	373	65	374	66
rect	373	66	374	67
rect	373	67	374	68
rect	373	68	374	69
rect	373	69	374	70
rect	373	70	374	71
rect	373	71	374	72
rect	373	72	374	73
rect	373	73	374	74
rect	373	74	374	75
rect	373	75	374	76
rect	373	76	374	77
rect	373	77	374	78
rect	373	78	374	79
rect	373	79	374	80
rect	373	80	374	81
rect	373	81	374	82
rect	373	82	374	83
rect	373	83	374	84
rect	373	84	374	85
rect	373	85	374	86
rect	373	86	374	87
rect	373	87	374	88
rect	373	88	374	89
rect	373	89	374	90
rect	373	90	374	91
rect	373	91	374	92
rect	373	92	374	93
rect	373	93	374	94
rect	373	94	374	95
rect	373	95	374	96
rect	373	96	374	97
rect	373	97	374	98
rect	373	98	374	99
rect	373	99	374	100
rect	373	100	374	101
rect	373	101	374	102
rect	373	102	374	103
rect	373	103	374	104
rect	373	104	374	105
rect	373	105	374	106
rect	373	106	374	107
rect	373	107	374	108
rect	373	108	374	109
rect	373	109	374	110
rect	373	110	374	111
rect	373	111	374	112
rect	373	112	374	113
rect	373	113	374	114
rect	373	114	374	115
rect	373	115	374	116
rect	373	116	374	117
rect	373	117	374	118
rect	373	118	374	119
rect	373	119	374	120
rect	373	120	374	121
rect	373	121	374	122
rect	373	122	374	123
rect	373	123	374	124
rect	373	124	374	125
rect	373	125	374	126
rect	373	126	374	127
rect	373	127	374	128
rect	373	128	374	129
rect	373	129	374	130
rect	373	130	374	131
rect	373	131	374	132
rect	373	132	374	133
rect	373	133	374	134
rect	373	134	374	135
rect	373	135	374	136
rect	373	136	374	137
rect	373	137	374	138
rect	373	138	374	139
rect	373	139	374	140
rect	373	140	374	141
rect	373	141	374	142
rect	373	142	374	143
rect	373	143	374	144
rect	373	144	374	145
rect	373	145	374	146
rect	373	146	374	147
rect	373	147	374	148
rect	373	148	374	149
rect	373	149	374	150
rect	373	150	374	151
rect	373	151	374	152
rect	373	152	374	153
rect	373	153	374	154
rect	373	154	374	155
rect	373	155	374	156
rect	373	156	374	157
rect	373	157	374	158
rect	373	158	374	159
rect	373	159	374	160
rect	373	160	374	161
rect	373	161	374	162
rect	373	162	374	163
rect	373	163	374	164
rect	373	164	374	165
rect	373	165	374	166
rect	373	166	374	167
rect	373	167	374	168
rect	373	168	374	169
rect	373	169	374	170
rect	373	170	374	171
rect	373	171	374	172
rect	373	172	374	173
rect	373	173	374	174
rect	373	174	374	175
rect	373	175	374	176
rect	373	176	374	177
rect	373	177	374	178
rect	373	178	374	179
rect	373	179	374	180
rect	373	180	374	181
rect	373	181	374	182
rect	373	182	374	183
rect	373	183	374	184
rect	373	184	374	185
rect	373	185	374	186
rect	373	186	374	187
rect	373	187	374	188
rect	373	188	374	189
rect	373	189	374	190
rect	373	190	374	191
rect	373	191	374	192
rect	373	192	374	193
rect	373	193	374	194
rect	373	194	374	195
rect	373	195	374	196
rect	373	196	374	197
rect	373	197	374	198
rect	373	198	374	199
rect	373	199	374	200
rect	373	200	374	201
rect	373	201	374	202
rect	373	202	374	203
rect	373	203	374	204
rect	373	204	374	205
rect	373	205	374	206
rect	373	206	374	207
rect	373	207	374	208
rect	373	208	374	209
rect	373	209	374	210
rect	373	210	374	211
rect	373	211	374	212
rect	373	212	374	213
rect	373	213	374	214
rect	373	214	374	215
rect	373	215	374	216
rect	373	216	374	217
rect	373	217	374	218
rect	373	218	374	219
rect	373	219	374	220
rect	373	220	374	221
rect	373	221	374	222
rect	373	222	374	223
rect	373	223	374	224
rect	373	224	374	225
rect	373	225	374	226
rect	373	226	374	227
rect	373	227	374	228
rect	373	228	374	229
rect	373	229	374	230
rect	373	230	374	231
rect	373	231	374	232
rect	373	232	374	233
rect	373	233	374	234
rect	373	234	374	235
rect	373	235	374	236
rect	373	236	374	237
rect	373	237	374	238
rect	373	238	374	239
rect	373	239	374	240
rect	373	240	374	241
rect	373	241	374	242
rect	373	242	374	243
rect	373	243	374	244
rect	373	244	374	245
rect	373	245	374	246
rect	373	246	374	247
rect	373	247	374	248
rect	373	248	374	249
rect	373	249	374	250
rect	373	250	374	251
rect	373	251	374	252
rect	373	252	374	253
rect	373	253	374	254
rect	373	254	374	255
rect	373	255	374	256
rect	373	256	374	257
rect	373	257	374	258
rect	373	258	374	259
rect	373	259	374	260
rect	373	260	374	261
rect	373	261	374	262
rect	373	262	374	263
rect	373	263	374	264
rect	373	264	374	265
rect	373	265	374	266
rect	373	266	374	267
rect	373	267	374	268
rect	373	268	374	269
rect	373	269	374	270
rect	373	270	374	271
rect	373	271	374	272
rect	373	272	374	273
rect	373	273	374	274
rect	373	274	374	275
rect	373	275	374	276
rect	373	276	374	277
rect	373	277	374	278
rect	373	278	374	279
rect	373	279	374	280
rect	373	280	374	281
rect	373	281	374	282
rect	373	282	374	283
rect	373	283	374	284
rect	373	284	374	285
rect	373	285	374	286
rect	373	286	374	287
rect	373	287	374	288
rect	373	288	374	289
rect	373	289	374	290
rect	373	290	374	291
rect	373	291	374	292
rect	373	292	374	293
rect	373	293	374	294
rect	373	294	374	295
rect	373	295	374	296
rect	373	296	374	297
rect	373	297	374	298
rect	373	298	374	299
rect	373	299	374	300
rect	373	300	374	301
rect	373	301	374	302
rect	373	302	374	303
rect	373	303	374	304
rect	373	304	374	305
rect	373	305	374	306
rect	373	306	374	307
rect	373	307	374	308
rect	373	308	374	309
rect	373	309	374	310
rect	373	310	374	311
rect	373	311	374	312
rect	373	312	374	313
rect	373	313	374	314
rect	373	314	374	315
rect	373	315	374	316
rect	373	316	374	317
rect	373	317	374	318
rect	373	318	374	319
rect	373	319	374	320
rect	373	320	374	321
rect	373	321	374	322
rect	373	322	374	323
rect	373	323	374	324
rect	373	324	374	325
rect	373	325	374	326
rect	373	326	374	327
rect	373	327	374	328
rect	373	328	374	329
rect	373	329	374	330
rect	373	330	374	331
rect	373	331	374	332
rect	373	332	374	333
rect	373	333	374	334
rect	373	334	374	335
rect	373	335	374	336
rect	373	336	374	337
rect	373	337	374	338
rect	373	338	374	339
rect	373	339	374	340
rect	373	340	374	341
rect	373	341	374	342
rect	373	342	374	343
rect	373	343	374	344
rect	373	344	374	345
rect	373	345	374	346
rect	373	346	374	347
rect	373	347	374	348
rect	373	348	374	349
rect	373	349	374	350
rect	373	350	374	351
rect	373	351	374	352
rect	373	352	374	353
rect	373	353	374	354
rect	373	354	374	355
rect	373	355	374	356
rect	373	356	374	357
rect	373	357	374	358
rect	373	358	374	359
rect	373	359	374	360
rect	373	360	374	361
rect	373	361	374	362
rect	373	362	374	363
rect	373	363	374	364
rect	373	364	374	365
rect	373	365	374	366
rect	373	366	374	367
rect	373	367	374	368
rect	373	368	374	369
rect	374	0	375	1
rect	374	1	375	2
rect	374	2	375	3
rect	374	3	375	4
rect	374	4	375	5
rect	374	5	375	6
rect	374	6	375	7
rect	374	7	375	8
rect	374	8	375	9
rect	374	9	375	10
rect	374	10	375	11
rect	374	11	375	12
rect	374	12	375	13
rect	374	13	375	14
rect	374	14	375	15
rect	374	15	375	16
rect	374	16	375	17
rect	374	17	375	18
rect	374	18	375	19
rect	374	19	375	20
rect	374	20	375	21
rect	374	21	375	22
rect	374	22	375	23
rect	374	23	375	24
rect	374	24	375	25
rect	374	25	375	26
rect	374	26	375	27
rect	374	27	375	28
rect	374	28	375	29
rect	374	29	375	30
rect	374	30	375	31
rect	374	31	375	32
rect	374	32	375	33
rect	374	33	375	34
rect	374	34	375	35
rect	374	35	375	36
rect	374	36	375	37
rect	374	37	375	38
rect	374	38	375	39
rect	374	39	375	40
rect	374	40	375	41
rect	374	41	375	42
rect	374	42	375	43
rect	374	43	375	44
rect	374	44	375	45
rect	374	45	375	46
rect	374	46	375	47
rect	374	47	375	48
rect	374	48	375	49
rect	374	49	375	50
rect	374	50	375	51
rect	374	51	375	52
rect	374	52	375	53
rect	374	53	375	54
rect	374	54	375	55
rect	374	55	375	56
rect	374	56	375	57
rect	374	57	375	58
rect	374	58	375	59
rect	374	59	375	60
rect	374	60	375	61
rect	374	61	375	62
rect	374	62	375	63
rect	374	63	375	64
rect	374	64	375	65
rect	374	65	375	66
rect	374	66	375	67
rect	374	67	375	68
rect	374	68	375	69
rect	374	69	375	70
rect	374	70	375	71
rect	374	71	375	72
rect	374	72	375	73
rect	374	73	375	74
rect	374	74	375	75
rect	374	75	375	76
rect	374	76	375	77
rect	374	77	375	78
rect	374	78	375	79
rect	374	79	375	80
rect	374	80	375	81
rect	374	81	375	82
rect	374	82	375	83
rect	374	83	375	84
rect	374	84	375	85
rect	374	85	375	86
rect	374	86	375	87
rect	374	87	375	88
rect	374	88	375	89
rect	374	89	375	90
rect	374	90	375	91
rect	374	91	375	92
rect	374	92	375	93
rect	374	93	375	94
rect	374	94	375	95
rect	374	95	375	96
rect	374	96	375	97
rect	374	97	375	98
rect	374	98	375	99
rect	374	99	375	100
rect	374	100	375	101
rect	374	101	375	102
rect	374	102	375	103
rect	374	103	375	104
rect	374	104	375	105
rect	374	105	375	106
rect	374	106	375	107
rect	374	107	375	108
rect	374	108	375	109
rect	374	109	375	110
rect	374	110	375	111
rect	374	111	375	112
rect	374	112	375	113
rect	374	113	375	114
rect	374	114	375	115
rect	374	115	375	116
rect	374	116	375	117
rect	374	117	375	118
rect	374	118	375	119
rect	374	119	375	120
rect	374	120	375	121
rect	374	121	375	122
rect	374	122	375	123
rect	374	123	375	124
rect	374	124	375	125
rect	374	125	375	126
rect	374	126	375	127
rect	374	127	375	128
rect	374	128	375	129
rect	374	129	375	130
rect	374	130	375	131
rect	374	131	375	132
rect	374	132	375	133
rect	374	133	375	134
rect	374	134	375	135
rect	374	135	375	136
rect	374	136	375	137
rect	374	137	375	138
rect	374	138	375	139
rect	374	139	375	140
rect	374	140	375	141
rect	374	141	375	142
rect	374	142	375	143
rect	374	143	375	144
rect	374	144	375	145
rect	374	145	375	146
rect	374	146	375	147
rect	374	147	375	148
rect	374	148	375	149
rect	374	149	375	150
rect	374	150	375	151
rect	374	151	375	152
rect	374	152	375	153
rect	374	153	375	154
rect	374	154	375	155
rect	374	155	375	156
rect	374	156	375	157
rect	374	157	375	158
rect	374	158	375	159
rect	374	159	375	160
rect	374	160	375	161
rect	374	161	375	162
rect	374	162	375	163
rect	374	163	375	164
rect	374	164	375	165
rect	374	165	375	166
rect	374	166	375	167
rect	374	167	375	168
rect	374	168	375	169
rect	374	169	375	170
rect	374	170	375	171
rect	374	171	375	172
rect	374	172	375	173
rect	374	173	375	174
rect	374	174	375	175
rect	374	175	375	176
rect	374	176	375	177
rect	374	177	375	178
rect	374	178	375	179
rect	374	179	375	180
rect	374	180	375	181
rect	374	181	375	182
rect	374	182	375	183
rect	374	183	375	184
rect	374	184	375	185
rect	374	185	375	186
rect	374	186	375	187
rect	374	187	375	188
rect	374	188	375	189
rect	374	189	375	190
rect	374	190	375	191
rect	374	191	375	192
rect	374	192	375	193
rect	374	193	375	194
rect	374	194	375	195
rect	374	195	375	196
rect	374	196	375	197
rect	374	197	375	198
rect	374	198	375	199
rect	374	199	375	200
rect	374	200	375	201
rect	374	201	375	202
rect	374	202	375	203
rect	374	203	375	204
rect	374	204	375	205
rect	374	205	375	206
rect	374	206	375	207
rect	374	207	375	208
rect	374	208	375	209
rect	374	209	375	210
rect	374	210	375	211
rect	374	211	375	212
rect	374	212	375	213
rect	374	213	375	214
rect	374	214	375	215
rect	374	215	375	216
rect	374	216	375	217
rect	374	217	375	218
rect	374	218	375	219
rect	374	219	375	220
rect	374	220	375	221
rect	374	221	375	222
rect	374	222	375	223
rect	374	223	375	224
rect	374	224	375	225
rect	374	225	375	226
rect	374	226	375	227
rect	374	227	375	228
rect	374	228	375	229
rect	374	229	375	230
rect	374	230	375	231
rect	374	231	375	232
rect	374	232	375	233
rect	374	233	375	234
rect	374	234	375	235
rect	374	235	375	236
rect	374	236	375	237
rect	374	237	375	238
rect	374	238	375	239
rect	374	239	375	240
rect	374	240	375	241
rect	374	241	375	242
rect	374	242	375	243
rect	374	243	375	244
rect	374	244	375	245
rect	374	245	375	246
rect	374	246	375	247
rect	374	247	375	248
rect	374	248	375	249
rect	374	249	375	250
rect	374	250	375	251
rect	374	251	375	252
rect	374	252	375	253
rect	374	253	375	254
rect	374	254	375	255
rect	374	255	375	256
rect	374	256	375	257
rect	374	257	375	258
rect	374	258	375	259
rect	374	259	375	260
rect	374	260	375	261
rect	374	261	375	262
rect	374	262	375	263
rect	374	263	375	264
rect	374	264	375	265
rect	374	265	375	266
rect	374	266	375	267
rect	374	267	375	268
rect	374	268	375	269
rect	374	269	375	270
rect	374	270	375	271
rect	374	271	375	272
rect	374	272	375	273
rect	374	273	375	274
rect	374	274	375	275
rect	374	275	375	276
rect	374	276	375	277
rect	374	277	375	278
rect	374	278	375	279
rect	374	279	375	280
rect	374	280	375	281
rect	374	281	375	282
rect	374	282	375	283
rect	374	283	375	284
rect	374	284	375	285
rect	374	285	375	286
rect	374	286	375	287
rect	374	287	375	288
rect	374	288	375	289
rect	374	289	375	290
rect	374	290	375	291
rect	374	291	375	292
rect	374	292	375	293
rect	374	293	375	294
rect	374	294	375	295
rect	374	295	375	296
rect	374	296	375	297
rect	374	297	375	298
rect	374	298	375	299
rect	374	299	375	300
rect	374	300	375	301
rect	374	301	375	302
rect	374	302	375	303
rect	374	303	375	304
rect	374	304	375	305
rect	374	305	375	306
rect	374	306	375	307
rect	374	307	375	308
rect	374	308	375	309
rect	374	309	375	310
rect	374	310	375	311
rect	374	311	375	312
rect	374	312	375	313
rect	374	313	375	314
rect	374	314	375	315
rect	374	315	375	316
rect	374	316	375	317
rect	374	317	375	318
rect	374	318	375	319
rect	374	319	375	320
rect	374	320	375	321
rect	374	321	375	322
rect	374	322	375	323
rect	374	323	375	324
rect	374	324	375	325
rect	374	325	375	326
rect	374	326	375	327
rect	374	327	375	328
rect	374	328	375	329
rect	374	329	375	330
rect	374	330	375	331
rect	374	331	375	332
rect	374	332	375	333
rect	374	333	375	334
rect	374	334	375	335
rect	374	335	375	336
rect	374	336	375	337
rect	374	337	375	338
rect	374	338	375	339
rect	374	339	375	340
rect	374	340	375	341
rect	374	341	375	342
rect	374	342	375	343
rect	374	343	375	344
rect	374	344	375	345
rect	374	345	375	346
rect	374	346	375	347
rect	374	347	375	348
rect	374	348	375	349
rect	374	349	375	350
rect	374	350	375	351
rect	374	351	375	352
rect	374	352	375	353
rect	374	353	375	354
rect	374	354	375	355
rect	374	355	375	356
rect	374	356	375	357
rect	374	357	375	358
rect	374	358	375	359
rect	374	359	375	360
rect	374	360	375	361
rect	374	361	375	362
rect	374	362	375	363
rect	374	363	375	364
rect	374	364	375	365
rect	374	365	375	366
rect	374	366	375	367
rect	374	367	375	368
rect	374	368	375	369
rect	375	0	376	1
rect	375	1	376	2
rect	375	2	376	3
rect	375	3	376	4
rect	375	4	376	5
rect	375	5	376	6
rect	375	6	376	7
rect	375	7	376	8
rect	375	8	376	9
rect	375	9	376	10
rect	375	10	376	11
rect	375	11	376	12
rect	375	12	376	13
rect	375	13	376	14
rect	375	14	376	15
rect	375	15	376	16
rect	375	16	376	17
rect	375	17	376	18
rect	375	18	376	19
rect	375	19	376	20
rect	375	20	376	21
rect	375	21	376	22
rect	375	22	376	23
rect	375	23	376	24
rect	375	24	376	25
rect	375	25	376	26
rect	375	26	376	27
rect	375	27	376	28
rect	375	28	376	29
rect	375	29	376	30
rect	375	30	376	31
rect	375	31	376	32
rect	375	32	376	33
rect	375	33	376	34
rect	375	34	376	35
rect	375	35	376	36
rect	375	36	376	37
rect	375	37	376	38
rect	375	38	376	39
rect	375	39	376	40
rect	375	40	376	41
rect	375	41	376	42
rect	375	42	376	43
rect	375	43	376	44
rect	375	44	376	45
rect	375	45	376	46
rect	375	46	376	47
rect	375	47	376	48
rect	375	48	376	49
rect	375	49	376	50
rect	375	50	376	51
rect	375	51	376	52
rect	375	52	376	53
rect	375	53	376	54
rect	375	54	376	55
rect	375	55	376	56
rect	375	56	376	57
rect	375	57	376	58
rect	375	58	376	59
rect	375	59	376	60
rect	375	60	376	61
rect	375	61	376	62
rect	375	62	376	63
rect	375	63	376	64
rect	375	64	376	65
rect	375	65	376	66
rect	375	66	376	67
rect	375	67	376	68
rect	375	68	376	69
rect	375	69	376	70
rect	375	70	376	71
rect	375	71	376	72
rect	375	72	376	73
rect	375	73	376	74
rect	375	74	376	75
rect	375	75	376	76
rect	375	76	376	77
rect	375	77	376	78
rect	375	78	376	79
rect	375	79	376	80
rect	375	80	376	81
rect	375	81	376	82
rect	375	82	376	83
rect	375	83	376	84
rect	375	84	376	85
rect	375	85	376	86
rect	375	86	376	87
rect	375	87	376	88
rect	375	88	376	89
rect	375	89	376	90
rect	375	90	376	91
rect	375	91	376	92
rect	375	92	376	93
rect	375	93	376	94
rect	375	94	376	95
rect	375	95	376	96
rect	375	96	376	97
rect	375	97	376	98
rect	375	98	376	99
rect	375	99	376	100
rect	375	100	376	101
rect	375	101	376	102
rect	375	102	376	103
rect	375	103	376	104
rect	375	104	376	105
rect	375	105	376	106
rect	375	106	376	107
rect	375	107	376	108
rect	375	108	376	109
rect	375	109	376	110
rect	375	110	376	111
rect	375	111	376	112
rect	375	112	376	113
rect	375	113	376	114
rect	375	114	376	115
rect	375	115	376	116
rect	375	116	376	117
rect	375	117	376	118
rect	375	118	376	119
rect	375	119	376	120
rect	375	120	376	121
rect	375	121	376	122
rect	375	122	376	123
rect	375	123	376	124
rect	375	124	376	125
rect	375	125	376	126
rect	375	126	376	127
rect	375	127	376	128
rect	375	128	376	129
rect	375	129	376	130
rect	375	130	376	131
rect	375	131	376	132
rect	375	132	376	133
rect	375	133	376	134
rect	375	134	376	135
rect	375	135	376	136
rect	375	136	376	137
rect	375	137	376	138
rect	375	138	376	139
rect	375	139	376	140
rect	375	140	376	141
rect	375	141	376	142
rect	375	142	376	143
rect	375	143	376	144
rect	375	144	376	145
rect	375	145	376	146
rect	375	146	376	147
rect	375	147	376	148
rect	375	148	376	149
rect	375	149	376	150
rect	375	150	376	151
rect	375	151	376	152
rect	375	152	376	153
rect	375	153	376	154
rect	375	154	376	155
rect	375	155	376	156
rect	375	156	376	157
rect	375	157	376	158
rect	375	158	376	159
rect	375	159	376	160
rect	375	160	376	161
rect	375	161	376	162
rect	375	162	376	163
rect	375	163	376	164
rect	375	164	376	165
rect	375	165	376	166
rect	375	166	376	167
rect	375	167	376	168
rect	375	168	376	169
rect	375	169	376	170
rect	375	170	376	171
rect	375	171	376	172
rect	375	172	376	173
rect	375	173	376	174
rect	375	174	376	175
rect	375	175	376	176
rect	375	176	376	177
rect	375	177	376	178
rect	375	178	376	179
rect	375	179	376	180
rect	375	180	376	181
rect	375	181	376	182
rect	375	182	376	183
rect	375	183	376	184
rect	375	184	376	185
rect	375	185	376	186
rect	375	186	376	187
rect	375	187	376	188
rect	375	188	376	189
rect	375	189	376	190
rect	375	190	376	191
rect	375	191	376	192
rect	375	192	376	193
rect	375	193	376	194
rect	375	194	376	195
rect	375	195	376	196
rect	375	196	376	197
rect	375	197	376	198
rect	375	198	376	199
rect	375	199	376	200
rect	375	200	376	201
rect	375	201	376	202
rect	375	202	376	203
rect	375	203	376	204
rect	375	204	376	205
rect	375	205	376	206
rect	375	206	376	207
rect	375	207	376	208
rect	375	208	376	209
rect	375	209	376	210
rect	375	210	376	211
rect	375	211	376	212
rect	375	212	376	213
rect	375	213	376	214
rect	375	214	376	215
rect	375	215	376	216
rect	375	216	376	217
rect	375	217	376	218
rect	375	218	376	219
rect	375	219	376	220
rect	375	220	376	221
rect	375	221	376	222
rect	375	222	376	223
rect	375	223	376	224
rect	375	224	376	225
rect	375	225	376	226
rect	375	226	376	227
rect	375	227	376	228
rect	375	228	376	229
rect	375	229	376	230
rect	375	230	376	231
rect	375	231	376	232
rect	375	232	376	233
rect	375	233	376	234
rect	375	234	376	235
rect	375	235	376	236
rect	375	236	376	237
rect	375	237	376	238
rect	375	238	376	239
rect	375	239	376	240
rect	375	240	376	241
rect	375	241	376	242
rect	375	242	376	243
rect	375	243	376	244
rect	375	244	376	245
rect	375	245	376	246
rect	375	246	376	247
rect	375	247	376	248
rect	375	248	376	249
rect	375	249	376	250
rect	375	250	376	251
rect	375	251	376	252
rect	375	252	376	253
rect	375	253	376	254
rect	375	254	376	255
rect	375	255	376	256
rect	375	256	376	257
rect	375	257	376	258
rect	375	258	376	259
rect	375	259	376	260
rect	375	260	376	261
rect	375	261	376	262
rect	375	262	376	263
rect	375	263	376	264
rect	375	264	376	265
rect	375	265	376	266
rect	375	266	376	267
rect	375	267	376	268
rect	375	268	376	269
rect	375	269	376	270
rect	375	270	376	271
rect	375	271	376	272
rect	375	272	376	273
rect	375	273	376	274
rect	375	274	376	275
rect	375	275	376	276
rect	375	276	376	277
rect	375	277	376	278
rect	375	278	376	279
rect	375	279	376	280
rect	375	280	376	281
rect	375	281	376	282
rect	375	282	376	283
rect	375	283	376	284
rect	375	284	376	285
rect	375	285	376	286
rect	375	286	376	287
rect	375	287	376	288
rect	375	288	376	289
rect	375	289	376	290
rect	375	290	376	291
rect	375	291	376	292
rect	375	292	376	293
rect	375	293	376	294
rect	375	294	376	295
rect	375	295	376	296
rect	375	296	376	297
rect	375	297	376	298
rect	375	298	376	299
rect	375	299	376	300
rect	375	300	376	301
rect	375	301	376	302
rect	375	302	376	303
rect	375	303	376	304
rect	375	304	376	305
rect	375	305	376	306
rect	375	306	376	307
rect	375	307	376	308
rect	375	308	376	309
rect	375	309	376	310
rect	375	310	376	311
rect	375	311	376	312
rect	375	312	376	313
rect	375	313	376	314
rect	375	314	376	315
rect	375	315	376	316
rect	375	316	376	317
rect	375	317	376	318
rect	375	318	376	319
rect	375	319	376	320
rect	375	320	376	321
rect	375	321	376	322
rect	375	322	376	323
rect	375	323	376	324
rect	375	324	376	325
rect	375	325	376	326
rect	375	326	376	327
rect	375	327	376	328
rect	375	328	376	329
rect	375	329	376	330
rect	375	330	376	331
rect	375	331	376	332
rect	375	332	376	333
rect	375	333	376	334
rect	375	334	376	335
rect	375	335	376	336
rect	375	336	376	337
rect	375	337	376	338
rect	375	338	376	339
rect	375	339	376	340
rect	375	340	376	341
rect	375	341	376	342
rect	375	342	376	343
rect	375	343	376	344
rect	375	344	376	345
rect	375	345	376	346
rect	375	346	376	347
rect	375	347	376	348
rect	375	348	376	349
rect	375	349	376	350
rect	375	350	376	351
rect	375	351	376	352
rect	375	352	376	353
rect	375	353	376	354
rect	375	354	376	355
rect	375	355	376	356
rect	375	356	376	357
rect	375	357	376	358
rect	375	358	376	359
rect	375	359	376	360
rect	375	360	376	361
rect	375	361	376	362
rect	375	362	376	363
rect	375	363	376	364
rect	375	364	376	365
rect	375	365	376	366
rect	375	366	376	367
rect	375	367	376	368
rect	375	368	376	369
rect	421	0	422	1
rect	421	1	422	2
rect	421	2	422	3
rect	421	3	422	4
rect	421	4	422	5
rect	421	5	422	6
rect	421	6	422	7
rect	421	7	422	8
rect	421	8	422	9
rect	421	9	422	10
rect	421	10	422	11
rect	421	11	422	12
rect	421	12	422	13
rect	421	13	422	14
rect	421	14	422	15
rect	421	15	422	16
rect	421	16	422	17
rect	421	17	422	18
rect	421	18	422	19
rect	421	19	422	20
rect	421	20	422	21
rect	421	21	422	22
rect	421	22	422	23
rect	421	23	422	24
rect	421	24	422	25
rect	421	25	422	26
rect	421	26	422	27
rect	421	27	422	28
rect	421	28	422	29
rect	421	29	422	30
rect	421	30	422	31
rect	421	31	422	32
rect	421	32	422	33
rect	421	33	422	34
rect	421	34	422	35
rect	421	35	422	36
rect	421	36	422	37
rect	421	37	422	38
rect	421	38	422	39
rect	421	39	422	40
rect	421	40	422	41
rect	421	41	422	42
rect	421	42	422	43
rect	421	43	422	44
rect	421	44	422	45
rect	421	45	422	46
rect	421	46	422	47
rect	421	47	422	48
rect	421	48	422	49
rect	421	49	422	50
rect	421	50	422	51
rect	421	51	422	52
rect	421	52	422	53
rect	421	53	422	54
rect	421	54	422	55
rect	421	55	422	56
rect	421	56	422	57
rect	421	57	422	58
rect	421	58	422	59
rect	421	59	422	60
rect	421	60	422	61
rect	421	61	422	62
rect	421	62	422	63
rect	421	63	422	64
rect	421	64	422	65
rect	421	65	422	66
rect	421	66	422	67
rect	421	67	422	68
rect	421	68	422	69
rect	421	69	422	70
rect	421	70	422	71
rect	421	71	422	72
rect	421	72	422	73
rect	421	73	422	74
rect	421	74	422	75
rect	421	75	422	76
rect	421	76	422	77
rect	421	77	422	78
rect	421	78	422	79
rect	421	79	422	80
rect	421	80	422	81
rect	421	81	422	82
rect	421	82	422	83
rect	421	83	422	84
rect	421	84	422	85
rect	421	85	422	86
rect	421	86	422	87
rect	421	87	422	88
rect	421	88	422	89
rect	421	89	422	90
rect	421	90	422	91
rect	421	91	422	92
rect	421	92	422	93
rect	421	93	422	94
rect	421	94	422	95
rect	421	95	422	96
rect	421	96	422	97
rect	421	97	422	98
rect	421	98	422	99
rect	421	99	422	100
rect	421	100	422	101
rect	421	101	422	102
rect	421	102	422	103
rect	421	103	422	104
rect	421	104	422	105
rect	421	105	422	106
rect	421	106	422	107
rect	421	107	422	108
rect	421	108	422	109
rect	421	109	422	110
rect	421	110	422	111
rect	421	111	422	112
rect	421	112	422	113
rect	421	113	422	114
rect	421	114	422	115
rect	421	115	422	116
rect	421	116	422	117
rect	421	117	422	118
rect	421	118	422	119
rect	421	119	422	120
rect	421	120	422	121
rect	421	121	422	122
rect	421	122	422	123
rect	421	123	422	124
rect	421	124	422	125
rect	421	125	422	126
rect	421	126	422	127
rect	421	127	422	128
rect	421	128	422	129
rect	421	129	422	130
rect	421	130	422	131
rect	421	131	422	132
rect	421	132	422	133
rect	421	133	422	134
rect	421	134	422	135
rect	421	135	422	136
rect	421	136	422	137
rect	421	137	422	138
rect	421	138	422	139
rect	421	139	422	140
rect	421	140	422	141
rect	421	141	422	142
rect	421	142	422	143
rect	421	143	422	144
rect	421	144	422	145
rect	421	145	422	146
rect	421	146	422	147
rect	421	147	422	148
rect	421	148	422	149
rect	421	149	422	150
rect	421	150	422	151
rect	421	151	422	152
rect	421	152	422	153
rect	421	153	422	154
rect	421	154	422	155
rect	421	155	422	156
rect	421	156	422	157
rect	421	157	422	158
rect	421	158	422	159
rect	421	159	422	160
rect	421	160	422	161
rect	421	161	422	162
rect	421	162	422	163
rect	421	163	422	164
rect	421	164	422	165
rect	421	165	422	166
rect	421	166	422	167
rect	421	167	422	168
rect	421	168	422	169
rect	421	169	422	170
rect	421	170	422	171
rect	421	171	422	172
rect	421	172	422	173
rect	421	173	422	174
rect	421	174	422	175
rect	421	175	422	176
rect	421	176	422	177
rect	421	177	422	178
rect	421	178	422	179
rect	421	179	422	180
rect	421	180	422	181
rect	421	181	422	182
rect	421	182	422	183
rect	421	183	422	184
rect	421	184	422	185
rect	421	185	422	186
rect	421	186	422	187
rect	421	187	422	188
rect	421	188	422	189
rect	421	189	422	190
rect	421	190	422	191
rect	421	191	422	192
rect	421	192	422	193
rect	421	193	422	194
rect	421	194	422	195
rect	421	195	422	196
rect	421	196	422	197
rect	421	197	422	198
rect	421	198	422	199
rect	421	199	422	200
rect	421	200	422	201
rect	421	201	422	202
rect	421	202	422	203
rect	421	203	422	204
rect	421	204	422	205
rect	421	205	422	206
rect	421	206	422	207
rect	421	207	422	208
rect	421	208	422	209
rect	421	209	422	210
rect	421	210	422	211
rect	421	211	422	212
rect	421	212	422	213
rect	421	213	422	214
rect	421	214	422	215
rect	421	215	422	216
rect	421	216	422	217
rect	421	217	422	218
rect	421	218	422	219
rect	421	219	422	220
rect	421	220	422	221
rect	421	221	422	222
rect	421	222	422	223
rect	421	223	422	224
rect	421	224	422	225
rect	421	225	422	226
rect	421	226	422	227
rect	421	227	422	228
rect	421	228	422	229
rect	421	229	422	230
rect	421	230	422	231
rect	421	231	422	232
rect	421	232	422	233
rect	421	233	422	234
rect	421	234	422	235
rect	421	235	422	236
rect	421	236	422	237
rect	421	237	422	238
rect	421	238	422	239
rect	421	239	422	240
rect	421	240	422	241
rect	421	241	422	242
rect	421	242	422	243
rect	421	243	422	244
rect	421	244	422	245
rect	421	245	422	246
rect	421	246	422	247
rect	421	247	422	248
rect	421	248	422	249
rect	421	249	422	250
rect	421	250	422	251
rect	421	251	422	252
rect	421	252	422	253
rect	421	253	422	254
rect	421	254	422	255
rect	421	255	422	256
rect	421	256	422	257
rect	421	257	422	258
rect	421	258	422	259
rect	421	259	422	260
rect	421	260	422	261
rect	421	261	422	262
rect	421	262	422	263
rect	421	263	422	264
rect	421	264	422	265
rect	421	265	422	266
rect	421	266	422	267
rect	421	267	422	268
rect	421	268	422	269
rect	421	269	422	270
rect	421	270	422	271
rect	421	271	422	272
rect	421	272	422	273
rect	421	273	422	274
rect	421	274	422	275
rect	421	275	422	276
rect	421	276	422	277
rect	421	277	422	278
rect	421	278	422	279
rect	421	279	422	280
rect	421	280	422	281
rect	421	281	422	282
rect	421	282	422	283
rect	421	283	422	284
rect	421	284	422	285
rect	421	285	422	286
rect	421	286	422	287
rect	421	287	422	288
rect	421	288	422	289
rect	421	289	422	290
rect	421	290	422	291
rect	421	291	422	292
rect	421	292	422	293
rect	421	293	422	294
rect	421	294	422	295
rect	421	295	422	296
rect	421	296	422	297
rect	421	297	422	298
rect	421	298	422	299
rect	421	299	422	300
rect	421	300	422	301
rect	421	301	422	302
rect	421	302	422	303
rect	421	303	422	304
rect	421	304	422	305
rect	421	305	422	306
rect	421	306	422	307
rect	421	307	422	308
rect	421	308	422	309
rect	421	309	422	310
rect	421	310	422	311
rect	421	311	422	312
rect	421	312	422	313
rect	421	313	422	314
rect	421	314	422	315
rect	421	315	422	316
rect	421	316	422	317
rect	421	317	422	318
rect	421	318	422	319
rect	421	319	422	320
rect	421	320	422	321
rect	421	321	422	322
rect	421	322	422	323
rect	421	323	422	324
rect	421	324	422	325
rect	421	325	422	326
rect	421	326	422	327
rect	421	327	422	328
rect	421	328	422	329
rect	421	329	422	330
rect	421	330	422	331
rect	421	331	422	332
rect	421	332	422	333
rect	421	333	422	334
rect	421	334	422	335
rect	421	335	422	336
rect	421	336	422	337
rect	421	337	422	338
rect	421	338	422	339
rect	421	339	422	340
rect	421	340	422	341
rect	421	341	422	342
rect	421	342	422	343
rect	421	343	422	344
rect	421	344	422	345
rect	421	345	422	346
rect	421	346	422	347
rect	421	347	422	348
rect	421	348	422	349
rect	421	349	422	350
rect	421	350	422	351
rect	421	351	422	352
rect	421	352	422	353
rect	421	353	422	354
rect	421	354	422	355
rect	421	355	422	356
rect	421	356	422	357
rect	421	357	422	358
rect	421	358	422	359
rect	421	359	422	360
rect	421	360	422	361
rect	421	361	422	362
rect	421	362	422	363
rect	421	363	422	364
rect	421	364	422	365
rect	421	365	422	366
rect	421	366	422	367
rect	421	367	422	368
rect	421	368	422	369
rect	422	0	423	1
rect	422	1	423	2
rect	422	2	423	3
rect	422	3	423	4
rect	422	4	423	5
rect	422	5	423	6
rect	422	6	423	7
rect	422	7	423	8
rect	422	8	423	9
rect	422	9	423	10
rect	422	10	423	11
rect	422	11	423	12
rect	422	12	423	13
rect	422	13	423	14
rect	422	14	423	15
rect	422	15	423	16
rect	422	16	423	17
rect	422	17	423	18
rect	422	18	423	19
rect	422	19	423	20
rect	422	20	423	21
rect	422	21	423	22
rect	422	22	423	23
rect	422	23	423	24
rect	422	24	423	25
rect	422	25	423	26
rect	422	26	423	27
rect	422	27	423	28
rect	422	28	423	29
rect	422	29	423	30
rect	422	30	423	31
rect	422	31	423	32
rect	422	32	423	33
rect	422	33	423	34
rect	422	34	423	35
rect	422	35	423	36
rect	422	36	423	37
rect	422	37	423	38
rect	422	38	423	39
rect	422	39	423	40
rect	422	40	423	41
rect	422	41	423	42
rect	422	42	423	43
rect	422	43	423	44
rect	422	44	423	45
rect	422	45	423	46
rect	422	46	423	47
rect	422	47	423	48
rect	422	48	423	49
rect	422	49	423	50
rect	422	50	423	51
rect	422	51	423	52
rect	422	52	423	53
rect	422	53	423	54
rect	422	54	423	55
rect	422	55	423	56
rect	422	56	423	57
rect	422	57	423	58
rect	422	58	423	59
rect	422	59	423	60
rect	422	60	423	61
rect	422	61	423	62
rect	422	62	423	63
rect	422	63	423	64
rect	422	64	423	65
rect	422	65	423	66
rect	422	66	423	67
rect	422	67	423	68
rect	422	68	423	69
rect	422	69	423	70
rect	422	70	423	71
rect	422	71	423	72
rect	422	72	423	73
rect	422	73	423	74
rect	422	74	423	75
rect	422	75	423	76
rect	422	76	423	77
rect	422	77	423	78
rect	422	78	423	79
rect	422	79	423	80
rect	422	80	423	81
rect	422	81	423	82
rect	422	82	423	83
rect	422	83	423	84
rect	422	84	423	85
rect	422	85	423	86
rect	422	86	423	87
rect	422	87	423	88
rect	422	88	423	89
rect	422	89	423	90
rect	422	90	423	91
rect	422	91	423	92
rect	422	92	423	93
rect	422	93	423	94
rect	422	94	423	95
rect	422	95	423	96
rect	422	96	423	97
rect	422	97	423	98
rect	422	98	423	99
rect	422	99	423	100
rect	422	100	423	101
rect	422	101	423	102
rect	422	102	423	103
rect	422	103	423	104
rect	422	104	423	105
rect	422	105	423	106
rect	422	106	423	107
rect	422	107	423	108
rect	422	108	423	109
rect	422	109	423	110
rect	422	110	423	111
rect	422	111	423	112
rect	422	112	423	113
rect	422	113	423	114
rect	422	114	423	115
rect	422	115	423	116
rect	422	116	423	117
rect	422	117	423	118
rect	422	118	423	119
rect	422	119	423	120
rect	422	120	423	121
rect	422	121	423	122
rect	422	122	423	123
rect	422	123	423	124
rect	422	124	423	125
rect	422	125	423	126
rect	422	126	423	127
rect	422	127	423	128
rect	422	128	423	129
rect	422	129	423	130
rect	422	130	423	131
rect	422	131	423	132
rect	422	132	423	133
rect	422	133	423	134
rect	422	134	423	135
rect	422	135	423	136
rect	422	136	423	137
rect	422	137	423	138
rect	422	138	423	139
rect	422	139	423	140
rect	422	140	423	141
rect	422	141	423	142
rect	422	142	423	143
rect	422	143	423	144
rect	422	144	423	145
rect	422	145	423	146
rect	422	146	423	147
rect	422	147	423	148
rect	422	148	423	149
rect	422	149	423	150
rect	422	150	423	151
rect	422	151	423	152
rect	422	152	423	153
rect	422	153	423	154
rect	422	154	423	155
rect	422	155	423	156
rect	422	156	423	157
rect	422	157	423	158
rect	422	158	423	159
rect	422	159	423	160
rect	422	160	423	161
rect	422	161	423	162
rect	422	162	423	163
rect	422	163	423	164
rect	422	164	423	165
rect	422	165	423	166
rect	422	166	423	167
rect	422	167	423	168
rect	422	168	423	169
rect	422	169	423	170
rect	422	170	423	171
rect	422	171	423	172
rect	422	172	423	173
rect	422	173	423	174
rect	422	174	423	175
rect	422	175	423	176
rect	422	176	423	177
rect	422	177	423	178
rect	422	178	423	179
rect	422	179	423	180
rect	422	180	423	181
rect	422	181	423	182
rect	422	182	423	183
rect	422	183	423	184
rect	422	184	423	185
rect	422	185	423	186
rect	422	186	423	187
rect	422	187	423	188
rect	422	188	423	189
rect	422	189	423	190
rect	422	190	423	191
rect	422	191	423	192
rect	422	192	423	193
rect	422	193	423	194
rect	422	194	423	195
rect	422	195	423	196
rect	422	196	423	197
rect	422	197	423	198
rect	422	198	423	199
rect	422	199	423	200
rect	422	200	423	201
rect	422	201	423	202
rect	422	202	423	203
rect	422	203	423	204
rect	422	204	423	205
rect	422	205	423	206
rect	422	206	423	207
rect	422	207	423	208
rect	422	208	423	209
rect	422	209	423	210
rect	422	210	423	211
rect	422	211	423	212
rect	422	212	423	213
rect	422	213	423	214
rect	422	214	423	215
rect	422	215	423	216
rect	422	216	423	217
rect	422	217	423	218
rect	422	218	423	219
rect	422	219	423	220
rect	422	220	423	221
rect	422	221	423	222
rect	422	222	423	223
rect	422	223	423	224
rect	422	224	423	225
rect	422	225	423	226
rect	422	226	423	227
rect	422	227	423	228
rect	422	228	423	229
rect	422	229	423	230
rect	422	230	423	231
rect	422	231	423	232
rect	422	232	423	233
rect	422	233	423	234
rect	422	234	423	235
rect	422	235	423	236
rect	422	236	423	237
rect	422	237	423	238
rect	422	238	423	239
rect	422	239	423	240
rect	422	240	423	241
rect	422	241	423	242
rect	422	242	423	243
rect	422	243	423	244
rect	422	244	423	245
rect	422	245	423	246
rect	422	246	423	247
rect	422	247	423	248
rect	422	248	423	249
rect	422	249	423	250
rect	422	250	423	251
rect	422	251	423	252
rect	422	252	423	253
rect	422	253	423	254
rect	422	254	423	255
rect	422	255	423	256
rect	422	256	423	257
rect	422	257	423	258
rect	422	258	423	259
rect	422	259	423	260
rect	422	260	423	261
rect	422	261	423	262
rect	422	262	423	263
rect	422	263	423	264
rect	422	264	423	265
rect	422	265	423	266
rect	422	266	423	267
rect	422	267	423	268
rect	422	268	423	269
rect	422	269	423	270
rect	422	270	423	271
rect	422	271	423	272
rect	422	272	423	273
rect	422	273	423	274
rect	422	274	423	275
rect	422	275	423	276
rect	422	276	423	277
rect	422	277	423	278
rect	422	278	423	279
rect	422	279	423	280
rect	422	280	423	281
rect	422	281	423	282
rect	422	282	423	283
rect	422	283	423	284
rect	422	284	423	285
rect	422	285	423	286
rect	422	286	423	287
rect	422	287	423	288
rect	422	288	423	289
rect	422	289	423	290
rect	422	290	423	291
rect	422	291	423	292
rect	422	292	423	293
rect	422	293	423	294
rect	422	294	423	295
rect	422	295	423	296
rect	422	296	423	297
rect	422	297	423	298
rect	422	298	423	299
rect	422	299	423	300
rect	422	300	423	301
rect	422	301	423	302
rect	422	302	423	303
rect	422	303	423	304
rect	422	304	423	305
rect	422	305	423	306
rect	422	306	423	307
rect	422	307	423	308
rect	422	308	423	309
rect	422	309	423	310
rect	422	310	423	311
rect	422	311	423	312
rect	422	312	423	313
rect	422	313	423	314
rect	422	314	423	315
rect	422	315	423	316
rect	422	316	423	317
rect	422	317	423	318
rect	422	318	423	319
rect	422	319	423	320
rect	422	320	423	321
rect	422	321	423	322
rect	422	322	423	323
rect	422	323	423	324
rect	422	324	423	325
rect	422	325	423	326
rect	422	326	423	327
rect	422	327	423	328
rect	422	328	423	329
rect	422	329	423	330
rect	422	330	423	331
rect	422	331	423	332
rect	422	332	423	333
rect	422	333	423	334
rect	422	334	423	335
rect	422	335	423	336
rect	422	336	423	337
rect	422	337	423	338
rect	422	338	423	339
rect	422	339	423	340
rect	422	340	423	341
rect	422	341	423	342
rect	422	342	423	343
rect	422	343	423	344
rect	422	344	423	345
rect	422	345	423	346
rect	422	346	423	347
rect	422	347	423	348
rect	422	348	423	349
rect	422	349	423	350
rect	422	350	423	351
rect	422	351	423	352
rect	422	352	423	353
rect	422	353	423	354
rect	422	354	423	355
rect	422	355	423	356
rect	422	356	423	357
rect	422	357	423	358
rect	422	358	423	359
rect	422	359	423	360
rect	422	360	423	361
rect	422	361	423	362
rect	422	362	423	363
rect	422	363	423	364
rect	422	364	423	365
rect	422	365	423	366
rect	422	366	423	367
rect	422	367	423	368
rect	422	368	423	369
rect	423	0	424	1
rect	423	1	424	2
rect	423	2	424	3
rect	423	3	424	4
rect	423	4	424	5
rect	423	5	424	6
rect	423	6	424	7
rect	423	7	424	8
rect	423	8	424	9
rect	423	9	424	10
rect	423	10	424	11
rect	423	11	424	12
rect	423	12	424	13
rect	423	13	424	14
rect	423	14	424	15
rect	423	15	424	16
rect	423	16	424	17
rect	423	17	424	18
rect	423	18	424	19
rect	423	19	424	20
rect	423	20	424	21
rect	423	21	424	22
rect	423	22	424	23
rect	423	23	424	24
rect	423	24	424	25
rect	423	25	424	26
rect	423	26	424	27
rect	423	27	424	28
rect	423	28	424	29
rect	423	29	424	30
rect	423	30	424	31
rect	423	31	424	32
rect	423	32	424	33
rect	423	33	424	34
rect	423	34	424	35
rect	423	35	424	36
rect	423	36	424	37
rect	423	37	424	38
rect	423	38	424	39
rect	423	39	424	40
rect	423	40	424	41
rect	423	41	424	42
rect	423	42	424	43
rect	423	43	424	44
rect	423	44	424	45
rect	423	45	424	46
rect	423	46	424	47
rect	423	47	424	48
rect	423	48	424	49
rect	423	49	424	50
rect	423	50	424	51
rect	423	51	424	52
rect	423	52	424	53
rect	423	53	424	54
rect	423	54	424	55
rect	423	55	424	56
rect	423	56	424	57
rect	423	57	424	58
rect	423	58	424	59
rect	423	59	424	60
rect	423	60	424	61
rect	423	61	424	62
rect	423	62	424	63
rect	423	63	424	64
rect	423	64	424	65
rect	423	65	424	66
rect	423	66	424	67
rect	423	67	424	68
rect	423	68	424	69
rect	423	69	424	70
rect	423	70	424	71
rect	423	71	424	72
rect	423	72	424	73
rect	423	73	424	74
rect	423	74	424	75
rect	423	75	424	76
rect	423	76	424	77
rect	423	77	424	78
rect	423	78	424	79
rect	423	79	424	80
rect	423	80	424	81
rect	423	81	424	82
rect	423	82	424	83
rect	423	83	424	84
rect	423	84	424	85
rect	423	85	424	86
rect	423	86	424	87
rect	423	87	424	88
rect	423	88	424	89
rect	423	89	424	90
rect	423	90	424	91
rect	423	91	424	92
rect	423	92	424	93
rect	423	93	424	94
rect	423	94	424	95
rect	423	95	424	96
rect	423	96	424	97
rect	423	97	424	98
rect	423	98	424	99
rect	423	99	424	100
rect	423	100	424	101
rect	423	101	424	102
rect	423	102	424	103
rect	423	103	424	104
rect	423	104	424	105
rect	423	105	424	106
rect	423	106	424	107
rect	423	107	424	108
rect	423	108	424	109
rect	423	109	424	110
rect	423	110	424	111
rect	423	111	424	112
rect	423	112	424	113
rect	423	113	424	114
rect	423	114	424	115
rect	423	115	424	116
rect	423	116	424	117
rect	423	117	424	118
rect	423	118	424	119
rect	423	119	424	120
rect	423	120	424	121
rect	423	121	424	122
rect	423	122	424	123
rect	423	123	424	124
rect	423	124	424	125
rect	423	125	424	126
rect	423	126	424	127
rect	423	127	424	128
rect	423	128	424	129
rect	423	129	424	130
rect	423	130	424	131
rect	423	131	424	132
rect	423	132	424	133
rect	423	133	424	134
rect	423	134	424	135
rect	423	135	424	136
rect	423	136	424	137
rect	423	137	424	138
rect	423	138	424	139
rect	423	139	424	140
rect	423	140	424	141
rect	423	141	424	142
rect	423	142	424	143
rect	423	143	424	144
rect	423	144	424	145
rect	423	145	424	146
rect	423	146	424	147
rect	423	147	424	148
rect	423	148	424	149
rect	423	149	424	150
rect	423	150	424	151
rect	423	151	424	152
rect	423	152	424	153
rect	423	153	424	154
rect	423	154	424	155
rect	423	155	424	156
rect	423	156	424	157
rect	423	157	424	158
rect	423	158	424	159
rect	423	159	424	160
rect	423	160	424	161
rect	423	161	424	162
rect	423	162	424	163
rect	423	163	424	164
rect	423	164	424	165
rect	423	165	424	166
rect	423	166	424	167
rect	423	167	424	168
rect	423	168	424	169
rect	423	169	424	170
rect	423	170	424	171
rect	423	171	424	172
rect	423	172	424	173
rect	423	173	424	174
rect	423	174	424	175
rect	423	175	424	176
rect	423	176	424	177
rect	423	177	424	178
rect	423	178	424	179
rect	423	179	424	180
rect	423	180	424	181
rect	423	181	424	182
rect	423	182	424	183
rect	423	183	424	184
rect	423	184	424	185
rect	423	185	424	186
rect	423	186	424	187
rect	423	187	424	188
rect	423	188	424	189
rect	423	189	424	190
rect	423	190	424	191
rect	423	191	424	192
rect	423	192	424	193
rect	423	193	424	194
rect	423	194	424	195
rect	423	195	424	196
rect	423	196	424	197
rect	423	197	424	198
rect	423	198	424	199
rect	423	199	424	200
rect	423	200	424	201
rect	423	201	424	202
rect	423	202	424	203
rect	423	203	424	204
rect	423	204	424	205
rect	423	205	424	206
rect	423	206	424	207
rect	423	207	424	208
rect	423	208	424	209
rect	423	209	424	210
rect	423	210	424	211
rect	423	211	424	212
rect	423	212	424	213
rect	423	213	424	214
rect	423	214	424	215
rect	423	215	424	216
rect	423	216	424	217
rect	423	217	424	218
rect	423	218	424	219
rect	423	219	424	220
rect	423	220	424	221
rect	423	221	424	222
rect	423	222	424	223
rect	423	223	424	224
rect	423	224	424	225
rect	423	225	424	226
rect	423	226	424	227
rect	423	227	424	228
rect	423	228	424	229
rect	423	229	424	230
rect	423	230	424	231
rect	423	231	424	232
rect	423	232	424	233
rect	423	233	424	234
rect	423	234	424	235
rect	423	235	424	236
rect	423	236	424	237
rect	423	237	424	238
rect	423	238	424	239
rect	423	239	424	240
rect	423	240	424	241
rect	423	241	424	242
rect	423	242	424	243
rect	423	243	424	244
rect	423	244	424	245
rect	423	245	424	246
rect	423	246	424	247
rect	423	247	424	248
rect	423	248	424	249
rect	423	249	424	250
rect	423	250	424	251
rect	423	251	424	252
rect	423	252	424	253
rect	423	253	424	254
rect	423	254	424	255
rect	423	255	424	256
rect	423	256	424	257
rect	423	257	424	258
rect	423	258	424	259
rect	423	259	424	260
rect	423	260	424	261
rect	423	261	424	262
rect	423	262	424	263
rect	423	263	424	264
rect	423	264	424	265
rect	423	265	424	266
rect	423	266	424	267
rect	423	267	424	268
rect	423	268	424	269
rect	423	269	424	270
rect	423	270	424	271
rect	423	271	424	272
rect	423	272	424	273
rect	423	273	424	274
rect	423	274	424	275
rect	423	275	424	276
rect	423	276	424	277
rect	423	277	424	278
rect	423	278	424	279
rect	423	279	424	280
rect	423	280	424	281
rect	423	281	424	282
rect	423	282	424	283
rect	423	283	424	284
rect	423	284	424	285
rect	423	285	424	286
rect	423	286	424	287
rect	423	287	424	288
rect	423	288	424	289
rect	423	289	424	290
rect	423	290	424	291
rect	423	291	424	292
rect	423	292	424	293
rect	423	293	424	294
rect	423	294	424	295
rect	423	295	424	296
rect	423	296	424	297
rect	423	297	424	298
rect	423	298	424	299
rect	423	299	424	300
rect	423	300	424	301
rect	423	301	424	302
rect	423	302	424	303
rect	423	303	424	304
rect	423	304	424	305
rect	423	305	424	306
rect	423	306	424	307
rect	423	307	424	308
rect	423	308	424	309
rect	423	309	424	310
rect	423	310	424	311
rect	423	311	424	312
rect	423	312	424	313
rect	423	313	424	314
rect	423	314	424	315
rect	423	315	424	316
rect	423	316	424	317
rect	423	317	424	318
rect	423	318	424	319
rect	423	319	424	320
rect	423	320	424	321
rect	423	321	424	322
rect	423	322	424	323
rect	423	323	424	324
rect	423	324	424	325
rect	423	325	424	326
rect	423	326	424	327
rect	423	327	424	328
rect	423	328	424	329
rect	423	329	424	330
rect	423	330	424	331
rect	423	331	424	332
rect	423	332	424	333
rect	423	333	424	334
rect	423	334	424	335
rect	423	335	424	336
rect	423	336	424	337
rect	423	337	424	338
rect	423	338	424	339
rect	423	339	424	340
rect	423	340	424	341
rect	423	341	424	342
rect	423	342	424	343
rect	423	343	424	344
rect	423	344	424	345
rect	423	345	424	346
rect	423	346	424	347
rect	423	347	424	348
rect	423	348	424	349
rect	423	349	424	350
rect	423	350	424	351
rect	423	351	424	352
rect	423	352	424	353
rect	423	353	424	354
rect	423	354	424	355
rect	423	355	424	356
rect	423	356	424	357
rect	423	357	424	358
rect	423	358	424	359
rect	423	359	424	360
rect	423	360	424	361
rect	423	361	424	362
rect	423	362	424	363
rect	423	363	424	364
rect	423	364	424	365
rect	423	365	424	366
rect	423	366	424	367
rect	423	367	424	368
rect	423	368	424	369
rect	424	0	425	1
rect	424	1	425	2
rect	424	2	425	3
rect	424	3	425	4
rect	424	4	425	5
rect	424	5	425	6
rect	424	6	425	7
rect	424	7	425	8
rect	424	8	425	9
rect	424	9	425	10
rect	424	10	425	11
rect	424	11	425	12
rect	424	12	425	13
rect	424	13	425	14
rect	424	14	425	15
rect	424	15	425	16
rect	424	16	425	17
rect	424	17	425	18
rect	424	18	425	19
rect	424	19	425	20
rect	424	20	425	21
rect	424	21	425	22
rect	424	22	425	23
rect	424	23	425	24
rect	424	24	425	25
rect	424	25	425	26
rect	424	26	425	27
rect	424	27	425	28
rect	424	28	425	29
rect	424	29	425	30
rect	424	30	425	31
rect	424	31	425	32
rect	424	32	425	33
rect	424	33	425	34
rect	424	34	425	35
rect	424	35	425	36
rect	424	36	425	37
rect	424	37	425	38
rect	424	38	425	39
rect	424	39	425	40
rect	424	40	425	41
rect	424	41	425	42
rect	424	42	425	43
rect	424	43	425	44
rect	424	44	425	45
rect	424	45	425	46
rect	424	46	425	47
rect	424	47	425	48
rect	424	48	425	49
rect	424	49	425	50
rect	424	50	425	51
rect	424	51	425	52
rect	424	52	425	53
rect	424	53	425	54
rect	424	54	425	55
rect	424	55	425	56
rect	424	56	425	57
rect	424	57	425	58
rect	424	58	425	59
rect	424	59	425	60
rect	424	60	425	61
rect	424	61	425	62
rect	424	62	425	63
rect	424	63	425	64
rect	424	64	425	65
rect	424	65	425	66
rect	424	66	425	67
rect	424	67	425	68
rect	424	68	425	69
rect	424	69	425	70
rect	424	70	425	71
rect	424	71	425	72
rect	424	72	425	73
rect	424	73	425	74
rect	424	74	425	75
rect	424	75	425	76
rect	424	76	425	77
rect	424	77	425	78
rect	424	78	425	79
rect	424	79	425	80
rect	424	80	425	81
rect	424	81	425	82
rect	424	82	425	83
rect	424	83	425	84
rect	424	84	425	85
rect	424	85	425	86
rect	424	86	425	87
rect	424	87	425	88
rect	424	88	425	89
rect	424	89	425	90
rect	424	90	425	91
rect	424	91	425	92
rect	424	92	425	93
rect	424	93	425	94
rect	424	94	425	95
rect	424	95	425	96
rect	424	96	425	97
rect	424	97	425	98
rect	424	98	425	99
rect	424	99	425	100
rect	424	100	425	101
rect	424	101	425	102
rect	424	102	425	103
rect	424	103	425	104
rect	424	104	425	105
rect	424	105	425	106
rect	424	106	425	107
rect	424	107	425	108
rect	424	108	425	109
rect	424	109	425	110
rect	424	110	425	111
rect	424	111	425	112
rect	424	112	425	113
rect	424	113	425	114
rect	424	114	425	115
rect	424	115	425	116
rect	424	116	425	117
rect	424	117	425	118
rect	424	118	425	119
rect	424	119	425	120
rect	424	120	425	121
rect	424	121	425	122
rect	424	122	425	123
rect	424	123	425	124
rect	424	124	425	125
rect	424	125	425	126
rect	424	126	425	127
rect	424	127	425	128
rect	424	128	425	129
rect	424	129	425	130
rect	424	130	425	131
rect	424	131	425	132
rect	424	132	425	133
rect	424	133	425	134
rect	424	134	425	135
rect	424	135	425	136
rect	424	136	425	137
rect	424	137	425	138
rect	424	138	425	139
rect	424	139	425	140
rect	424	140	425	141
rect	424	141	425	142
rect	424	142	425	143
rect	424	143	425	144
rect	424	144	425	145
rect	424	145	425	146
rect	424	146	425	147
rect	424	147	425	148
rect	424	148	425	149
rect	424	149	425	150
rect	424	150	425	151
rect	424	151	425	152
rect	424	152	425	153
rect	424	153	425	154
rect	424	154	425	155
rect	424	155	425	156
rect	424	156	425	157
rect	424	157	425	158
rect	424	158	425	159
rect	424	159	425	160
rect	424	160	425	161
rect	424	161	425	162
rect	424	162	425	163
rect	424	163	425	164
rect	424	164	425	165
rect	424	165	425	166
rect	424	166	425	167
rect	424	167	425	168
rect	424	168	425	169
rect	424	169	425	170
rect	424	170	425	171
rect	424	171	425	172
rect	424	172	425	173
rect	424	173	425	174
rect	424	174	425	175
rect	424	175	425	176
rect	424	176	425	177
rect	424	177	425	178
rect	424	178	425	179
rect	424	179	425	180
rect	424	180	425	181
rect	424	181	425	182
rect	424	182	425	183
rect	424	183	425	184
rect	424	184	425	185
rect	424	185	425	186
rect	424	186	425	187
rect	424	187	425	188
rect	424	188	425	189
rect	424	189	425	190
rect	424	190	425	191
rect	424	191	425	192
rect	424	192	425	193
rect	424	193	425	194
rect	424	194	425	195
rect	424	195	425	196
rect	424	196	425	197
rect	424	197	425	198
rect	424	198	425	199
rect	424	199	425	200
rect	424	200	425	201
rect	424	201	425	202
rect	424	202	425	203
rect	424	203	425	204
rect	424	204	425	205
rect	424	205	425	206
rect	424	206	425	207
rect	424	207	425	208
rect	424	208	425	209
rect	424	209	425	210
rect	424	210	425	211
rect	424	211	425	212
rect	424	212	425	213
rect	424	213	425	214
rect	424	214	425	215
rect	424	215	425	216
rect	424	216	425	217
rect	424	217	425	218
rect	424	218	425	219
rect	424	219	425	220
rect	424	220	425	221
rect	424	221	425	222
rect	424	222	425	223
rect	424	223	425	224
rect	424	224	425	225
rect	424	225	425	226
rect	424	226	425	227
rect	424	227	425	228
rect	424	228	425	229
rect	424	229	425	230
rect	424	230	425	231
rect	424	231	425	232
rect	424	232	425	233
rect	424	233	425	234
rect	424	234	425	235
rect	424	235	425	236
rect	424	236	425	237
rect	424	237	425	238
rect	424	238	425	239
rect	424	239	425	240
rect	424	240	425	241
rect	424	241	425	242
rect	424	242	425	243
rect	424	243	425	244
rect	424	244	425	245
rect	424	245	425	246
rect	424	246	425	247
rect	424	247	425	248
rect	424	248	425	249
rect	424	249	425	250
rect	424	250	425	251
rect	424	251	425	252
rect	424	252	425	253
rect	424	253	425	254
rect	424	254	425	255
rect	424	255	425	256
rect	424	256	425	257
rect	424	257	425	258
rect	424	258	425	259
rect	424	259	425	260
rect	424	260	425	261
rect	424	261	425	262
rect	424	262	425	263
rect	424	263	425	264
rect	424	264	425	265
rect	424	265	425	266
rect	424	266	425	267
rect	424	267	425	268
rect	424	268	425	269
rect	424	269	425	270
rect	424	270	425	271
rect	424	271	425	272
rect	424	272	425	273
rect	424	273	425	274
rect	424	274	425	275
rect	424	275	425	276
rect	424	276	425	277
rect	424	277	425	278
rect	424	278	425	279
rect	424	279	425	280
rect	424	280	425	281
rect	424	281	425	282
rect	424	282	425	283
rect	424	283	425	284
rect	424	284	425	285
rect	424	285	425	286
rect	424	286	425	287
rect	424	287	425	288
rect	424	288	425	289
rect	424	289	425	290
rect	424	290	425	291
rect	424	291	425	292
rect	424	292	425	293
rect	424	293	425	294
rect	424	294	425	295
rect	424	295	425	296
rect	424	296	425	297
rect	424	297	425	298
rect	424	298	425	299
rect	424	299	425	300
rect	424	300	425	301
rect	424	301	425	302
rect	424	302	425	303
rect	424	303	425	304
rect	424	304	425	305
rect	424	305	425	306
rect	424	306	425	307
rect	424	307	425	308
rect	424	308	425	309
rect	424	309	425	310
rect	424	310	425	311
rect	424	311	425	312
rect	424	312	425	313
rect	424	313	425	314
rect	424	314	425	315
rect	424	315	425	316
rect	424	316	425	317
rect	424	317	425	318
rect	424	318	425	319
rect	424	319	425	320
rect	424	320	425	321
rect	424	321	425	322
rect	424	322	425	323
rect	424	323	425	324
rect	424	324	425	325
rect	424	325	425	326
rect	424	326	425	327
rect	424	327	425	328
rect	424	328	425	329
rect	424	329	425	330
rect	424	330	425	331
rect	424	331	425	332
rect	424	332	425	333
rect	424	333	425	334
rect	424	334	425	335
rect	424	335	425	336
rect	424	336	425	337
rect	424	337	425	338
rect	424	338	425	339
rect	424	339	425	340
rect	424	340	425	341
rect	424	341	425	342
rect	424	342	425	343
rect	424	343	425	344
rect	424	344	425	345
rect	424	345	425	346
rect	424	346	425	347
rect	424	347	425	348
rect	424	348	425	349
rect	424	349	425	350
rect	424	350	425	351
rect	424	351	425	352
rect	424	352	425	353
rect	424	353	425	354
rect	424	354	425	355
rect	424	355	425	356
rect	424	356	425	357
rect	424	357	425	358
rect	424	358	425	359
rect	424	359	425	360
rect	424	360	425	361
rect	424	361	425	362
rect	424	362	425	363
rect	424	363	425	364
rect	424	364	425	365
rect	424	365	425	366
rect	424	366	425	367
rect	424	367	425	368
rect	424	368	425	369
rect	425	0	426	1
rect	425	1	426	2
rect	425	2	426	3
rect	425	3	426	4
rect	425	4	426	5
rect	425	5	426	6
rect	425	6	426	7
rect	425	7	426	8
rect	425	8	426	9
rect	425	9	426	10
rect	425	10	426	11
rect	425	11	426	12
rect	425	12	426	13
rect	425	13	426	14
rect	425	14	426	15
rect	425	15	426	16
rect	425	16	426	17
rect	425	17	426	18
rect	425	18	426	19
rect	425	19	426	20
rect	425	20	426	21
rect	425	21	426	22
rect	425	22	426	23
rect	425	23	426	24
rect	425	24	426	25
rect	425	25	426	26
rect	425	26	426	27
rect	425	27	426	28
rect	425	28	426	29
rect	425	29	426	30
rect	425	30	426	31
rect	425	31	426	32
rect	425	32	426	33
rect	425	33	426	34
rect	425	34	426	35
rect	425	35	426	36
rect	425	36	426	37
rect	425	37	426	38
rect	425	38	426	39
rect	425	39	426	40
rect	425	40	426	41
rect	425	41	426	42
rect	425	42	426	43
rect	425	43	426	44
rect	425	44	426	45
rect	425	45	426	46
rect	425	46	426	47
rect	425	47	426	48
rect	425	48	426	49
rect	425	49	426	50
rect	425	50	426	51
rect	425	51	426	52
rect	425	52	426	53
rect	425	53	426	54
rect	425	54	426	55
rect	425	55	426	56
rect	425	56	426	57
rect	425	57	426	58
rect	425	58	426	59
rect	425	59	426	60
rect	425	60	426	61
rect	425	61	426	62
rect	425	62	426	63
rect	425	63	426	64
rect	425	64	426	65
rect	425	65	426	66
rect	425	66	426	67
rect	425	67	426	68
rect	425	68	426	69
rect	425	69	426	70
rect	425	70	426	71
rect	425	71	426	72
rect	425	72	426	73
rect	425	73	426	74
rect	425	74	426	75
rect	425	75	426	76
rect	425	76	426	77
rect	425	77	426	78
rect	425	78	426	79
rect	425	79	426	80
rect	425	80	426	81
rect	425	81	426	82
rect	425	82	426	83
rect	425	83	426	84
rect	425	84	426	85
rect	425	85	426	86
rect	425	86	426	87
rect	425	87	426	88
rect	425	88	426	89
rect	425	89	426	90
rect	425	90	426	91
rect	425	91	426	92
rect	425	92	426	93
rect	425	93	426	94
rect	425	94	426	95
rect	425	95	426	96
rect	425	96	426	97
rect	425	97	426	98
rect	425	98	426	99
rect	425	99	426	100
rect	425	100	426	101
rect	425	101	426	102
rect	425	102	426	103
rect	425	103	426	104
rect	425	104	426	105
rect	425	105	426	106
rect	425	106	426	107
rect	425	107	426	108
rect	425	108	426	109
rect	425	109	426	110
rect	425	110	426	111
rect	425	111	426	112
rect	425	112	426	113
rect	425	113	426	114
rect	425	114	426	115
rect	425	115	426	116
rect	425	116	426	117
rect	425	117	426	118
rect	425	118	426	119
rect	425	119	426	120
rect	425	120	426	121
rect	425	121	426	122
rect	425	122	426	123
rect	425	123	426	124
rect	425	124	426	125
rect	425	125	426	126
rect	425	126	426	127
rect	425	127	426	128
rect	425	128	426	129
rect	425	129	426	130
rect	425	130	426	131
rect	425	131	426	132
rect	425	132	426	133
rect	425	133	426	134
rect	425	134	426	135
rect	425	135	426	136
rect	425	136	426	137
rect	425	137	426	138
rect	425	138	426	139
rect	425	139	426	140
rect	425	140	426	141
rect	425	141	426	142
rect	425	142	426	143
rect	425	143	426	144
rect	425	144	426	145
rect	425	145	426	146
rect	425	146	426	147
rect	425	147	426	148
rect	425	148	426	149
rect	425	149	426	150
rect	425	150	426	151
rect	425	151	426	152
rect	425	152	426	153
rect	425	153	426	154
rect	425	154	426	155
rect	425	155	426	156
rect	425	156	426	157
rect	425	157	426	158
rect	425	158	426	159
rect	425	159	426	160
rect	425	160	426	161
rect	425	161	426	162
rect	425	162	426	163
rect	425	163	426	164
rect	425	164	426	165
rect	425	165	426	166
rect	425	166	426	167
rect	425	167	426	168
rect	425	168	426	169
rect	425	169	426	170
rect	425	170	426	171
rect	425	171	426	172
rect	425	172	426	173
rect	425	173	426	174
rect	425	174	426	175
rect	425	175	426	176
rect	425	176	426	177
rect	425	177	426	178
rect	425	178	426	179
rect	425	179	426	180
rect	425	180	426	181
rect	425	181	426	182
rect	425	182	426	183
rect	425	183	426	184
rect	425	184	426	185
rect	425	185	426	186
rect	425	186	426	187
rect	425	187	426	188
rect	425	188	426	189
rect	425	189	426	190
rect	425	190	426	191
rect	425	191	426	192
rect	425	192	426	193
rect	425	193	426	194
rect	425	194	426	195
rect	425	195	426	196
rect	425	196	426	197
rect	425	197	426	198
rect	425	198	426	199
rect	425	199	426	200
rect	425	200	426	201
rect	425	201	426	202
rect	425	202	426	203
rect	425	203	426	204
rect	425	204	426	205
rect	425	205	426	206
rect	425	206	426	207
rect	425	207	426	208
rect	425	208	426	209
rect	425	209	426	210
rect	425	210	426	211
rect	425	211	426	212
rect	425	212	426	213
rect	425	213	426	214
rect	425	214	426	215
rect	425	215	426	216
rect	425	216	426	217
rect	425	217	426	218
rect	425	218	426	219
rect	425	219	426	220
rect	425	220	426	221
rect	425	221	426	222
rect	425	222	426	223
rect	425	223	426	224
rect	425	224	426	225
rect	425	225	426	226
rect	425	226	426	227
rect	425	227	426	228
rect	425	228	426	229
rect	425	229	426	230
rect	425	230	426	231
rect	425	231	426	232
rect	425	232	426	233
rect	425	233	426	234
rect	425	234	426	235
rect	425	235	426	236
rect	425	236	426	237
rect	425	237	426	238
rect	425	238	426	239
rect	425	239	426	240
rect	425	240	426	241
rect	425	241	426	242
rect	425	242	426	243
rect	425	243	426	244
rect	425	244	426	245
rect	425	245	426	246
rect	425	246	426	247
rect	425	247	426	248
rect	425	248	426	249
rect	425	249	426	250
rect	425	250	426	251
rect	425	251	426	252
rect	425	252	426	253
rect	425	253	426	254
rect	425	254	426	255
rect	425	255	426	256
rect	425	256	426	257
rect	425	257	426	258
rect	425	258	426	259
rect	425	259	426	260
rect	425	260	426	261
rect	425	261	426	262
rect	425	262	426	263
rect	425	263	426	264
rect	425	264	426	265
rect	425	265	426	266
rect	425	266	426	267
rect	425	267	426	268
rect	425	268	426	269
rect	425	269	426	270
rect	425	270	426	271
rect	425	271	426	272
rect	425	272	426	273
rect	425	273	426	274
rect	425	274	426	275
rect	425	275	426	276
rect	425	276	426	277
rect	425	277	426	278
rect	425	278	426	279
rect	425	279	426	280
rect	425	280	426	281
rect	425	281	426	282
rect	425	282	426	283
rect	425	283	426	284
rect	425	284	426	285
rect	425	285	426	286
rect	425	286	426	287
rect	425	287	426	288
rect	425	288	426	289
rect	425	289	426	290
rect	425	290	426	291
rect	425	291	426	292
rect	425	292	426	293
rect	425	293	426	294
rect	425	294	426	295
rect	425	295	426	296
rect	425	296	426	297
rect	425	297	426	298
rect	425	298	426	299
rect	425	299	426	300
rect	425	300	426	301
rect	425	301	426	302
rect	425	302	426	303
rect	425	303	426	304
rect	425	304	426	305
rect	425	305	426	306
rect	425	306	426	307
rect	425	307	426	308
rect	425	308	426	309
rect	425	309	426	310
rect	425	310	426	311
rect	425	311	426	312
rect	425	312	426	313
rect	425	313	426	314
rect	425	314	426	315
rect	425	315	426	316
rect	425	316	426	317
rect	425	317	426	318
rect	425	318	426	319
rect	425	319	426	320
rect	425	320	426	321
rect	425	321	426	322
rect	425	322	426	323
rect	425	323	426	324
rect	425	324	426	325
rect	425	325	426	326
rect	425	326	426	327
rect	425	327	426	328
rect	425	328	426	329
rect	425	329	426	330
rect	425	330	426	331
rect	425	331	426	332
rect	425	332	426	333
rect	425	333	426	334
rect	425	334	426	335
rect	425	335	426	336
rect	425	336	426	337
rect	425	337	426	338
rect	425	338	426	339
rect	425	339	426	340
rect	425	340	426	341
rect	425	341	426	342
rect	425	342	426	343
rect	425	343	426	344
rect	425	344	426	345
rect	425	345	426	346
rect	425	346	426	347
rect	425	347	426	348
rect	425	348	426	349
rect	425	349	426	350
rect	425	350	426	351
rect	425	351	426	352
rect	425	352	426	353
rect	425	353	426	354
rect	425	354	426	355
rect	425	355	426	356
rect	425	356	426	357
rect	425	357	426	358
rect	425	358	426	359
rect	425	359	426	360
rect	425	360	426	361
rect	425	361	426	362
rect	425	362	426	363
rect	425	363	426	364
rect	425	364	426	365
rect	425	365	426	366
rect	425	366	426	367
rect	425	367	426	368
rect	425	368	426	369
rect	426	0	427	1
rect	426	1	427	2
rect	426	2	427	3
rect	426	3	427	4
rect	426	4	427	5
rect	426	5	427	6
rect	426	6	427	7
rect	426	7	427	8
rect	426	8	427	9
rect	426	9	427	10
rect	426	10	427	11
rect	426	11	427	12
rect	426	12	427	13
rect	426	13	427	14
rect	426	14	427	15
rect	426	15	427	16
rect	426	16	427	17
rect	426	17	427	18
rect	426	18	427	19
rect	426	19	427	20
rect	426	20	427	21
rect	426	21	427	22
rect	426	22	427	23
rect	426	23	427	24
rect	426	24	427	25
rect	426	25	427	26
rect	426	26	427	27
rect	426	27	427	28
rect	426	28	427	29
rect	426	29	427	30
rect	426	30	427	31
rect	426	31	427	32
rect	426	32	427	33
rect	426	33	427	34
rect	426	34	427	35
rect	426	35	427	36
rect	426	36	427	37
rect	426	37	427	38
rect	426	38	427	39
rect	426	39	427	40
rect	426	40	427	41
rect	426	41	427	42
rect	426	42	427	43
rect	426	43	427	44
rect	426	44	427	45
rect	426	45	427	46
rect	426	46	427	47
rect	426	47	427	48
rect	426	48	427	49
rect	426	49	427	50
rect	426	50	427	51
rect	426	51	427	52
rect	426	52	427	53
rect	426	53	427	54
rect	426	54	427	55
rect	426	55	427	56
rect	426	56	427	57
rect	426	57	427	58
rect	426	58	427	59
rect	426	59	427	60
rect	426	60	427	61
rect	426	61	427	62
rect	426	62	427	63
rect	426	63	427	64
rect	426	64	427	65
rect	426	65	427	66
rect	426	66	427	67
rect	426	67	427	68
rect	426	68	427	69
rect	426	69	427	70
rect	426	70	427	71
rect	426	71	427	72
rect	426	72	427	73
rect	426	73	427	74
rect	426	74	427	75
rect	426	75	427	76
rect	426	76	427	77
rect	426	77	427	78
rect	426	78	427	79
rect	426	79	427	80
rect	426	80	427	81
rect	426	81	427	82
rect	426	82	427	83
rect	426	83	427	84
rect	426	84	427	85
rect	426	85	427	86
rect	426	86	427	87
rect	426	87	427	88
rect	426	88	427	89
rect	426	89	427	90
rect	426	90	427	91
rect	426	91	427	92
rect	426	92	427	93
rect	426	93	427	94
rect	426	94	427	95
rect	426	95	427	96
rect	426	96	427	97
rect	426	97	427	98
rect	426	98	427	99
rect	426	99	427	100
rect	426	100	427	101
rect	426	101	427	102
rect	426	102	427	103
rect	426	103	427	104
rect	426	104	427	105
rect	426	105	427	106
rect	426	106	427	107
rect	426	107	427	108
rect	426	108	427	109
rect	426	109	427	110
rect	426	110	427	111
rect	426	111	427	112
rect	426	112	427	113
rect	426	113	427	114
rect	426	114	427	115
rect	426	115	427	116
rect	426	116	427	117
rect	426	117	427	118
rect	426	118	427	119
rect	426	119	427	120
rect	426	120	427	121
rect	426	121	427	122
rect	426	122	427	123
rect	426	123	427	124
rect	426	124	427	125
rect	426	125	427	126
rect	426	126	427	127
rect	426	127	427	128
rect	426	128	427	129
rect	426	129	427	130
rect	426	130	427	131
rect	426	131	427	132
rect	426	132	427	133
rect	426	133	427	134
rect	426	134	427	135
rect	426	135	427	136
rect	426	136	427	137
rect	426	137	427	138
rect	426	138	427	139
rect	426	139	427	140
rect	426	140	427	141
rect	426	141	427	142
rect	426	142	427	143
rect	426	143	427	144
rect	426	144	427	145
rect	426	145	427	146
rect	426	146	427	147
rect	426	147	427	148
rect	426	148	427	149
rect	426	149	427	150
rect	426	150	427	151
rect	426	151	427	152
rect	426	152	427	153
rect	426	153	427	154
rect	426	154	427	155
rect	426	155	427	156
rect	426	156	427	157
rect	426	157	427	158
rect	426	158	427	159
rect	426	159	427	160
rect	426	160	427	161
rect	426	161	427	162
rect	426	162	427	163
rect	426	163	427	164
rect	426	164	427	165
rect	426	165	427	166
rect	426	166	427	167
rect	426	167	427	168
rect	426	168	427	169
rect	426	169	427	170
rect	426	170	427	171
rect	426	171	427	172
rect	426	172	427	173
rect	426	173	427	174
rect	426	174	427	175
rect	426	175	427	176
rect	426	176	427	177
rect	426	177	427	178
rect	426	178	427	179
rect	426	179	427	180
rect	426	180	427	181
rect	426	181	427	182
rect	426	182	427	183
rect	426	183	427	184
rect	426	184	427	185
rect	426	185	427	186
rect	426	186	427	187
rect	426	187	427	188
rect	426	188	427	189
rect	426	189	427	190
rect	426	190	427	191
rect	426	191	427	192
rect	426	192	427	193
rect	426	193	427	194
rect	426	194	427	195
rect	426	195	427	196
rect	426	196	427	197
rect	426	197	427	198
rect	426	198	427	199
rect	426	199	427	200
rect	426	200	427	201
rect	426	201	427	202
rect	426	202	427	203
rect	426	203	427	204
rect	426	204	427	205
rect	426	205	427	206
rect	426	206	427	207
rect	426	207	427	208
rect	426	208	427	209
rect	426	209	427	210
rect	426	210	427	211
rect	426	211	427	212
rect	426	212	427	213
rect	426	213	427	214
rect	426	214	427	215
rect	426	215	427	216
rect	426	216	427	217
rect	426	217	427	218
rect	426	218	427	219
rect	426	219	427	220
rect	426	220	427	221
rect	426	221	427	222
rect	426	222	427	223
rect	426	223	427	224
rect	426	224	427	225
rect	426	225	427	226
rect	426	226	427	227
rect	426	227	427	228
rect	426	228	427	229
rect	426	229	427	230
rect	426	230	427	231
rect	426	231	427	232
rect	426	232	427	233
rect	426	233	427	234
rect	426	234	427	235
rect	426	235	427	236
rect	426	236	427	237
rect	426	237	427	238
rect	426	238	427	239
rect	426	239	427	240
rect	426	240	427	241
rect	426	241	427	242
rect	426	242	427	243
rect	426	243	427	244
rect	426	244	427	245
rect	426	245	427	246
rect	426	246	427	247
rect	426	247	427	248
rect	426	248	427	249
rect	426	249	427	250
rect	426	250	427	251
rect	426	251	427	252
rect	426	252	427	253
rect	426	253	427	254
rect	426	254	427	255
rect	426	255	427	256
rect	426	256	427	257
rect	426	257	427	258
rect	426	258	427	259
rect	426	259	427	260
rect	426	260	427	261
rect	426	261	427	262
rect	426	262	427	263
rect	426	263	427	264
rect	426	264	427	265
rect	426	265	427	266
rect	426	266	427	267
rect	426	267	427	268
rect	426	268	427	269
rect	426	269	427	270
rect	426	270	427	271
rect	426	271	427	272
rect	426	272	427	273
rect	426	273	427	274
rect	426	274	427	275
rect	426	275	427	276
rect	426	276	427	277
rect	426	277	427	278
rect	426	278	427	279
rect	426	279	427	280
rect	426	280	427	281
rect	426	281	427	282
rect	426	282	427	283
rect	426	283	427	284
rect	426	284	427	285
rect	426	285	427	286
rect	426	286	427	287
rect	426	287	427	288
rect	426	288	427	289
rect	426	289	427	290
rect	426	290	427	291
rect	426	291	427	292
rect	426	292	427	293
rect	426	293	427	294
rect	426	294	427	295
rect	426	295	427	296
rect	426	296	427	297
rect	426	297	427	298
rect	426	298	427	299
rect	426	299	427	300
rect	426	300	427	301
rect	426	301	427	302
rect	426	302	427	303
rect	426	303	427	304
rect	426	304	427	305
rect	426	305	427	306
rect	426	306	427	307
rect	426	307	427	308
rect	426	308	427	309
rect	426	309	427	310
rect	426	310	427	311
rect	426	311	427	312
rect	426	312	427	313
rect	426	313	427	314
rect	426	314	427	315
rect	426	315	427	316
rect	426	316	427	317
rect	426	317	427	318
rect	426	318	427	319
rect	426	319	427	320
rect	426	320	427	321
rect	426	321	427	322
rect	426	322	427	323
rect	426	323	427	324
rect	426	324	427	325
rect	426	325	427	326
rect	426	326	427	327
rect	426	327	427	328
rect	426	328	427	329
rect	426	329	427	330
rect	426	330	427	331
rect	426	331	427	332
rect	426	332	427	333
rect	426	333	427	334
rect	426	334	427	335
rect	426	335	427	336
rect	426	336	427	337
rect	426	337	427	338
rect	426	338	427	339
rect	426	339	427	340
rect	426	340	427	341
rect	426	341	427	342
rect	426	342	427	343
rect	426	343	427	344
rect	426	344	427	345
rect	426	345	427	346
rect	426	346	427	347
rect	426	347	427	348
rect	426	348	427	349
rect	426	349	427	350
rect	426	350	427	351
rect	426	351	427	352
rect	426	352	427	353
rect	426	353	427	354
rect	426	354	427	355
rect	426	355	427	356
rect	426	356	427	357
rect	426	357	427	358
rect	426	358	427	359
rect	426	359	427	360
rect	426	360	427	361
rect	426	361	427	362
rect	426	362	427	363
rect	426	363	427	364
rect	426	364	427	365
rect	426	365	427	366
rect	426	366	427	367
rect	426	367	427	368
rect	426	368	427	369
rect	452	0	453	1
rect	452	1	453	2
rect	452	2	453	3
rect	452	3	453	4
rect	452	4	453	5
rect	452	5	453	6
rect	452	6	453	7
rect	452	7	453	8
rect	452	8	453	9
rect	452	9	453	10
rect	452	10	453	11
rect	452	11	453	12
rect	452	12	453	13
rect	452	13	453	14
rect	452	14	453	15
rect	452	15	453	16
rect	452	16	453	17
rect	452	17	453	18
rect	452	18	453	19
rect	452	19	453	20
rect	452	20	453	21
rect	452	21	453	22
rect	452	22	453	23
rect	452	23	453	24
rect	452	24	453	25
rect	452	25	453	26
rect	452	26	453	27
rect	452	27	453	28
rect	452	28	453	29
rect	452	29	453	30
rect	452	30	453	31
rect	452	31	453	32
rect	452	32	453	33
rect	452	33	453	34
rect	452	34	453	35
rect	452	35	453	36
rect	452	36	453	37
rect	452	37	453	38
rect	452	38	453	39
rect	452	39	453	40
rect	452	40	453	41
rect	452	41	453	42
rect	452	42	453	43
rect	452	43	453	44
rect	452	44	453	45
rect	452	45	453	46
rect	452	46	453	47
rect	452	47	453	48
rect	452	48	453	49
rect	452	49	453	50
rect	452	50	453	51
rect	452	51	453	52
rect	452	52	453	53
rect	452	53	453	54
rect	452	54	453	55
rect	452	55	453	56
rect	452	56	453	57
rect	452	57	453	58
rect	452	58	453	59
rect	452	59	453	60
rect	452	60	453	61
rect	452	61	453	62
rect	452	62	453	63
rect	452	63	453	64
rect	452	64	453	65
rect	452	65	453	66
rect	452	66	453	67
rect	452	67	453	68
rect	452	68	453	69
rect	452	69	453	70
rect	452	70	453	71
rect	452	71	453	72
rect	452	72	453	73
rect	452	73	453	74
rect	452	74	453	75
rect	452	75	453	76
rect	452	76	453	77
rect	452	77	453	78
rect	452	78	453	79
rect	452	79	453	80
rect	452	80	453	81
rect	452	81	453	82
rect	452	82	453	83
rect	452	83	453	84
rect	452	84	453	85
rect	452	85	453	86
rect	452	86	453	87
rect	452	87	453	88
rect	452	88	453	89
rect	452	89	453	90
rect	452	90	453	91
rect	452	91	453	92
rect	452	92	453	93
rect	452	93	453	94
rect	452	94	453	95
rect	452	95	453	96
rect	452	96	453	97
rect	452	97	453	98
rect	452	98	453	99
rect	452	99	453	100
rect	452	100	453	101
rect	452	101	453	102
rect	452	102	453	103
rect	452	103	453	104
rect	452	104	453	105
rect	452	105	453	106
rect	452	106	453	107
rect	452	107	453	108
rect	452	108	453	109
rect	452	109	453	110
rect	452	110	453	111
rect	452	111	453	112
rect	452	112	453	113
rect	452	113	453	114
rect	452	114	453	115
rect	452	115	453	116
rect	452	116	453	117
rect	452	117	453	118
rect	452	118	453	119
rect	452	119	453	120
rect	452	120	453	121
rect	452	121	453	122
rect	452	122	453	123
rect	452	123	453	124
rect	452	124	453	125
rect	452	125	453	126
rect	452	126	453	127
rect	452	127	453	128
rect	452	128	453	129
rect	452	129	453	130
rect	452	130	453	131
rect	452	131	453	132
rect	452	132	453	133
rect	452	133	453	134
rect	452	134	453	135
rect	452	135	453	136
rect	452	136	453	137
rect	452	137	453	138
rect	452	138	453	139
rect	452	139	453	140
rect	452	140	453	141
rect	452	141	453	142
rect	452	142	453	143
rect	452	143	453	144
rect	452	144	453	145
rect	452	145	453	146
rect	452	146	453	147
rect	452	147	453	148
rect	452	148	453	149
rect	452	149	453	150
rect	452	150	453	151
rect	452	151	453	152
rect	452	152	453	153
rect	452	153	453	154
rect	452	154	453	155
rect	452	155	453	156
rect	452	156	453	157
rect	452	157	453	158
rect	452	158	453	159
rect	452	159	453	160
rect	452	160	453	161
rect	452	161	453	162
rect	452	162	453	163
rect	452	163	453	164
rect	452	164	453	165
rect	452	165	453	166
rect	452	166	453	167
rect	452	167	453	168
rect	452	168	453	169
rect	452	169	453	170
rect	452	170	453	171
rect	452	171	453	172
rect	452	172	453	173
rect	452	173	453	174
rect	452	174	453	175
rect	452	175	453	176
rect	452	176	453	177
rect	452	177	453	178
rect	452	178	453	179
rect	452	179	453	180
rect	452	180	453	181
rect	452	181	453	182
rect	452	182	453	183
rect	452	183	453	184
rect	452	184	453	185
rect	452	185	453	186
rect	452	186	453	187
rect	452	187	453	188
rect	452	188	453	189
rect	452	189	453	190
rect	452	190	453	191
rect	452	191	453	192
rect	452	192	453	193
rect	452	193	453	194
rect	452	194	453	195
rect	452	195	453	196
rect	452	196	453	197
rect	452	197	453	198
rect	452	198	453	199
rect	452	199	453	200
rect	452	200	453	201
rect	452	201	453	202
rect	452	202	453	203
rect	452	203	453	204
rect	452	204	453	205
rect	452	205	453	206
rect	452	206	453	207
rect	452	207	453	208
rect	452	208	453	209
rect	452	209	453	210
rect	452	210	453	211
rect	452	211	453	212
rect	452	212	453	213
rect	452	213	453	214
rect	452	214	453	215
rect	452	215	453	216
rect	452	216	453	217
rect	452	217	453	218
rect	452	218	453	219
rect	452	219	453	220
rect	452	220	453	221
rect	452	221	453	222
rect	452	222	453	223
rect	452	223	453	224
rect	452	224	453	225
rect	452	225	453	226
rect	452	226	453	227
rect	452	227	453	228
rect	452	228	453	229
rect	452	229	453	230
rect	452	230	453	231
rect	452	231	453	232
rect	452	232	453	233
rect	452	233	453	234
rect	452	234	453	235
rect	452	235	453	236
rect	452	236	453	237
rect	452	237	453	238
rect	452	238	453	239
rect	452	239	453	240
rect	452	240	453	241
rect	452	241	453	242
rect	452	242	453	243
rect	452	243	453	244
rect	452	244	453	245
rect	452	245	453	246
rect	452	246	453	247
rect	452	247	453	248
rect	452	248	453	249
rect	452	249	453	250
rect	452	250	453	251
rect	452	251	453	252
rect	452	252	453	253
rect	452	253	453	254
rect	452	254	453	255
rect	452	255	453	256
rect	452	256	453	257
rect	452	257	453	258
rect	452	258	453	259
rect	452	259	453	260
rect	452	260	453	261
rect	452	261	453	262
rect	452	262	453	263
rect	452	263	453	264
rect	452	264	453	265
rect	452	265	453	266
rect	452	266	453	267
rect	452	267	453	268
rect	452	268	453	269
rect	452	269	453	270
rect	452	270	453	271
rect	452	271	453	272
rect	452	272	453	273
rect	452	273	453	274
rect	452	274	453	275
rect	452	275	453	276
rect	452	276	453	277
rect	452	277	453	278
rect	452	278	453	279
rect	452	279	453	280
rect	452	280	453	281
rect	452	281	453	282
rect	452	282	453	283
rect	452	283	453	284
rect	452	284	453	285
rect	452	285	453	286
rect	452	286	453	287
rect	452	287	453	288
rect	452	288	453	289
rect	452	289	453	290
rect	452	290	453	291
rect	452	291	453	292
rect	452	292	453	293
rect	452	293	453	294
rect	452	294	453	295
rect	452	295	453	296
rect	452	296	453	297
rect	452	297	453	298
rect	452	298	453	299
rect	452	299	453	300
rect	452	300	453	301
rect	452	301	453	302
rect	452	302	453	303
rect	452	303	453	304
rect	452	304	453	305
rect	452	305	453	306
rect	452	306	453	307
rect	452	307	453	308
rect	452	308	453	309
rect	452	309	453	310
rect	452	310	453	311
rect	452	311	453	312
rect	452	312	453	313
rect	452	313	453	314
rect	452	314	453	315
rect	452	315	453	316
rect	452	316	453	317
rect	452	317	453	318
rect	452	318	453	319
rect	452	319	453	320
rect	452	320	453	321
rect	452	321	453	322
rect	452	322	453	323
rect	452	323	453	324
rect	452	324	453	325
rect	452	325	453	326
rect	452	326	453	327
rect	452	327	453	328
rect	452	328	453	329
rect	452	329	453	330
rect	452	330	453	331
rect	452	331	453	332
rect	452	332	453	333
rect	452	333	453	334
rect	452	334	453	335
rect	452	335	453	336
rect	452	336	453	337
rect	452	337	453	338
rect	452	338	453	339
rect	452	339	453	340
rect	452	340	453	341
rect	452	341	453	342
rect	452	342	453	343
rect	452	343	453	344
rect	452	344	453	345
rect	452	345	453	346
rect	452	346	453	347
rect	452	347	453	348
rect	453	0	454	1
rect	453	1	454	2
rect	453	2	454	3
rect	453	3	454	4
rect	453	4	454	5
rect	453	5	454	6
rect	453	6	454	7
rect	453	7	454	8
rect	453	8	454	9
rect	453	9	454	10
rect	453	10	454	11
rect	453	11	454	12
rect	453	12	454	13
rect	453	13	454	14
rect	453	14	454	15
rect	453	15	454	16
rect	453	16	454	17
rect	453	17	454	18
rect	453	18	454	19
rect	453	19	454	20
rect	453	20	454	21
rect	453	21	454	22
rect	453	22	454	23
rect	453	23	454	24
rect	453	24	454	25
rect	453	25	454	26
rect	453	26	454	27
rect	453	27	454	28
rect	453	28	454	29
rect	453	29	454	30
rect	453	30	454	31
rect	453	31	454	32
rect	453	32	454	33
rect	453	33	454	34
rect	453	34	454	35
rect	453	35	454	36
rect	453	36	454	37
rect	453	37	454	38
rect	453	38	454	39
rect	453	39	454	40
rect	453	40	454	41
rect	453	41	454	42
rect	453	42	454	43
rect	453	43	454	44
rect	453	44	454	45
rect	453	45	454	46
rect	453	46	454	47
rect	453	47	454	48
rect	453	48	454	49
rect	453	49	454	50
rect	453	50	454	51
rect	453	51	454	52
rect	453	52	454	53
rect	453	53	454	54
rect	453	54	454	55
rect	453	55	454	56
rect	453	56	454	57
rect	453	57	454	58
rect	453	58	454	59
rect	453	59	454	60
rect	453	60	454	61
rect	453	61	454	62
rect	453	62	454	63
rect	453	63	454	64
rect	453	64	454	65
rect	453	65	454	66
rect	453	66	454	67
rect	453	67	454	68
rect	453	68	454	69
rect	453	69	454	70
rect	453	70	454	71
rect	453	71	454	72
rect	453	72	454	73
rect	453	73	454	74
rect	453	74	454	75
rect	453	75	454	76
rect	453	76	454	77
rect	453	77	454	78
rect	453	78	454	79
rect	453	79	454	80
rect	453	80	454	81
rect	453	81	454	82
rect	453	82	454	83
rect	453	83	454	84
rect	453	84	454	85
rect	453	85	454	86
rect	453	86	454	87
rect	453	87	454	88
rect	453	88	454	89
rect	453	89	454	90
rect	453	90	454	91
rect	453	91	454	92
rect	453	92	454	93
rect	453	93	454	94
rect	453	94	454	95
rect	453	95	454	96
rect	453	96	454	97
rect	453	97	454	98
rect	453	98	454	99
rect	453	99	454	100
rect	453	100	454	101
rect	453	101	454	102
rect	453	102	454	103
rect	453	103	454	104
rect	453	104	454	105
rect	453	105	454	106
rect	453	106	454	107
rect	453	107	454	108
rect	453	108	454	109
rect	453	109	454	110
rect	453	110	454	111
rect	453	111	454	112
rect	453	112	454	113
rect	453	113	454	114
rect	453	114	454	115
rect	453	115	454	116
rect	453	116	454	117
rect	453	117	454	118
rect	453	118	454	119
rect	453	119	454	120
rect	453	120	454	121
rect	453	121	454	122
rect	453	122	454	123
rect	453	123	454	124
rect	453	124	454	125
rect	453	125	454	126
rect	453	126	454	127
rect	453	127	454	128
rect	453	128	454	129
rect	453	129	454	130
rect	453	130	454	131
rect	453	131	454	132
rect	453	132	454	133
rect	453	133	454	134
rect	453	134	454	135
rect	453	135	454	136
rect	453	136	454	137
rect	453	137	454	138
rect	453	138	454	139
rect	453	139	454	140
rect	453	140	454	141
rect	453	141	454	142
rect	453	142	454	143
rect	453	143	454	144
rect	453	144	454	145
rect	453	145	454	146
rect	453	146	454	147
rect	453	147	454	148
rect	453	148	454	149
rect	453	149	454	150
rect	453	150	454	151
rect	453	151	454	152
rect	453	152	454	153
rect	453	153	454	154
rect	453	154	454	155
rect	453	155	454	156
rect	453	156	454	157
rect	453	157	454	158
rect	453	158	454	159
rect	453	159	454	160
rect	453	160	454	161
rect	453	161	454	162
rect	453	162	454	163
rect	453	163	454	164
rect	453	164	454	165
rect	453	165	454	166
rect	453	166	454	167
rect	453	167	454	168
rect	453	168	454	169
rect	453	169	454	170
rect	453	170	454	171
rect	453	171	454	172
rect	453	172	454	173
rect	453	173	454	174
rect	453	174	454	175
rect	453	175	454	176
rect	453	176	454	177
rect	453	177	454	178
rect	453	178	454	179
rect	453	179	454	180
rect	453	180	454	181
rect	453	181	454	182
rect	453	182	454	183
rect	453	183	454	184
rect	453	184	454	185
rect	453	185	454	186
rect	453	186	454	187
rect	453	187	454	188
rect	453	188	454	189
rect	453	189	454	190
rect	453	190	454	191
rect	453	191	454	192
rect	453	192	454	193
rect	453	193	454	194
rect	453	194	454	195
rect	453	195	454	196
rect	453	196	454	197
rect	453	197	454	198
rect	453	198	454	199
rect	453	199	454	200
rect	453	200	454	201
rect	453	201	454	202
rect	453	202	454	203
rect	453	203	454	204
rect	453	204	454	205
rect	453	205	454	206
rect	453	206	454	207
rect	453	207	454	208
rect	453	208	454	209
rect	453	209	454	210
rect	453	210	454	211
rect	453	211	454	212
rect	453	212	454	213
rect	453	213	454	214
rect	453	214	454	215
rect	453	215	454	216
rect	453	216	454	217
rect	453	217	454	218
rect	453	218	454	219
rect	453	219	454	220
rect	453	220	454	221
rect	453	221	454	222
rect	453	222	454	223
rect	453	223	454	224
rect	453	224	454	225
rect	453	225	454	226
rect	453	226	454	227
rect	453	227	454	228
rect	453	228	454	229
rect	453	229	454	230
rect	453	230	454	231
rect	453	231	454	232
rect	453	232	454	233
rect	453	233	454	234
rect	453	234	454	235
rect	453	235	454	236
rect	453	236	454	237
rect	453	237	454	238
rect	453	238	454	239
rect	453	239	454	240
rect	453	240	454	241
rect	453	241	454	242
rect	453	242	454	243
rect	453	243	454	244
rect	453	244	454	245
rect	453	245	454	246
rect	453	246	454	247
rect	453	247	454	248
rect	453	248	454	249
rect	453	249	454	250
rect	453	250	454	251
rect	453	251	454	252
rect	453	252	454	253
rect	453	253	454	254
rect	453	254	454	255
rect	453	255	454	256
rect	453	256	454	257
rect	453	257	454	258
rect	453	258	454	259
rect	453	259	454	260
rect	453	260	454	261
rect	453	261	454	262
rect	453	262	454	263
rect	453	263	454	264
rect	453	264	454	265
rect	453	265	454	266
rect	453	266	454	267
rect	453	267	454	268
rect	453	268	454	269
rect	453	269	454	270
rect	453	270	454	271
rect	453	271	454	272
rect	453	272	454	273
rect	453	273	454	274
rect	453	274	454	275
rect	453	275	454	276
rect	453	276	454	277
rect	453	277	454	278
rect	453	278	454	279
rect	453	279	454	280
rect	453	280	454	281
rect	453	281	454	282
rect	453	282	454	283
rect	453	283	454	284
rect	453	284	454	285
rect	453	285	454	286
rect	453	286	454	287
rect	453	287	454	288
rect	453	288	454	289
rect	453	289	454	290
rect	453	290	454	291
rect	453	291	454	292
rect	453	292	454	293
rect	453	293	454	294
rect	453	294	454	295
rect	453	295	454	296
rect	453	296	454	297
rect	453	297	454	298
rect	453	298	454	299
rect	453	299	454	300
rect	453	300	454	301
rect	453	301	454	302
rect	453	302	454	303
rect	453	303	454	304
rect	453	304	454	305
rect	453	305	454	306
rect	453	306	454	307
rect	453	307	454	308
rect	453	308	454	309
rect	453	309	454	310
rect	453	310	454	311
rect	453	311	454	312
rect	453	312	454	313
rect	453	313	454	314
rect	453	314	454	315
rect	453	315	454	316
rect	453	316	454	317
rect	453	317	454	318
rect	453	318	454	319
rect	453	319	454	320
rect	453	320	454	321
rect	453	321	454	322
rect	453	322	454	323
rect	453	323	454	324
rect	453	324	454	325
rect	453	325	454	326
rect	453	326	454	327
rect	453	327	454	328
rect	453	328	454	329
rect	453	329	454	330
rect	453	330	454	331
rect	453	331	454	332
rect	453	332	454	333
rect	453	333	454	334
rect	453	334	454	335
rect	453	335	454	336
rect	453	336	454	337
rect	453	337	454	338
rect	453	338	454	339
rect	453	339	454	340
rect	453	340	454	341
rect	453	341	454	342
rect	453	342	454	343
rect	453	343	454	344
rect	453	344	454	345
rect	453	345	454	346
rect	453	346	454	347
rect	453	347	454	348
rect	454	0	455	1
rect	454	1	455	2
rect	454	2	455	3
rect	454	3	455	4
rect	454	4	455	5
rect	454	5	455	6
rect	454	6	455	7
rect	454	7	455	8
rect	454	8	455	9
rect	454	9	455	10
rect	454	10	455	11
rect	454	11	455	12
rect	454	12	455	13
rect	454	13	455	14
rect	454	14	455	15
rect	454	15	455	16
rect	454	16	455	17
rect	454	17	455	18
rect	454	18	455	19
rect	454	19	455	20
rect	454	20	455	21
rect	454	21	455	22
rect	454	22	455	23
rect	454	23	455	24
rect	454	24	455	25
rect	454	25	455	26
rect	454	26	455	27
rect	454	27	455	28
rect	454	28	455	29
rect	454	29	455	30
rect	454	30	455	31
rect	454	31	455	32
rect	454	32	455	33
rect	454	33	455	34
rect	454	34	455	35
rect	454	35	455	36
rect	454	36	455	37
rect	454	37	455	38
rect	454	38	455	39
rect	454	39	455	40
rect	454	40	455	41
rect	454	41	455	42
rect	454	42	455	43
rect	454	43	455	44
rect	454	44	455	45
rect	454	45	455	46
rect	454	46	455	47
rect	454	47	455	48
rect	454	48	455	49
rect	454	49	455	50
rect	454	50	455	51
rect	454	51	455	52
rect	454	52	455	53
rect	454	53	455	54
rect	454	54	455	55
rect	454	55	455	56
rect	454	56	455	57
rect	454	57	455	58
rect	454	58	455	59
rect	454	59	455	60
rect	454	60	455	61
rect	454	61	455	62
rect	454	62	455	63
rect	454	63	455	64
rect	454	64	455	65
rect	454	65	455	66
rect	454	66	455	67
rect	454	67	455	68
rect	454	68	455	69
rect	454	69	455	70
rect	454	70	455	71
rect	454	71	455	72
rect	454	72	455	73
rect	454	73	455	74
rect	454	74	455	75
rect	454	75	455	76
rect	454	76	455	77
rect	454	77	455	78
rect	454	78	455	79
rect	454	79	455	80
rect	454	80	455	81
rect	454	81	455	82
rect	454	82	455	83
rect	454	83	455	84
rect	454	84	455	85
rect	454	85	455	86
rect	454	86	455	87
rect	454	87	455	88
rect	454	88	455	89
rect	454	89	455	90
rect	454	90	455	91
rect	454	91	455	92
rect	454	92	455	93
rect	454	93	455	94
rect	454	94	455	95
rect	454	95	455	96
rect	454	96	455	97
rect	454	97	455	98
rect	454	98	455	99
rect	454	99	455	100
rect	454	100	455	101
rect	454	101	455	102
rect	454	102	455	103
rect	454	103	455	104
rect	454	104	455	105
rect	454	105	455	106
rect	454	106	455	107
rect	454	107	455	108
rect	454	108	455	109
rect	454	109	455	110
rect	454	110	455	111
rect	454	111	455	112
rect	454	112	455	113
rect	454	113	455	114
rect	454	114	455	115
rect	454	115	455	116
rect	454	116	455	117
rect	454	117	455	118
rect	454	118	455	119
rect	454	119	455	120
rect	454	120	455	121
rect	454	121	455	122
rect	454	122	455	123
rect	454	123	455	124
rect	454	124	455	125
rect	454	125	455	126
rect	454	126	455	127
rect	454	127	455	128
rect	454	128	455	129
rect	454	129	455	130
rect	454	130	455	131
rect	454	131	455	132
rect	454	132	455	133
rect	454	133	455	134
rect	454	134	455	135
rect	454	135	455	136
rect	454	136	455	137
rect	454	137	455	138
rect	454	138	455	139
rect	454	139	455	140
rect	454	140	455	141
rect	454	141	455	142
rect	454	142	455	143
rect	454	143	455	144
rect	454	144	455	145
rect	454	145	455	146
rect	454	146	455	147
rect	454	147	455	148
rect	454	148	455	149
rect	454	149	455	150
rect	454	150	455	151
rect	454	151	455	152
rect	454	152	455	153
rect	454	153	455	154
rect	454	154	455	155
rect	454	155	455	156
rect	454	156	455	157
rect	454	157	455	158
rect	454	158	455	159
rect	454	159	455	160
rect	454	160	455	161
rect	454	161	455	162
rect	454	162	455	163
rect	454	163	455	164
rect	454	164	455	165
rect	454	165	455	166
rect	454	166	455	167
rect	454	167	455	168
rect	454	168	455	169
rect	454	169	455	170
rect	454	170	455	171
rect	454	171	455	172
rect	454	172	455	173
rect	454	173	455	174
rect	454	174	455	175
rect	454	175	455	176
rect	454	176	455	177
rect	454	177	455	178
rect	454	178	455	179
rect	454	179	455	180
rect	454	180	455	181
rect	454	181	455	182
rect	454	182	455	183
rect	454	183	455	184
rect	454	184	455	185
rect	454	185	455	186
rect	454	186	455	187
rect	454	187	455	188
rect	454	188	455	189
rect	454	189	455	190
rect	454	190	455	191
rect	454	191	455	192
rect	454	192	455	193
rect	454	193	455	194
rect	454	194	455	195
rect	454	195	455	196
rect	454	196	455	197
rect	454	197	455	198
rect	454	198	455	199
rect	454	199	455	200
rect	454	200	455	201
rect	454	201	455	202
rect	454	202	455	203
rect	454	203	455	204
rect	454	204	455	205
rect	454	205	455	206
rect	454	206	455	207
rect	454	207	455	208
rect	454	208	455	209
rect	454	209	455	210
rect	454	210	455	211
rect	454	211	455	212
rect	454	212	455	213
rect	454	213	455	214
rect	454	214	455	215
rect	454	215	455	216
rect	454	216	455	217
rect	454	217	455	218
rect	454	218	455	219
rect	454	219	455	220
rect	454	220	455	221
rect	454	221	455	222
rect	454	222	455	223
rect	454	223	455	224
rect	454	224	455	225
rect	454	225	455	226
rect	454	226	455	227
rect	454	227	455	228
rect	454	228	455	229
rect	454	229	455	230
rect	454	230	455	231
rect	454	231	455	232
rect	454	232	455	233
rect	454	233	455	234
rect	454	234	455	235
rect	454	235	455	236
rect	454	236	455	237
rect	454	237	455	238
rect	454	238	455	239
rect	454	239	455	240
rect	454	240	455	241
rect	454	241	455	242
rect	454	242	455	243
rect	454	243	455	244
rect	454	244	455	245
rect	454	245	455	246
rect	454	246	455	247
rect	454	247	455	248
rect	454	248	455	249
rect	454	249	455	250
rect	454	250	455	251
rect	454	251	455	252
rect	454	252	455	253
rect	454	253	455	254
rect	454	254	455	255
rect	454	255	455	256
rect	454	256	455	257
rect	454	257	455	258
rect	454	258	455	259
rect	454	259	455	260
rect	454	260	455	261
rect	454	261	455	262
rect	454	262	455	263
rect	454	263	455	264
rect	454	264	455	265
rect	454	265	455	266
rect	454	266	455	267
rect	454	267	455	268
rect	454	268	455	269
rect	454	269	455	270
rect	454	270	455	271
rect	454	271	455	272
rect	454	272	455	273
rect	454	273	455	274
rect	454	274	455	275
rect	454	275	455	276
rect	454	276	455	277
rect	454	277	455	278
rect	454	278	455	279
rect	454	279	455	280
rect	454	280	455	281
rect	454	281	455	282
rect	454	282	455	283
rect	454	283	455	284
rect	454	284	455	285
rect	454	285	455	286
rect	454	286	455	287
rect	454	287	455	288
rect	454	288	455	289
rect	454	289	455	290
rect	454	290	455	291
rect	454	291	455	292
rect	454	292	455	293
rect	454	293	455	294
rect	454	294	455	295
rect	454	295	455	296
rect	454	296	455	297
rect	454	297	455	298
rect	454	298	455	299
rect	454	299	455	300
rect	454	300	455	301
rect	454	301	455	302
rect	454	302	455	303
rect	454	303	455	304
rect	454	304	455	305
rect	454	305	455	306
rect	454	306	455	307
rect	454	307	455	308
rect	454	308	455	309
rect	454	309	455	310
rect	454	310	455	311
rect	454	311	455	312
rect	454	312	455	313
rect	454	313	455	314
rect	454	314	455	315
rect	454	315	455	316
rect	454	316	455	317
rect	454	317	455	318
rect	454	318	455	319
rect	454	319	455	320
rect	454	320	455	321
rect	454	321	455	322
rect	454	322	455	323
rect	454	323	455	324
rect	454	324	455	325
rect	454	325	455	326
rect	454	326	455	327
rect	454	327	455	328
rect	454	328	455	329
rect	454	329	455	330
rect	454	330	455	331
rect	454	331	455	332
rect	454	332	455	333
rect	454	333	455	334
rect	454	334	455	335
rect	454	335	455	336
rect	454	336	455	337
rect	454	337	455	338
rect	454	338	455	339
rect	454	339	455	340
rect	454	340	455	341
rect	454	341	455	342
rect	454	342	455	343
rect	454	343	455	344
rect	454	344	455	345
rect	454	345	455	346
rect	454	346	455	347
rect	454	347	455	348
rect	455	0	456	1
rect	455	1	456	2
rect	455	2	456	3
rect	455	3	456	4
rect	455	4	456	5
rect	455	5	456	6
rect	455	6	456	7
rect	455	7	456	8
rect	455	8	456	9
rect	455	9	456	10
rect	455	10	456	11
rect	455	11	456	12
rect	455	12	456	13
rect	455	13	456	14
rect	455	14	456	15
rect	455	15	456	16
rect	455	16	456	17
rect	455	17	456	18
rect	455	18	456	19
rect	455	19	456	20
rect	455	20	456	21
rect	455	21	456	22
rect	455	22	456	23
rect	455	23	456	24
rect	455	24	456	25
rect	455	25	456	26
rect	455	26	456	27
rect	455	27	456	28
rect	455	28	456	29
rect	455	29	456	30
rect	455	30	456	31
rect	455	31	456	32
rect	455	32	456	33
rect	455	33	456	34
rect	455	34	456	35
rect	455	35	456	36
rect	455	36	456	37
rect	455	37	456	38
rect	455	38	456	39
rect	455	39	456	40
rect	455	40	456	41
rect	455	41	456	42
rect	455	42	456	43
rect	455	43	456	44
rect	455	44	456	45
rect	455	45	456	46
rect	455	46	456	47
rect	455	47	456	48
rect	455	48	456	49
rect	455	49	456	50
rect	455	50	456	51
rect	455	51	456	52
rect	455	52	456	53
rect	455	53	456	54
rect	455	54	456	55
rect	455	55	456	56
rect	455	56	456	57
rect	455	57	456	58
rect	455	58	456	59
rect	455	59	456	60
rect	455	60	456	61
rect	455	61	456	62
rect	455	62	456	63
rect	455	63	456	64
rect	455	64	456	65
rect	455	65	456	66
rect	455	66	456	67
rect	455	67	456	68
rect	455	68	456	69
rect	455	69	456	70
rect	455	70	456	71
rect	455	71	456	72
rect	455	72	456	73
rect	455	73	456	74
rect	455	74	456	75
rect	455	75	456	76
rect	455	76	456	77
rect	455	77	456	78
rect	455	78	456	79
rect	455	79	456	80
rect	455	80	456	81
rect	455	81	456	82
rect	455	82	456	83
rect	455	83	456	84
rect	455	84	456	85
rect	455	85	456	86
rect	455	86	456	87
rect	455	87	456	88
rect	455	88	456	89
rect	455	89	456	90
rect	455	90	456	91
rect	455	91	456	92
rect	455	92	456	93
rect	455	93	456	94
rect	455	94	456	95
rect	455	95	456	96
rect	455	96	456	97
rect	455	97	456	98
rect	455	98	456	99
rect	455	99	456	100
rect	455	100	456	101
rect	455	101	456	102
rect	455	102	456	103
rect	455	103	456	104
rect	455	104	456	105
rect	455	105	456	106
rect	455	106	456	107
rect	455	107	456	108
rect	455	108	456	109
rect	455	109	456	110
rect	455	110	456	111
rect	455	111	456	112
rect	455	112	456	113
rect	455	113	456	114
rect	455	114	456	115
rect	455	115	456	116
rect	455	116	456	117
rect	455	117	456	118
rect	455	118	456	119
rect	455	119	456	120
rect	455	120	456	121
rect	455	121	456	122
rect	455	122	456	123
rect	455	123	456	124
rect	455	124	456	125
rect	455	125	456	126
rect	455	126	456	127
rect	455	127	456	128
rect	455	128	456	129
rect	455	129	456	130
rect	455	130	456	131
rect	455	131	456	132
rect	455	132	456	133
rect	455	133	456	134
rect	455	134	456	135
rect	455	135	456	136
rect	455	136	456	137
rect	455	137	456	138
rect	455	138	456	139
rect	455	139	456	140
rect	455	140	456	141
rect	455	141	456	142
rect	455	142	456	143
rect	455	143	456	144
rect	455	144	456	145
rect	455	145	456	146
rect	455	146	456	147
rect	455	147	456	148
rect	455	148	456	149
rect	455	149	456	150
rect	455	150	456	151
rect	455	151	456	152
rect	455	152	456	153
rect	455	153	456	154
rect	455	154	456	155
rect	455	155	456	156
rect	455	156	456	157
rect	455	157	456	158
rect	455	158	456	159
rect	455	159	456	160
rect	455	160	456	161
rect	455	161	456	162
rect	455	162	456	163
rect	455	163	456	164
rect	455	164	456	165
rect	455	165	456	166
rect	455	166	456	167
rect	455	167	456	168
rect	455	168	456	169
rect	455	169	456	170
rect	455	170	456	171
rect	455	171	456	172
rect	455	172	456	173
rect	455	173	456	174
rect	455	174	456	175
rect	455	175	456	176
rect	455	176	456	177
rect	455	177	456	178
rect	455	178	456	179
rect	455	179	456	180
rect	455	180	456	181
rect	455	181	456	182
rect	455	182	456	183
rect	455	183	456	184
rect	455	184	456	185
rect	455	185	456	186
rect	455	186	456	187
rect	455	187	456	188
rect	455	188	456	189
rect	455	189	456	190
rect	455	190	456	191
rect	455	191	456	192
rect	455	192	456	193
rect	455	193	456	194
rect	455	194	456	195
rect	455	195	456	196
rect	455	196	456	197
rect	455	197	456	198
rect	455	198	456	199
rect	455	199	456	200
rect	455	200	456	201
rect	455	201	456	202
rect	455	202	456	203
rect	455	203	456	204
rect	455	204	456	205
rect	455	205	456	206
rect	455	206	456	207
rect	455	207	456	208
rect	455	208	456	209
rect	455	209	456	210
rect	455	210	456	211
rect	455	211	456	212
rect	455	212	456	213
rect	455	213	456	214
rect	455	214	456	215
rect	455	215	456	216
rect	455	216	456	217
rect	455	217	456	218
rect	455	218	456	219
rect	455	219	456	220
rect	455	220	456	221
rect	455	221	456	222
rect	455	222	456	223
rect	455	223	456	224
rect	455	224	456	225
rect	455	225	456	226
rect	455	226	456	227
rect	455	227	456	228
rect	455	228	456	229
rect	455	229	456	230
rect	455	230	456	231
rect	455	231	456	232
rect	455	232	456	233
rect	455	233	456	234
rect	455	234	456	235
rect	455	235	456	236
rect	455	236	456	237
rect	455	237	456	238
rect	455	238	456	239
rect	455	239	456	240
rect	455	240	456	241
rect	455	241	456	242
rect	455	242	456	243
rect	455	243	456	244
rect	455	244	456	245
rect	455	245	456	246
rect	455	246	456	247
rect	455	247	456	248
rect	455	248	456	249
rect	455	249	456	250
rect	455	250	456	251
rect	455	251	456	252
rect	455	252	456	253
rect	455	253	456	254
rect	455	254	456	255
rect	455	255	456	256
rect	455	256	456	257
rect	455	257	456	258
rect	455	258	456	259
rect	455	259	456	260
rect	455	260	456	261
rect	455	261	456	262
rect	455	262	456	263
rect	455	263	456	264
rect	455	264	456	265
rect	455	265	456	266
rect	455	266	456	267
rect	455	267	456	268
rect	455	268	456	269
rect	455	269	456	270
rect	455	270	456	271
rect	455	271	456	272
rect	455	272	456	273
rect	455	273	456	274
rect	455	274	456	275
rect	455	275	456	276
rect	455	276	456	277
rect	455	277	456	278
rect	455	278	456	279
rect	455	279	456	280
rect	455	280	456	281
rect	455	281	456	282
rect	455	282	456	283
rect	455	283	456	284
rect	455	284	456	285
rect	455	285	456	286
rect	455	286	456	287
rect	455	287	456	288
rect	455	288	456	289
rect	455	289	456	290
rect	455	290	456	291
rect	455	291	456	292
rect	455	292	456	293
rect	455	293	456	294
rect	455	294	456	295
rect	455	295	456	296
rect	455	296	456	297
rect	455	297	456	298
rect	455	298	456	299
rect	455	299	456	300
rect	455	300	456	301
rect	455	301	456	302
rect	455	302	456	303
rect	455	303	456	304
rect	455	304	456	305
rect	455	305	456	306
rect	455	306	456	307
rect	455	307	456	308
rect	455	308	456	309
rect	455	309	456	310
rect	455	310	456	311
rect	455	311	456	312
rect	455	312	456	313
rect	455	313	456	314
rect	455	314	456	315
rect	455	315	456	316
rect	455	316	456	317
rect	455	317	456	318
rect	455	318	456	319
rect	455	319	456	320
rect	455	320	456	321
rect	455	321	456	322
rect	455	322	456	323
rect	455	323	456	324
rect	455	324	456	325
rect	455	325	456	326
rect	455	326	456	327
rect	455	327	456	328
rect	455	328	456	329
rect	455	329	456	330
rect	455	330	456	331
rect	455	331	456	332
rect	455	332	456	333
rect	455	333	456	334
rect	455	334	456	335
rect	455	335	456	336
rect	455	336	456	337
rect	455	337	456	338
rect	455	338	456	339
rect	455	339	456	340
rect	455	340	456	341
rect	455	341	456	342
rect	455	342	456	343
rect	455	343	456	344
rect	455	344	456	345
rect	455	345	456	346
rect	455	346	456	347
rect	455	347	456	348
rect	456	0	457	1
rect	456	1	457	2
rect	456	2	457	3
rect	456	3	457	4
rect	456	4	457	5
rect	456	5	457	6
rect	456	6	457	7
rect	456	7	457	8
rect	456	8	457	9
rect	456	9	457	10
rect	456	10	457	11
rect	456	11	457	12
rect	456	12	457	13
rect	456	13	457	14
rect	456	14	457	15
rect	456	15	457	16
rect	456	16	457	17
rect	456	17	457	18
rect	456	18	457	19
rect	456	19	457	20
rect	456	20	457	21
rect	456	21	457	22
rect	456	22	457	23
rect	456	23	457	24
rect	456	24	457	25
rect	456	25	457	26
rect	456	26	457	27
rect	456	27	457	28
rect	456	28	457	29
rect	456	29	457	30
rect	456	30	457	31
rect	456	31	457	32
rect	456	32	457	33
rect	456	33	457	34
rect	456	34	457	35
rect	456	35	457	36
rect	456	36	457	37
rect	456	37	457	38
rect	456	38	457	39
rect	456	39	457	40
rect	456	40	457	41
rect	456	41	457	42
rect	456	42	457	43
rect	456	43	457	44
rect	456	44	457	45
rect	456	45	457	46
rect	456	46	457	47
rect	456	47	457	48
rect	456	48	457	49
rect	456	49	457	50
rect	456	50	457	51
rect	456	51	457	52
rect	456	52	457	53
rect	456	53	457	54
rect	456	54	457	55
rect	456	55	457	56
rect	456	56	457	57
rect	456	57	457	58
rect	456	58	457	59
rect	456	59	457	60
rect	456	60	457	61
rect	456	61	457	62
rect	456	62	457	63
rect	456	63	457	64
rect	456	64	457	65
rect	456	65	457	66
rect	456	66	457	67
rect	456	67	457	68
rect	456	68	457	69
rect	456	69	457	70
rect	456	70	457	71
rect	456	71	457	72
rect	456	72	457	73
rect	456	73	457	74
rect	456	74	457	75
rect	456	75	457	76
rect	456	76	457	77
rect	456	77	457	78
rect	456	78	457	79
rect	456	79	457	80
rect	456	80	457	81
rect	456	81	457	82
rect	456	82	457	83
rect	456	83	457	84
rect	456	84	457	85
rect	456	85	457	86
rect	456	86	457	87
rect	456	87	457	88
rect	456	88	457	89
rect	456	89	457	90
rect	456	90	457	91
rect	456	91	457	92
rect	456	92	457	93
rect	456	93	457	94
rect	456	94	457	95
rect	456	95	457	96
rect	456	96	457	97
rect	456	97	457	98
rect	456	98	457	99
rect	456	99	457	100
rect	456	100	457	101
rect	456	101	457	102
rect	456	102	457	103
rect	456	103	457	104
rect	456	104	457	105
rect	456	105	457	106
rect	456	106	457	107
rect	456	107	457	108
rect	456	108	457	109
rect	456	109	457	110
rect	456	110	457	111
rect	456	111	457	112
rect	456	112	457	113
rect	456	113	457	114
rect	456	114	457	115
rect	456	115	457	116
rect	456	116	457	117
rect	456	117	457	118
rect	456	118	457	119
rect	456	119	457	120
rect	456	120	457	121
rect	456	121	457	122
rect	456	122	457	123
rect	456	123	457	124
rect	456	124	457	125
rect	456	125	457	126
rect	456	126	457	127
rect	456	127	457	128
rect	456	128	457	129
rect	456	129	457	130
rect	456	130	457	131
rect	456	131	457	132
rect	456	132	457	133
rect	456	133	457	134
rect	456	134	457	135
rect	456	135	457	136
rect	456	136	457	137
rect	456	137	457	138
rect	456	138	457	139
rect	456	139	457	140
rect	456	140	457	141
rect	456	141	457	142
rect	456	142	457	143
rect	456	143	457	144
rect	456	144	457	145
rect	456	145	457	146
rect	456	146	457	147
rect	456	147	457	148
rect	456	148	457	149
rect	456	149	457	150
rect	456	150	457	151
rect	456	151	457	152
rect	456	152	457	153
rect	456	153	457	154
rect	456	154	457	155
rect	456	155	457	156
rect	456	156	457	157
rect	456	157	457	158
rect	456	158	457	159
rect	456	159	457	160
rect	456	160	457	161
rect	456	161	457	162
rect	456	162	457	163
rect	456	163	457	164
rect	456	164	457	165
rect	456	165	457	166
rect	456	166	457	167
rect	456	167	457	168
rect	456	168	457	169
rect	456	169	457	170
rect	456	170	457	171
rect	456	171	457	172
rect	456	172	457	173
rect	456	173	457	174
rect	456	174	457	175
rect	456	175	457	176
rect	456	176	457	177
rect	456	177	457	178
rect	456	178	457	179
rect	456	179	457	180
rect	456	180	457	181
rect	456	181	457	182
rect	456	182	457	183
rect	456	183	457	184
rect	456	184	457	185
rect	456	185	457	186
rect	456	186	457	187
rect	456	187	457	188
rect	456	188	457	189
rect	456	189	457	190
rect	456	190	457	191
rect	456	191	457	192
rect	456	192	457	193
rect	456	193	457	194
rect	456	194	457	195
rect	456	195	457	196
rect	456	196	457	197
rect	456	197	457	198
rect	456	198	457	199
rect	456	199	457	200
rect	456	200	457	201
rect	456	201	457	202
rect	456	202	457	203
rect	456	203	457	204
rect	456	204	457	205
rect	456	205	457	206
rect	456	206	457	207
rect	456	207	457	208
rect	456	208	457	209
rect	456	209	457	210
rect	456	210	457	211
rect	456	211	457	212
rect	456	212	457	213
rect	456	213	457	214
rect	456	214	457	215
rect	456	215	457	216
rect	456	216	457	217
rect	456	217	457	218
rect	456	218	457	219
rect	456	219	457	220
rect	456	220	457	221
rect	456	221	457	222
rect	456	222	457	223
rect	456	223	457	224
rect	456	224	457	225
rect	456	225	457	226
rect	456	226	457	227
rect	456	227	457	228
rect	456	228	457	229
rect	456	229	457	230
rect	456	230	457	231
rect	456	231	457	232
rect	456	232	457	233
rect	456	233	457	234
rect	456	234	457	235
rect	456	235	457	236
rect	456	236	457	237
rect	456	237	457	238
rect	456	238	457	239
rect	456	239	457	240
rect	456	240	457	241
rect	456	241	457	242
rect	456	242	457	243
rect	456	243	457	244
rect	456	244	457	245
rect	456	245	457	246
rect	456	246	457	247
rect	456	247	457	248
rect	456	248	457	249
rect	456	249	457	250
rect	456	250	457	251
rect	456	251	457	252
rect	456	252	457	253
rect	456	253	457	254
rect	456	254	457	255
rect	456	255	457	256
rect	456	256	457	257
rect	456	257	457	258
rect	456	258	457	259
rect	456	259	457	260
rect	456	260	457	261
rect	456	261	457	262
rect	456	262	457	263
rect	456	263	457	264
rect	456	264	457	265
rect	456	265	457	266
rect	456	266	457	267
rect	456	267	457	268
rect	456	268	457	269
rect	456	269	457	270
rect	456	270	457	271
rect	456	271	457	272
rect	456	272	457	273
rect	456	273	457	274
rect	456	274	457	275
rect	456	275	457	276
rect	456	276	457	277
rect	456	277	457	278
rect	456	278	457	279
rect	456	279	457	280
rect	456	280	457	281
rect	456	281	457	282
rect	456	282	457	283
rect	456	283	457	284
rect	456	284	457	285
rect	456	285	457	286
rect	456	286	457	287
rect	456	287	457	288
rect	456	288	457	289
rect	456	289	457	290
rect	456	290	457	291
rect	456	291	457	292
rect	456	292	457	293
rect	456	293	457	294
rect	456	294	457	295
rect	456	295	457	296
rect	456	296	457	297
rect	456	297	457	298
rect	456	298	457	299
rect	456	299	457	300
rect	456	300	457	301
rect	456	301	457	302
rect	456	302	457	303
rect	456	303	457	304
rect	456	304	457	305
rect	456	305	457	306
rect	456	306	457	307
rect	456	307	457	308
rect	456	308	457	309
rect	456	309	457	310
rect	456	310	457	311
rect	456	311	457	312
rect	456	312	457	313
rect	456	313	457	314
rect	456	314	457	315
rect	456	315	457	316
rect	456	316	457	317
rect	456	317	457	318
rect	456	318	457	319
rect	456	319	457	320
rect	456	320	457	321
rect	456	321	457	322
rect	456	322	457	323
rect	456	323	457	324
rect	456	324	457	325
rect	456	325	457	326
rect	456	326	457	327
rect	456	327	457	328
rect	456	328	457	329
rect	456	329	457	330
rect	456	330	457	331
rect	456	331	457	332
rect	456	332	457	333
rect	456	333	457	334
rect	456	334	457	335
rect	456	335	457	336
rect	456	336	457	337
rect	456	337	457	338
rect	456	338	457	339
rect	456	339	457	340
rect	456	340	457	341
rect	456	341	457	342
rect	456	342	457	343
rect	456	343	457	344
rect	456	344	457	345
rect	456	345	457	346
rect	456	346	457	347
rect	456	347	457	348
rect	457	0	458	1
rect	457	1	458	2
rect	457	2	458	3
rect	457	3	458	4
rect	457	4	458	5
rect	457	5	458	6
rect	457	6	458	7
rect	457	7	458	8
rect	457	8	458	9
rect	457	9	458	10
rect	457	10	458	11
rect	457	11	458	12
rect	457	12	458	13
rect	457	13	458	14
rect	457	14	458	15
rect	457	15	458	16
rect	457	16	458	17
rect	457	17	458	18
rect	457	18	458	19
rect	457	19	458	20
rect	457	20	458	21
rect	457	21	458	22
rect	457	22	458	23
rect	457	23	458	24
rect	457	24	458	25
rect	457	25	458	26
rect	457	26	458	27
rect	457	27	458	28
rect	457	28	458	29
rect	457	29	458	30
rect	457	30	458	31
rect	457	31	458	32
rect	457	32	458	33
rect	457	33	458	34
rect	457	34	458	35
rect	457	35	458	36
rect	457	36	458	37
rect	457	37	458	38
rect	457	38	458	39
rect	457	39	458	40
rect	457	40	458	41
rect	457	41	458	42
rect	457	42	458	43
rect	457	43	458	44
rect	457	44	458	45
rect	457	45	458	46
rect	457	46	458	47
rect	457	47	458	48
rect	457	48	458	49
rect	457	49	458	50
rect	457	50	458	51
rect	457	51	458	52
rect	457	52	458	53
rect	457	53	458	54
rect	457	54	458	55
rect	457	55	458	56
rect	457	56	458	57
rect	457	57	458	58
rect	457	58	458	59
rect	457	59	458	60
rect	457	60	458	61
rect	457	61	458	62
rect	457	62	458	63
rect	457	63	458	64
rect	457	64	458	65
rect	457	65	458	66
rect	457	66	458	67
rect	457	67	458	68
rect	457	68	458	69
rect	457	69	458	70
rect	457	70	458	71
rect	457	71	458	72
rect	457	72	458	73
rect	457	73	458	74
rect	457	74	458	75
rect	457	75	458	76
rect	457	76	458	77
rect	457	77	458	78
rect	457	78	458	79
rect	457	79	458	80
rect	457	80	458	81
rect	457	81	458	82
rect	457	82	458	83
rect	457	83	458	84
rect	457	84	458	85
rect	457	85	458	86
rect	457	86	458	87
rect	457	87	458	88
rect	457	88	458	89
rect	457	89	458	90
rect	457	90	458	91
rect	457	91	458	92
rect	457	92	458	93
rect	457	93	458	94
rect	457	94	458	95
rect	457	95	458	96
rect	457	96	458	97
rect	457	97	458	98
rect	457	98	458	99
rect	457	99	458	100
rect	457	100	458	101
rect	457	101	458	102
rect	457	102	458	103
rect	457	103	458	104
rect	457	104	458	105
rect	457	105	458	106
rect	457	106	458	107
rect	457	107	458	108
rect	457	108	458	109
rect	457	109	458	110
rect	457	110	458	111
rect	457	111	458	112
rect	457	112	458	113
rect	457	113	458	114
rect	457	114	458	115
rect	457	115	458	116
rect	457	116	458	117
rect	457	117	458	118
rect	457	118	458	119
rect	457	119	458	120
rect	457	120	458	121
rect	457	121	458	122
rect	457	122	458	123
rect	457	123	458	124
rect	457	124	458	125
rect	457	125	458	126
rect	457	126	458	127
rect	457	127	458	128
rect	457	128	458	129
rect	457	129	458	130
rect	457	130	458	131
rect	457	131	458	132
rect	457	132	458	133
rect	457	133	458	134
rect	457	134	458	135
rect	457	135	458	136
rect	457	136	458	137
rect	457	137	458	138
rect	457	138	458	139
rect	457	139	458	140
rect	457	140	458	141
rect	457	141	458	142
rect	457	142	458	143
rect	457	143	458	144
rect	457	144	458	145
rect	457	145	458	146
rect	457	146	458	147
rect	457	147	458	148
rect	457	148	458	149
rect	457	149	458	150
rect	457	150	458	151
rect	457	151	458	152
rect	457	152	458	153
rect	457	153	458	154
rect	457	154	458	155
rect	457	155	458	156
rect	457	156	458	157
rect	457	157	458	158
rect	457	158	458	159
rect	457	159	458	160
rect	457	160	458	161
rect	457	161	458	162
rect	457	162	458	163
rect	457	163	458	164
rect	457	164	458	165
rect	457	165	458	166
rect	457	166	458	167
rect	457	167	458	168
rect	457	168	458	169
rect	457	169	458	170
rect	457	170	458	171
rect	457	171	458	172
rect	457	172	458	173
rect	457	173	458	174
rect	457	174	458	175
rect	457	175	458	176
rect	457	176	458	177
rect	457	177	458	178
rect	457	178	458	179
rect	457	179	458	180
rect	457	180	458	181
rect	457	181	458	182
rect	457	182	458	183
rect	457	183	458	184
rect	457	184	458	185
rect	457	185	458	186
rect	457	186	458	187
rect	457	187	458	188
rect	457	188	458	189
rect	457	189	458	190
rect	457	190	458	191
rect	457	191	458	192
rect	457	192	458	193
rect	457	193	458	194
rect	457	194	458	195
rect	457	195	458	196
rect	457	196	458	197
rect	457	197	458	198
rect	457	198	458	199
rect	457	199	458	200
rect	457	200	458	201
rect	457	201	458	202
rect	457	202	458	203
rect	457	203	458	204
rect	457	204	458	205
rect	457	205	458	206
rect	457	206	458	207
rect	457	207	458	208
rect	457	208	458	209
rect	457	209	458	210
rect	457	210	458	211
rect	457	211	458	212
rect	457	212	458	213
rect	457	213	458	214
rect	457	214	458	215
rect	457	215	458	216
rect	457	216	458	217
rect	457	217	458	218
rect	457	218	458	219
rect	457	219	458	220
rect	457	220	458	221
rect	457	221	458	222
rect	457	222	458	223
rect	457	223	458	224
rect	457	224	458	225
rect	457	225	458	226
rect	457	226	458	227
rect	457	227	458	228
rect	457	228	458	229
rect	457	229	458	230
rect	457	230	458	231
rect	457	231	458	232
rect	457	232	458	233
rect	457	233	458	234
rect	457	234	458	235
rect	457	235	458	236
rect	457	236	458	237
rect	457	237	458	238
rect	457	238	458	239
rect	457	239	458	240
rect	457	240	458	241
rect	457	241	458	242
rect	457	242	458	243
rect	457	243	458	244
rect	457	244	458	245
rect	457	245	458	246
rect	457	246	458	247
rect	457	247	458	248
rect	457	248	458	249
rect	457	249	458	250
rect	457	250	458	251
rect	457	251	458	252
rect	457	252	458	253
rect	457	253	458	254
rect	457	254	458	255
rect	457	255	458	256
rect	457	256	458	257
rect	457	257	458	258
rect	457	258	458	259
rect	457	259	458	260
rect	457	260	458	261
rect	457	261	458	262
rect	457	262	458	263
rect	457	263	458	264
rect	457	264	458	265
rect	457	265	458	266
rect	457	266	458	267
rect	457	267	458	268
rect	457	268	458	269
rect	457	269	458	270
rect	457	270	458	271
rect	457	271	458	272
rect	457	272	458	273
rect	457	273	458	274
rect	457	274	458	275
rect	457	275	458	276
rect	457	276	458	277
rect	457	277	458	278
rect	457	278	458	279
rect	457	279	458	280
rect	457	280	458	281
rect	457	281	458	282
rect	457	282	458	283
rect	457	283	458	284
rect	457	284	458	285
rect	457	285	458	286
rect	457	286	458	287
rect	457	287	458	288
rect	457	288	458	289
rect	457	289	458	290
rect	457	290	458	291
rect	457	291	458	292
rect	457	292	458	293
rect	457	293	458	294
rect	457	294	458	295
rect	457	295	458	296
rect	457	296	458	297
rect	457	297	458	298
rect	457	298	458	299
rect	457	299	458	300
rect	457	300	458	301
rect	457	301	458	302
rect	457	302	458	303
rect	457	303	458	304
rect	457	304	458	305
rect	457	305	458	306
rect	457	306	458	307
rect	457	307	458	308
rect	457	308	458	309
rect	457	309	458	310
rect	457	310	458	311
rect	457	311	458	312
rect	457	312	458	313
rect	457	313	458	314
rect	457	314	458	315
rect	457	315	458	316
rect	457	316	458	317
rect	457	317	458	318
rect	457	318	458	319
rect	457	319	458	320
rect	457	320	458	321
rect	457	321	458	322
rect	457	322	458	323
rect	457	323	458	324
rect	457	324	458	325
rect	457	325	458	326
rect	457	326	458	327
rect	457	327	458	328
rect	457	328	458	329
rect	457	329	458	330
rect	457	330	458	331
rect	457	331	458	332
rect	457	332	458	333
rect	457	333	458	334
rect	457	334	458	335
rect	457	335	458	336
rect	457	336	458	337
rect	457	337	458	338
rect	457	338	458	339
rect	457	339	458	340
rect	457	340	458	341
rect	457	341	458	342
rect	457	342	458	343
rect	457	343	458	344
rect	457	344	458	345
rect	457	345	458	346
rect	457	346	458	347
rect	457	347	458	348
rect	475	257	476	258
rect	475	258	476	259
rect	475	260	476	261
rect	475	261	476	262
rect	475	262	476	263
rect	475	263	476	264
rect	475	264	476	265
rect	489	0	490	1
rect	489	1	490	2
rect	489	2	490	3
rect	489	3	490	4
rect	489	4	490	5
rect	489	5	490	6
rect	489	6	490	7
rect	489	7	490	8
rect	489	8	490	9
rect	489	9	490	10
rect	489	10	490	11
rect	489	11	490	12
rect	489	12	490	13
rect	489	13	490	14
rect	489	14	490	15
rect	489	15	490	16
rect	489	16	490	17
rect	489	17	490	18
rect	489	18	490	19
rect	489	19	490	20
rect	489	20	490	21
rect	489	21	490	22
rect	489	22	490	23
rect	489	23	490	24
rect	489	24	490	25
rect	489	25	490	26
rect	489	26	490	27
rect	489	27	490	28
rect	489	28	490	29
rect	489	29	490	30
rect	489	30	490	31
rect	489	31	490	32
rect	489	32	490	33
rect	489	33	490	34
rect	489	34	490	35
rect	489	35	490	36
rect	489	36	490	37
rect	489	37	490	38
rect	489	38	490	39
rect	489	39	490	40
rect	489	40	490	41
rect	489	41	490	42
rect	489	42	490	43
rect	489	43	490	44
rect	489	44	490	45
rect	489	45	490	46
rect	489	46	490	47
rect	489	47	490	48
rect	489	48	490	49
rect	489	49	490	50
rect	489	50	490	51
rect	489	51	490	52
rect	489	52	490	53
rect	489	53	490	54
rect	489	54	490	55
rect	489	55	490	56
rect	489	56	490	57
rect	489	57	490	58
rect	489	58	490	59
rect	489	59	490	60
rect	489	60	490	61
rect	489	61	490	62
rect	489	62	490	63
rect	489	63	490	64
rect	489	64	490	65
rect	489	65	490	66
rect	489	66	490	67
rect	489	67	490	68
rect	489	68	490	69
rect	489	69	490	70
rect	489	70	490	71
rect	489	71	490	72
rect	489	72	490	73
rect	489	73	490	74
rect	489	74	490	75
rect	489	75	490	76
rect	489	76	490	77
rect	489	77	490	78
rect	489	78	490	79
rect	489	79	490	80
rect	489	80	490	81
rect	489	81	490	82
rect	489	82	490	83
rect	489	83	490	84
rect	489	84	490	85
rect	489	85	490	86
rect	489	86	490	87
rect	489	87	490	88
rect	489	88	490	89
rect	489	89	490	90
rect	489	90	490	91
rect	489	91	490	92
rect	489	92	490	93
rect	489	93	490	94
rect	489	94	490	95
rect	489	95	490	96
rect	489	96	490	97
rect	489	97	490	98
rect	489	98	490	99
rect	489	99	490	100
rect	489	100	490	101
rect	489	101	490	102
rect	489	102	490	103
rect	489	103	490	104
rect	489	104	490	105
rect	489	105	490	106
rect	489	106	490	107
rect	489	107	490	108
rect	489	108	490	109
rect	489	109	490	110
rect	489	110	490	111
rect	489	111	490	112
rect	489	112	490	113
rect	489	113	490	114
rect	489	114	490	115
rect	489	115	490	116
rect	489	116	490	117
rect	489	117	490	118
rect	489	118	490	119
rect	489	119	490	120
rect	489	120	490	121
rect	489	121	490	122
rect	489	122	490	123
rect	489	123	490	124
rect	489	124	490	125
rect	489	125	490	126
rect	489	126	490	127
rect	489	127	490	128
rect	489	128	490	129
rect	489	129	490	130
rect	489	130	490	131
rect	489	131	490	132
rect	489	132	490	133
rect	489	133	490	134
rect	489	134	490	135
rect	489	135	490	136
rect	489	136	490	137
rect	489	137	490	138
rect	489	138	490	139
rect	489	139	490	140
rect	489	140	490	141
rect	489	141	490	142
rect	489	142	490	143
rect	489	143	490	144
rect	489	144	490	145
rect	489	145	490	146
rect	489	146	490	147
rect	489	147	490	148
rect	489	148	490	149
rect	489	149	490	150
rect	489	150	490	151
rect	489	151	490	152
rect	489	152	490	153
rect	489	153	490	154
rect	489	154	490	155
rect	489	155	490	156
rect	489	156	490	157
rect	489	157	490	158
rect	489	158	490	159
rect	489	159	490	160
rect	489	160	490	161
rect	489	161	490	162
rect	489	162	490	163
rect	489	163	490	164
rect	489	164	490	165
rect	489	165	490	166
rect	489	166	490	167
rect	489	167	490	168
rect	489	168	490	169
rect	489	169	490	170
rect	489	170	490	171
rect	489	171	490	172
rect	489	172	490	173
rect	489	173	490	174
rect	489	174	490	175
rect	489	175	490	176
rect	489	176	490	177
rect	489	177	490	178
rect	489	178	490	179
rect	489	179	490	180
rect	489	180	490	181
rect	489	181	490	182
rect	489	182	490	183
rect	489	183	490	184
rect	489	184	490	185
rect	489	185	490	186
rect	489	186	490	187
rect	489	187	490	188
rect	489	188	490	189
rect	489	189	490	190
rect	489	190	490	191
rect	489	191	490	192
rect	489	192	490	193
rect	489	193	490	194
rect	489	194	490	195
rect	489	195	490	196
rect	489	196	490	197
rect	489	197	490	198
rect	489	198	490	199
rect	489	199	490	200
rect	489	200	490	201
rect	489	201	490	202
rect	489	202	490	203
rect	489	203	490	204
rect	489	204	490	205
rect	489	205	490	206
rect	489	206	490	207
rect	489	207	490	208
rect	489	208	490	209
rect	489	209	490	210
rect	489	210	490	211
rect	489	211	490	212
rect	489	212	490	213
rect	489	213	490	214
rect	489	214	490	215
rect	489	215	490	216
rect	489	216	490	217
rect	489	217	490	218
rect	489	218	490	219
rect	489	219	490	220
rect	489	220	490	221
rect	489	221	490	222
rect	489	222	490	223
rect	489	223	490	224
rect	489	224	490	225
rect	489	225	490	226
rect	489	226	490	227
rect	489	227	490	228
rect	489	228	490	229
rect	489	229	490	230
rect	489	230	490	231
rect	489	231	490	232
rect	489	232	490	233
rect	489	233	490	234
rect	489	234	490	235
rect	489	235	490	236
rect	489	236	490	237
rect	489	237	490	238
rect	489	238	490	239
rect	489	239	490	240
rect	489	240	490	241
rect	489	241	490	242
rect	489	242	490	243
rect	489	243	490	244
rect	489	244	490	245
rect	489	245	490	246
rect	489	246	490	247
rect	489	247	490	248
rect	489	248	490	249
rect	489	249	490	250
rect	489	250	490	251
rect	489	251	490	252
rect	489	252	490	253
rect	489	253	490	254
rect	489	254	490	255
rect	489	255	490	256
rect	489	256	490	257
rect	489	257	490	258
rect	489	258	490	259
rect	489	259	490	260
rect	489	260	490	261
rect	489	261	490	262
rect	489	262	490	263
rect	489	263	490	264
rect	489	264	490	265
rect	489	265	490	266
rect	489	266	490	267
rect	489	267	490	268
rect	489	268	490	269
rect	489	269	490	270
rect	489	270	490	271
rect	489	271	490	272
rect	489	272	490	273
rect	489	273	490	274
rect	489	274	490	275
rect	489	275	490	276
rect	489	276	490	277
rect	489	277	490	278
rect	489	278	490	279
rect	489	279	490	280
rect	489	280	490	281
rect	489	281	490	282
rect	489	282	490	283
rect	489	283	490	284
rect	489	284	490	285
rect	489	285	490	286
rect	489	286	490	287
rect	489	287	490	288
rect	489	288	490	289
rect	489	289	490	290
rect	489	290	490	291
rect	489	291	490	292
rect	489	292	490	293
rect	489	293	490	294
rect	489	294	490	295
rect	489	295	490	296
rect	489	296	490	297
rect	489	297	490	298
rect	489	298	490	299
rect	489	299	490	300
rect	489	300	490	301
rect	489	301	490	302
rect	489	302	490	303
rect	489	303	490	304
rect	489	304	490	305
rect	489	305	490	306
rect	489	306	490	307
rect	489	307	490	308
rect	489	308	490	309
rect	489	309	490	310
rect	489	310	490	311
rect	489	311	490	312
rect	489	312	490	313
rect	489	313	490	314
rect	489	314	490	315
rect	489	315	490	316
rect	489	316	490	317
rect	489	317	490	318
rect	489	318	490	319
rect	489	319	490	320
rect	489	320	490	321
rect	490	0	491	1
rect	490	1	491	2
rect	490	2	491	3
rect	490	3	491	4
rect	490	4	491	5
rect	490	5	491	6
rect	490	6	491	7
rect	490	7	491	8
rect	490	8	491	9
rect	490	9	491	10
rect	490	10	491	11
rect	490	11	491	12
rect	490	12	491	13
rect	490	13	491	14
rect	490	14	491	15
rect	490	15	491	16
rect	490	16	491	17
rect	490	17	491	18
rect	490	18	491	19
rect	490	19	491	20
rect	490	20	491	21
rect	490	21	491	22
rect	490	22	491	23
rect	490	23	491	24
rect	490	24	491	25
rect	490	25	491	26
rect	490	26	491	27
rect	490	27	491	28
rect	490	28	491	29
rect	490	29	491	30
rect	490	30	491	31
rect	490	31	491	32
rect	490	32	491	33
rect	490	33	491	34
rect	490	34	491	35
rect	490	35	491	36
rect	490	36	491	37
rect	490	37	491	38
rect	490	38	491	39
rect	490	39	491	40
rect	490	40	491	41
rect	490	41	491	42
rect	490	42	491	43
rect	490	43	491	44
rect	490	44	491	45
rect	490	45	491	46
rect	490	46	491	47
rect	490	47	491	48
rect	490	48	491	49
rect	490	49	491	50
rect	490	50	491	51
rect	490	51	491	52
rect	490	52	491	53
rect	490	53	491	54
rect	490	54	491	55
rect	490	55	491	56
rect	490	56	491	57
rect	490	57	491	58
rect	490	58	491	59
rect	490	59	491	60
rect	490	60	491	61
rect	490	61	491	62
rect	490	62	491	63
rect	490	63	491	64
rect	490	64	491	65
rect	490	65	491	66
rect	490	66	491	67
rect	490	67	491	68
rect	490	68	491	69
rect	490	69	491	70
rect	490	70	491	71
rect	490	71	491	72
rect	490	72	491	73
rect	490	73	491	74
rect	490	74	491	75
rect	490	75	491	76
rect	490	76	491	77
rect	490	77	491	78
rect	490	78	491	79
rect	490	79	491	80
rect	490	80	491	81
rect	490	81	491	82
rect	490	82	491	83
rect	490	83	491	84
rect	490	84	491	85
rect	490	85	491	86
rect	490	86	491	87
rect	490	87	491	88
rect	490	88	491	89
rect	490	89	491	90
rect	490	90	491	91
rect	490	91	491	92
rect	490	92	491	93
rect	490	93	491	94
rect	490	94	491	95
rect	490	95	491	96
rect	490	96	491	97
rect	490	97	491	98
rect	490	98	491	99
rect	490	99	491	100
rect	490	100	491	101
rect	490	101	491	102
rect	490	102	491	103
rect	490	103	491	104
rect	490	104	491	105
rect	490	105	491	106
rect	490	106	491	107
rect	490	107	491	108
rect	490	108	491	109
rect	490	109	491	110
rect	490	110	491	111
rect	490	111	491	112
rect	490	112	491	113
rect	490	113	491	114
rect	490	114	491	115
rect	490	115	491	116
rect	490	116	491	117
rect	490	117	491	118
rect	490	118	491	119
rect	490	119	491	120
rect	490	120	491	121
rect	490	121	491	122
rect	490	122	491	123
rect	490	123	491	124
rect	490	124	491	125
rect	490	125	491	126
rect	490	126	491	127
rect	490	127	491	128
rect	490	128	491	129
rect	490	129	491	130
rect	490	130	491	131
rect	490	131	491	132
rect	490	132	491	133
rect	490	133	491	134
rect	490	134	491	135
rect	490	135	491	136
rect	490	136	491	137
rect	490	137	491	138
rect	490	138	491	139
rect	490	139	491	140
rect	490	140	491	141
rect	490	141	491	142
rect	490	142	491	143
rect	490	143	491	144
rect	490	144	491	145
rect	490	145	491	146
rect	490	146	491	147
rect	490	147	491	148
rect	490	148	491	149
rect	490	149	491	150
rect	490	150	491	151
rect	490	151	491	152
rect	490	152	491	153
rect	490	153	491	154
rect	490	154	491	155
rect	490	155	491	156
rect	490	156	491	157
rect	490	157	491	158
rect	490	158	491	159
rect	490	159	491	160
rect	490	160	491	161
rect	490	161	491	162
rect	490	162	491	163
rect	490	163	491	164
rect	490	164	491	165
rect	490	165	491	166
rect	490	166	491	167
rect	490	167	491	168
rect	490	168	491	169
rect	490	169	491	170
rect	490	170	491	171
rect	490	171	491	172
rect	490	172	491	173
rect	490	173	491	174
rect	490	174	491	175
rect	490	175	491	176
rect	490	176	491	177
rect	490	177	491	178
rect	490	178	491	179
rect	490	179	491	180
rect	490	180	491	181
rect	490	181	491	182
rect	490	182	491	183
rect	490	183	491	184
rect	490	184	491	185
rect	490	185	491	186
rect	490	186	491	187
rect	490	187	491	188
rect	490	188	491	189
rect	490	189	491	190
rect	490	190	491	191
rect	490	191	491	192
rect	490	192	491	193
rect	490	193	491	194
rect	490	194	491	195
rect	490	195	491	196
rect	490	196	491	197
rect	490	197	491	198
rect	490	198	491	199
rect	490	199	491	200
rect	490	200	491	201
rect	490	201	491	202
rect	490	202	491	203
rect	490	203	491	204
rect	490	204	491	205
rect	490	205	491	206
rect	490	206	491	207
rect	490	207	491	208
rect	490	208	491	209
rect	490	209	491	210
rect	490	210	491	211
rect	490	211	491	212
rect	490	212	491	213
rect	490	213	491	214
rect	490	214	491	215
rect	490	215	491	216
rect	490	216	491	217
rect	490	217	491	218
rect	490	218	491	219
rect	490	219	491	220
rect	490	220	491	221
rect	490	221	491	222
rect	490	222	491	223
rect	490	223	491	224
rect	490	224	491	225
rect	490	225	491	226
rect	490	226	491	227
rect	490	227	491	228
rect	490	228	491	229
rect	490	229	491	230
rect	490	230	491	231
rect	490	231	491	232
rect	490	232	491	233
rect	490	233	491	234
rect	490	234	491	235
rect	490	235	491	236
rect	490	236	491	237
rect	490	237	491	238
rect	490	238	491	239
rect	490	239	491	240
rect	490	240	491	241
rect	490	241	491	242
rect	490	242	491	243
rect	490	243	491	244
rect	490	244	491	245
rect	490	245	491	246
rect	490	246	491	247
rect	490	247	491	248
rect	490	248	491	249
rect	490	249	491	250
rect	490	250	491	251
rect	490	251	491	252
rect	490	252	491	253
rect	490	253	491	254
rect	490	254	491	255
rect	490	255	491	256
rect	490	256	491	257
rect	490	257	491	258
rect	490	258	491	259
rect	490	259	491	260
rect	490	260	491	261
rect	490	261	491	262
rect	490	262	491	263
rect	490	263	491	264
rect	490	264	491	265
rect	490	265	491	266
rect	490	266	491	267
rect	490	267	491	268
rect	490	268	491	269
rect	490	269	491	270
rect	490	270	491	271
rect	490	271	491	272
rect	490	272	491	273
rect	490	273	491	274
rect	490	274	491	275
rect	490	275	491	276
rect	490	276	491	277
rect	490	277	491	278
rect	490	278	491	279
rect	490	279	491	280
rect	490	280	491	281
rect	490	281	491	282
rect	490	282	491	283
rect	490	283	491	284
rect	490	284	491	285
rect	490	285	491	286
rect	490	286	491	287
rect	490	287	491	288
rect	490	288	491	289
rect	490	289	491	290
rect	490	290	491	291
rect	490	291	491	292
rect	490	292	491	293
rect	490	293	491	294
rect	490	294	491	295
rect	490	295	491	296
rect	490	296	491	297
rect	490	297	491	298
rect	490	298	491	299
rect	490	299	491	300
rect	490	300	491	301
rect	490	301	491	302
rect	490	302	491	303
rect	490	303	491	304
rect	490	304	491	305
rect	490	305	491	306
rect	490	306	491	307
rect	490	307	491	308
rect	490	308	491	309
rect	490	309	491	310
rect	490	310	491	311
rect	490	311	491	312
rect	490	312	491	313
rect	490	313	491	314
rect	490	314	491	315
rect	490	315	491	316
rect	490	316	491	317
rect	490	317	491	318
rect	490	318	491	319
rect	490	319	491	320
rect	490	320	491	321
rect	491	0	492	1
rect	491	1	492	2
rect	491	2	492	3
rect	491	3	492	4
rect	491	4	492	5
rect	491	5	492	6
rect	491	6	492	7
rect	491	7	492	8
rect	491	8	492	9
rect	491	9	492	10
rect	491	10	492	11
rect	491	11	492	12
rect	491	12	492	13
rect	491	13	492	14
rect	491	14	492	15
rect	491	15	492	16
rect	491	16	492	17
rect	491	17	492	18
rect	491	18	492	19
rect	491	19	492	20
rect	491	20	492	21
rect	491	21	492	22
rect	491	22	492	23
rect	491	23	492	24
rect	491	24	492	25
rect	491	25	492	26
rect	491	26	492	27
rect	491	27	492	28
rect	491	28	492	29
rect	491	29	492	30
rect	491	30	492	31
rect	491	31	492	32
rect	491	32	492	33
rect	491	33	492	34
rect	491	34	492	35
rect	491	35	492	36
rect	491	36	492	37
rect	491	37	492	38
rect	491	38	492	39
rect	491	39	492	40
rect	491	40	492	41
rect	491	41	492	42
rect	491	42	492	43
rect	491	43	492	44
rect	491	44	492	45
rect	491	45	492	46
rect	491	46	492	47
rect	491	47	492	48
rect	491	48	492	49
rect	491	49	492	50
rect	491	50	492	51
rect	491	51	492	52
rect	491	52	492	53
rect	491	53	492	54
rect	491	54	492	55
rect	491	55	492	56
rect	491	56	492	57
rect	491	57	492	58
rect	491	58	492	59
rect	491	59	492	60
rect	491	60	492	61
rect	491	61	492	62
rect	491	62	492	63
rect	491	63	492	64
rect	491	64	492	65
rect	491	65	492	66
rect	491	66	492	67
rect	491	67	492	68
rect	491	68	492	69
rect	491	69	492	70
rect	491	70	492	71
rect	491	71	492	72
rect	491	72	492	73
rect	491	73	492	74
rect	491	74	492	75
rect	491	75	492	76
rect	491	76	492	77
rect	491	77	492	78
rect	491	78	492	79
rect	491	79	492	80
rect	491	80	492	81
rect	491	81	492	82
rect	491	82	492	83
rect	491	83	492	84
rect	491	84	492	85
rect	491	85	492	86
rect	491	86	492	87
rect	491	87	492	88
rect	491	88	492	89
rect	491	89	492	90
rect	491	90	492	91
rect	491	91	492	92
rect	491	92	492	93
rect	491	93	492	94
rect	491	94	492	95
rect	491	95	492	96
rect	491	96	492	97
rect	491	97	492	98
rect	491	98	492	99
rect	491	99	492	100
rect	491	100	492	101
rect	491	101	492	102
rect	491	102	492	103
rect	491	103	492	104
rect	491	104	492	105
rect	491	105	492	106
rect	491	106	492	107
rect	491	107	492	108
rect	491	108	492	109
rect	491	109	492	110
rect	491	110	492	111
rect	491	111	492	112
rect	491	112	492	113
rect	491	113	492	114
rect	491	114	492	115
rect	491	115	492	116
rect	491	116	492	117
rect	491	117	492	118
rect	491	118	492	119
rect	491	119	492	120
rect	491	120	492	121
rect	491	121	492	122
rect	491	122	492	123
rect	491	123	492	124
rect	491	124	492	125
rect	491	125	492	126
rect	491	126	492	127
rect	491	127	492	128
rect	491	128	492	129
rect	491	129	492	130
rect	491	130	492	131
rect	491	131	492	132
rect	491	132	492	133
rect	491	133	492	134
rect	491	134	492	135
rect	491	135	492	136
rect	491	136	492	137
rect	491	137	492	138
rect	491	138	492	139
rect	491	139	492	140
rect	491	140	492	141
rect	491	141	492	142
rect	491	142	492	143
rect	491	143	492	144
rect	491	144	492	145
rect	491	145	492	146
rect	491	146	492	147
rect	491	147	492	148
rect	491	148	492	149
rect	491	149	492	150
rect	491	150	492	151
rect	491	151	492	152
rect	491	152	492	153
rect	491	153	492	154
rect	491	154	492	155
rect	491	155	492	156
rect	491	156	492	157
rect	491	157	492	158
rect	491	158	492	159
rect	491	159	492	160
rect	491	160	492	161
rect	491	161	492	162
rect	491	162	492	163
rect	491	163	492	164
rect	491	164	492	165
rect	491	165	492	166
rect	491	166	492	167
rect	491	167	492	168
rect	491	168	492	169
rect	491	169	492	170
rect	491	170	492	171
rect	491	171	492	172
rect	491	172	492	173
rect	491	173	492	174
rect	491	174	492	175
rect	491	175	492	176
rect	491	176	492	177
rect	491	177	492	178
rect	491	178	492	179
rect	491	179	492	180
rect	491	180	492	181
rect	491	181	492	182
rect	491	182	492	183
rect	491	183	492	184
rect	491	184	492	185
rect	491	185	492	186
rect	491	186	492	187
rect	491	187	492	188
rect	491	188	492	189
rect	491	189	492	190
rect	491	190	492	191
rect	491	191	492	192
rect	491	192	492	193
rect	491	193	492	194
rect	491	194	492	195
rect	491	195	492	196
rect	491	196	492	197
rect	491	197	492	198
rect	491	198	492	199
rect	491	199	492	200
rect	491	200	492	201
rect	491	201	492	202
rect	491	202	492	203
rect	491	203	492	204
rect	491	204	492	205
rect	491	205	492	206
rect	491	206	492	207
rect	491	207	492	208
rect	491	208	492	209
rect	491	209	492	210
rect	491	210	492	211
rect	491	211	492	212
rect	491	212	492	213
rect	491	213	492	214
rect	491	214	492	215
rect	491	215	492	216
rect	491	216	492	217
rect	491	217	492	218
rect	491	218	492	219
rect	491	219	492	220
rect	491	220	492	221
rect	491	221	492	222
rect	491	222	492	223
rect	491	223	492	224
rect	491	224	492	225
rect	491	225	492	226
rect	491	226	492	227
rect	491	227	492	228
rect	491	228	492	229
rect	491	229	492	230
rect	491	230	492	231
rect	491	231	492	232
rect	491	232	492	233
rect	491	233	492	234
rect	491	234	492	235
rect	491	235	492	236
rect	491	236	492	237
rect	491	237	492	238
rect	491	238	492	239
rect	491	239	492	240
rect	491	240	492	241
rect	491	241	492	242
rect	491	242	492	243
rect	491	243	492	244
rect	491	244	492	245
rect	491	245	492	246
rect	491	246	492	247
rect	491	247	492	248
rect	491	248	492	249
rect	491	249	492	250
rect	491	250	492	251
rect	491	251	492	252
rect	491	252	492	253
rect	491	253	492	254
rect	491	254	492	255
rect	491	255	492	256
rect	491	256	492	257
rect	491	257	492	258
rect	491	258	492	259
rect	491	259	492	260
rect	491	260	492	261
rect	491	261	492	262
rect	491	262	492	263
rect	491	263	492	264
rect	491	264	492	265
rect	491	265	492	266
rect	491	266	492	267
rect	491	267	492	268
rect	491	268	492	269
rect	491	269	492	270
rect	491	270	492	271
rect	491	271	492	272
rect	491	272	492	273
rect	491	273	492	274
rect	491	274	492	275
rect	491	275	492	276
rect	491	276	492	277
rect	491	277	492	278
rect	491	278	492	279
rect	491	279	492	280
rect	491	280	492	281
rect	491	281	492	282
rect	491	282	492	283
rect	491	283	492	284
rect	491	284	492	285
rect	491	285	492	286
rect	491	286	492	287
rect	491	287	492	288
rect	491	288	492	289
rect	491	289	492	290
rect	491	290	492	291
rect	491	291	492	292
rect	491	292	492	293
rect	491	293	492	294
rect	491	294	492	295
rect	491	295	492	296
rect	491	296	492	297
rect	491	297	492	298
rect	491	298	492	299
rect	491	299	492	300
rect	491	300	492	301
rect	491	301	492	302
rect	491	302	492	303
rect	491	303	492	304
rect	491	304	492	305
rect	491	305	492	306
rect	491	306	492	307
rect	491	307	492	308
rect	491	308	492	309
rect	491	309	492	310
rect	491	310	492	311
rect	491	311	492	312
rect	491	312	492	313
rect	491	313	492	314
rect	491	314	492	315
rect	491	315	492	316
rect	491	316	492	317
rect	491	317	492	318
rect	491	318	492	319
rect	491	319	492	320
rect	491	320	492	321
rect	492	0	493	1
rect	492	1	493	2
rect	492	2	493	3
rect	492	3	493	4
rect	492	4	493	5
rect	492	5	493	6
rect	492	6	493	7
rect	492	7	493	8
rect	492	8	493	9
rect	492	9	493	10
rect	492	10	493	11
rect	492	11	493	12
rect	492	12	493	13
rect	492	13	493	14
rect	492	14	493	15
rect	492	15	493	16
rect	492	16	493	17
rect	492	17	493	18
rect	492	18	493	19
rect	492	19	493	20
rect	492	20	493	21
rect	492	21	493	22
rect	492	22	493	23
rect	492	23	493	24
rect	492	24	493	25
rect	492	25	493	26
rect	492	26	493	27
rect	492	27	493	28
rect	492	28	493	29
rect	492	29	493	30
rect	492	30	493	31
rect	492	31	493	32
rect	492	32	493	33
rect	492	33	493	34
rect	492	34	493	35
rect	492	35	493	36
rect	492	36	493	37
rect	492	37	493	38
rect	492	38	493	39
rect	492	39	493	40
rect	492	40	493	41
rect	492	41	493	42
rect	492	42	493	43
rect	492	43	493	44
rect	492	44	493	45
rect	492	45	493	46
rect	492	46	493	47
rect	492	47	493	48
rect	492	48	493	49
rect	492	49	493	50
rect	492	50	493	51
rect	492	51	493	52
rect	492	52	493	53
rect	492	53	493	54
rect	492	54	493	55
rect	492	55	493	56
rect	492	56	493	57
rect	492	57	493	58
rect	492	58	493	59
rect	492	59	493	60
rect	492	60	493	61
rect	492	61	493	62
rect	492	62	493	63
rect	492	63	493	64
rect	492	64	493	65
rect	492	65	493	66
rect	492	66	493	67
rect	492	67	493	68
rect	492	68	493	69
rect	492	69	493	70
rect	492	70	493	71
rect	492	71	493	72
rect	492	72	493	73
rect	492	73	493	74
rect	492	74	493	75
rect	492	75	493	76
rect	492	76	493	77
rect	492	77	493	78
rect	492	78	493	79
rect	492	79	493	80
rect	492	80	493	81
rect	492	81	493	82
rect	492	82	493	83
rect	492	83	493	84
rect	492	84	493	85
rect	492	85	493	86
rect	492	86	493	87
rect	492	87	493	88
rect	492	88	493	89
rect	492	89	493	90
rect	492	90	493	91
rect	492	91	493	92
rect	492	92	493	93
rect	492	93	493	94
rect	492	94	493	95
rect	492	95	493	96
rect	492	96	493	97
rect	492	97	493	98
rect	492	98	493	99
rect	492	99	493	100
rect	492	100	493	101
rect	492	101	493	102
rect	492	102	493	103
rect	492	103	493	104
rect	492	104	493	105
rect	492	105	493	106
rect	492	106	493	107
rect	492	107	493	108
rect	492	108	493	109
rect	492	109	493	110
rect	492	110	493	111
rect	492	111	493	112
rect	492	112	493	113
rect	492	113	493	114
rect	492	114	493	115
rect	492	115	493	116
rect	492	116	493	117
rect	492	117	493	118
rect	492	118	493	119
rect	492	119	493	120
rect	492	120	493	121
rect	492	121	493	122
rect	492	122	493	123
rect	492	123	493	124
rect	492	124	493	125
rect	492	125	493	126
rect	492	126	493	127
rect	492	127	493	128
rect	492	128	493	129
rect	492	129	493	130
rect	492	130	493	131
rect	492	131	493	132
rect	492	132	493	133
rect	492	133	493	134
rect	492	134	493	135
rect	492	135	493	136
rect	492	136	493	137
rect	492	137	493	138
rect	492	138	493	139
rect	492	139	493	140
rect	492	140	493	141
rect	492	141	493	142
rect	492	142	493	143
rect	492	143	493	144
rect	492	144	493	145
rect	492	145	493	146
rect	492	146	493	147
rect	492	147	493	148
rect	492	148	493	149
rect	492	149	493	150
rect	492	150	493	151
rect	492	151	493	152
rect	492	152	493	153
rect	492	153	493	154
rect	492	154	493	155
rect	492	155	493	156
rect	492	156	493	157
rect	492	157	493	158
rect	492	158	493	159
rect	492	159	493	160
rect	492	160	493	161
rect	492	161	493	162
rect	492	162	493	163
rect	492	163	493	164
rect	492	164	493	165
rect	492	165	493	166
rect	492	166	493	167
rect	492	167	493	168
rect	492	168	493	169
rect	492	169	493	170
rect	492	170	493	171
rect	492	171	493	172
rect	492	172	493	173
rect	492	173	493	174
rect	492	174	493	175
rect	492	175	493	176
rect	492	176	493	177
rect	492	177	493	178
rect	492	178	493	179
rect	492	179	493	180
rect	492	180	493	181
rect	492	181	493	182
rect	492	182	493	183
rect	492	183	493	184
rect	492	184	493	185
rect	492	185	493	186
rect	492	186	493	187
rect	492	187	493	188
rect	492	188	493	189
rect	492	189	493	190
rect	492	190	493	191
rect	492	191	493	192
rect	492	192	493	193
rect	492	193	493	194
rect	492	194	493	195
rect	492	195	493	196
rect	492	196	493	197
rect	492	197	493	198
rect	492	198	493	199
rect	492	199	493	200
rect	492	200	493	201
rect	492	201	493	202
rect	492	202	493	203
rect	492	203	493	204
rect	492	204	493	205
rect	492	205	493	206
rect	492	206	493	207
rect	492	207	493	208
rect	492	208	493	209
rect	492	209	493	210
rect	492	210	493	211
rect	492	211	493	212
rect	492	212	493	213
rect	492	213	493	214
rect	492	214	493	215
rect	492	215	493	216
rect	492	216	493	217
rect	492	217	493	218
rect	492	218	493	219
rect	492	219	493	220
rect	492	220	493	221
rect	492	221	493	222
rect	492	222	493	223
rect	492	223	493	224
rect	492	224	493	225
rect	492	225	493	226
rect	492	226	493	227
rect	492	227	493	228
rect	492	228	493	229
rect	492	229	493	230
rect	492	230	493	231
rect	492	231	493	232
rect	492	232	493	233
rect	492	233	493	234
rect	492	234	493	235
rect	492	235	493	236
rect	492	236	493	237
rect	492	237	493	238
rect	492	238	493	239
rect	492	239	493	240
rect	492	240	493	241
rect	492	241	493	242
rect	492	242	493	243
rect	492	243	493	244
rect	492	244	493	245
rect	492	245	493	246
rect	492	246	493	247
rect	492	247	493	248
rect	492	248	493	249
rect	492	249	493	250
rect	492	250	493	251
rect	492	251	493	252
rect	492	252	493	253
rect	492	253	493	254
rect	492	254	493	255
rect	492	255	493	256
rect	492	256	493	257
rect	492	257	493	258
rect	492	258	493	259
rect	492	259	493	260
rect	492	260	493	261
rect	492	261	493	262
rect	492	262	493	263
rect	492	263	493	264
rect	492	264	493	265
rect	492	265	493	266
rect	492	266	493	267
rect	492	267	493	268
rect	492	268	493	269
rect	492	269	493	270
rect	492	270	493	271
rect	492	271	493	272
rect	492	272	493	273
rect	492	273	493	274
rect	492	274	493	275
rect	492	275	493	276
rect	492	276	493	277
rect	492	277	493	278
rect	492	278	493	279
rect	492	279	493	280
rect	492	280	493	281
rect	492	281	493	282
rect	492	282	493	283
rect	492	283	493	284
rect	492	284	493	285
rect	492	285	493	286
rect	492	286	493	287
rect	492	287	493	288
rect	492	288	493	289
rect	492	289	493	290
rect	492	290	493	291
rect	492	291	493	292
rect	492	292	493	293
rect	492	293	493	294
rect	492	294	493	295
rect	492	295	493	296
rect	492	296	493	297
rect	492	297	493	298
rect	492	298	493	299
rect	492	299	493	300
rect	492	300	493	301
rect	492	301	493	302
rect	492	302	493	303
rect	492	303	493	304
rect	492	304	493	305
rect	492	305	493	306
rect	492	306	493	307
rect	492	307	493	308
rect	492	308	493	309
rect	492	309	493	310
rect	492	310	493	311
rect	492	311	493	312
rect	492	312	493	313
rect	492	313	493	314
rect	492	314	493	315
rect	492	315	493	316
rect	492	316	493	317
rect	492	317	493	318
rect	492	318	493	319
rect	492	319	493	320
rect	492	320	493	321
rect	493	0	494	1
rect	493	1	494	2
rect	493	2	494	3
rect	493	3	494	4
rect	493	4	494	5
rect	493	5	494	6
rect	493	6	494	7
rect	493	7	494	8
rect	493	8	494	9
rect	493	9	494	10
rect	493	10	494	11
rect	493	11	494	12
rect	493	12	494	13
rect	493	13	494	14
rect	493	14	494	15
rect	493	15	494	16
rect	493	16	494	17
rect	493	17	494	18
rect	493	18	494	19
rect	493	19	494	20
rect	493	20	494	21
rect	493	21	494	22
rect	493	22	494	23
rect	493	23	494	24
rect	493	24	494	25
rect	493	25	494	26
rect	493	26	494	27
rect	493	27	494	28
rect	493	28	494	29
rect	493	29	494	30
rect	493	30	494	31
rect	493	31	494	32
rect	493	32	494	33
rect	493	33	494	34
rect	493	34	494	35
rect	493	35	494	36
rect	493	36	494	37
rect	493	37	494	38
rect	493	38	494	39
rect	493	39	494	40
rect	493	40	494	41
rect	493	41	494	42
rect	493	42	494	43
rect	493	43	494	44
rect	493	44	494	45
rect	493	45	494	46
rect	493	46	494	47
rect	493	47	494	48
rect	493	48	494	49
rect	493	49	494	50
rect	493	50	494	51
rect	493	51	494	52
rect	493	52	494	53
rect	493	53	494	54
rect	493	54	494	55
rect	493	55	494	56
rect	493	56	494	57
rect	493	57	494	58
rect	493	58	494	59
rect	493	59	494	60
rect	493	60	494	61
rect	493	61	494	62
rect	493	62	494	63
rect	493	63	494	64
rect	493	64	494	65
rect	493	65	494	66
rect	493	66	494	67
rect	493	67	494	68
rect	493	68	494	69
rect	493	69	494	70
rect	493	70	494	71
rect	493	71	494	72
rect	493	72	494	73
rect	493	73	494	74
rect	493	74	494	75
rect	493	75	494	76
rect	493	76	494	77
rect	493	77	494	78
rect	493	78	494	79
rect	493	79	494	80
rect	493	80	494	81
rect	493	81	494	82
rect	493	82	494	83
rect	493	83	494	84
rect	493	84	494	85
rect	493	85	494	86
rect	493	86	494	87
rect	493	87	494	88
rect	493	88	494	89
rect	493	89	494	90
rect	493	90	494	91
rect	493	91	494	92
rect	493	92	494	93
rect	493	93	494	94
rect	493	94	494	95
rect	493	95	494	96
rect	493	96	494	97
rect	493	97	494	98
rect	493	98	494	99
rect	493	99	494	100
rect	493	100	494	101
rect	493	101	494	102
rect	493	102	494	103
rect	493	103	494	104
rect	493	104	494	105
rect	493	105	494	106
rect	493	106	494	107
rect	493	107	494	108
rect	493	108	494	109
rect	493	109	494	110
rect	493	110	494	111
rect	493	111	494	112
rect	493	112	494	113
rect	493	113	494	114
rect	493	114	494	115
rect	493	115	494	116
rect	493	116	494	117
rect	493	117	494	118
rect	493	118	494	119
rect	493	119	494	120
rect	493	120	494	121
rect	493	121	494	122
rect	493	122	494	123
rect	493	123	494	124
rect	493	124	494	125
rect	493	125	494	126
rect	493	126	494	127
rect	493	127	494	128
rect	493	128	494	129
rect	493	129	494	130
rect	493	130	494	131
rect	493	131	494	132
rect	493	132	494	133
rect	493	133	494	134
rect	493	134	494	135
rect	493	135	494	136
rect	493	136	494	137
rect	493	137	494	138
rect	493	138	494	139
rect	493	139	494	140
rect	493	140	494	141
rect	493	141	494	142
rect	493	142	494	143
rect	493	143	494	144
rect	493	144	494	145
rect	493	145	494	146
rect	493	146	494	147
rect	493	147	494	148
rect	493	148	494	149
rect	493	149	494	150
rect	493	150	494	151
rect	493	151	494	152
rect	493	152	494	153
rect	493	153	494	154
rect	493	154	494	155
rect	493	155	494	156
rect	493	156	494	157
rect	493	157	494	158
rect	493	158	494	159
rect	493	159	494	160
rect	493	160	494	161
rect	493	161	494	162
rect	493	162	494	163
rect	493	163	494	164
rect	493	164	494	165
rect	493	165	494	166
rect	493	166	494	167
rect	493	167	494	168
rect	493	168	494	169
rect	493	169	494	170
rect	493	170	494	171
rect	493	171	494	172
rect	493	172	494	173
rect	493	173	494	174
rect	493	174	494	175
rect	493	175	494	176
rect	493	176	494	177
rect	493	177	494	178
rect	493	178	494	179
rect	493	179	494	180
rect	493	180	494	181
rect	493	181	494	182
rect	493	182	494	183
rect	493	183	494	184
rect	493	184	494	185
rect	493	185	494	186
rect	493	186	494	187
rect	493	187	494	188
rect	493	188	494	189
rect	493	189	494	190
rect	493	190	494	191
rect	493	191	494	192
rect	493	192	494	193
rect	493	193	494	194
rect	493	194	494	195
rect	493	195	494	196
rect	493	196	494	197
rect	493	197	494	198
rect	493	198	494	199
rect	493	199	494	200
rect	493	200	494	201
rect	493	201	494	202
rect	493	202	494	203
rect	493	203	494	204
rect	493	204	494	205
rect	493	205	494	206
rect	493	206	494	207
rect	493	207	494	208
rect	493	208	494	209
rect	493	209	494	210
rect	493	210	494	211
rect	493	211	494	212
rect	493	212	494	213
rect	493	213	494	214
rect	493	214	494	215
rect	493	215	494	216
rect	493	216	494	217
rect	493	217	494	218
rect	493	218	494	219
rect	493	219	494	220
rect	493	220	494	221
rect	493	221	494	222
rect	493	222	494	223
rect	493	223	494	224
rect	493	224	494	225
rect	493	225	494	226
rect	493	226	494	227
rect	493	227	494	228
rect	493	228	494	229
rect	493	229	494	230
rect	493	230	494	231
rect	493	231	494	232
rect	493	232	494	233
rect	493	233	494	234
rect	493	234	494	235
rect	493	235	494	236
rect	493	236	494	237
rect	493	237	494	238
rect	493	238	494	239
rect	493	239	494	240
rect	493	240	494	241
rect	493	241	494	242
rect	493	242	494	243
rect	493	243	494	244
rect	493	244	494	245
rect	493	245	494	246
rect	493	246	494	247
rect	493	247	494	248
rect	493	248	494	249
rect	493	249	494	250
rect	493	250	494	251
rect	493	251	494	252
rect	493	252	494	253
rect	493	253	494	254
rect	493	254	494	255
rect	493	255	494	256
rect	493	256	494	257
rect	493	257	494	258
rect	493	258	494	259
rect	493	259	494	260
rect	493	260	494	261
rect	493	261	494	262
rect	493	262	494	263
rect	493	263	494	264
rect	493	264	494	265
rect	493	265	494	266
rect	493	266	494	267
rect	493	267	494	268
rect	493	268	494	269
rect	493	269	494	270
rect	493	270	494	271
rect	493	271	494	272
rect	493	272	494	273
rect	493	273	494	274
rect	493	274	494	275
rect	493	275	494	276
rect	493	276	494	277
rect	493	277	494	278
rect	493	278	494	279
rect	493	279	494	280
rect	493	280	494	281
rect	493	281	494	282
rect	493	282	494	283
rect	493	283	494	284
rect	493	284	494	285
rect	493	285	494	286
rect	493	286	494	287
rect	493	287	494	288
rect	493	288	494	289
rect	493	289	494	290
rect	493	290	494	291
rect	493	291	494	292
rect	493	292	494	293
rect	493	293	494	294
rect	493	294	494	295
rect	493	295	494	296
rect	493	296	494	297
rect	493	297	494	298
rect	493	298	494	299
rect	493	299	494	300
rect	493	300	494	301
rect	493	301	494	302
rect	493	302	494	303
rect	493	303	494	304
rect	493	304	494	305
rect	493	305	494	306
rect	493	306	494	307
rect	493	307	494	308
rect	493	308	494	309
rect	493	309	494	310
rect	493	310	494	311
rect	493	311	494	312
rect	493	312	494	313
rect	493	313	494	314
rect	493	314	494	315
rect	493	315	494	316
rect	493	316	494	317
rect	493	317	494	318
rect	493	318	494	319
rect	493	319	494	320
rect	493	320	494	321
rect	494	0	495	1
rect	494	1	495	2
rect	494	2	495	3
rect	494	3	495	4
rect	494	4	495	5
rect	494	5	495	6
rect	494	6	495	7
rect	494	7	495	8
rect	494	8	495	9
rect	494	9	495	10
rect	494	10	495	11
rect	494	11	495	12
rect	494	12	495	13
rect	494	13	495	14
rect	494	14	495	15
rect	494	15	495	16
rect	494	16	495	17
rect	494	17	495	18
rect	494	18	495	19
rect	494	19	495	20
rect	494	20	495	21
rect	494	21	495	22
rect	494	22	495	23
rect	494	23	495	24
rect	494	24	495	25
rect	494	25	495	26
rect	494	26	495	27
rect	494	27	495	28
rect	494	28	495	29
rect	494	29	495	30
rect	494	30	495	31
rect	494	31	495	32
rect	494	32	495	33
rect	494	33	495	34
rect	494	34	495	35
rect	494	35	495	36
rect	494	36	495	37
rect	494	37	495	38
rect	494	38	495	39
rect	494	39	495	40
rect	494	40	495	41
rect	494	41	495	42
rect	494	42	495	43
rect	494	43	495	44
rect	494	44	495	45
rect	494	45	495	46
rect	494	46	495	47
rect	494	47	495	48
rect	494	48	495	49
rect	494	49	495	50
rect	494	50	495	51
rect	494	51	495	52
rect	494	52	495	53
rect	494	53	495	54
rect	494	54	495	55
rect	494	55	495	56
rect	494	56	495	57
rect	494	57	495	58
rect	494	58	495	59
rect	494	59	495	60
rect	494	60	495	61
rect	494	61	495	62
rect	494	62	495	63
rect	494	63	495	64
rect	494	64	495	65
rect	494	65	495	66
rect	494	66	495	67
rect	494	67	495	68
rect	494	68	495	69
rect	494	69	495	70
rect	494	70	495	71
rect	494	71	495	72
rect	494	72	495	73
rect	494	73	495	74
rect	494	74	495	75
rect	494	75	495	76
rect	494	76	495	77
rect	494	77	495	78
rect	494	78	495	79
rect	494	79	495	80
rect	494	80	495	81
rect	494	81	495	82
rect	494	82	495	83
rect	494	83	495	84
rect	494	84	495	85
rect	494	85	495	86
rect	494	86	495	87
rect	494	87	495	88
rect	494	88	495	89
rect	494	89	495	90
rect	494	90	495	91
rect	494	91	495	92
rect	494	92	495	93
rect	494	93	495	94
rect	494	94	495	95
rect	494	95	495	96
rect	494	96	495	97
rect	494	97	495	98
rect	494	98	495	99
rect	494	99	495	100
rect	494	100	495	101
rect	494	101	495	102
rect	494	102	495	103
rect	494	103	495	104
rect	494	104	495	105
rect	494	105	495	106
rect	494	106	495	107
rect	494	107	495	108
rect	494	108	495	109
rect	494	109	495	110
rect	494	110	495	111
rect	494	111	495	112
rect	494	112	495	113
rect	494	113	495	114
rect	494	114	495	115
rect	494	115	495	116
rect	494	116	495	117
rect	494	117	495	118
rect	494	118	495	119
rect	494	119	495	120
rect	494	120	495	121
rect	494	121	495	122
rect	494	122	495	123
rect	494	123	495	124
rect	494	124	495	125
rect	494	125	495	126
rect	494	126	495	127
rect	494	127	495	128
rect	494	128	495	129
rect	494	129	495	130
rect	494	130	495	131
rect	494	131	495	132
rect	494	132	495	133
rect	494	133	495	134
rect	494	134	495	135
rect	494	135	495	136
rect	494	136	495	137
rect	494	137	495	138
rect	494	138	495	139
rect	494	139	495	140
rect	494	140	495	141
rect	494	141	495	142
rect	494	142	495	143
rect	494	143	495	144
rect	494	144	495	145
rect	494	145	495	146
rect	494	146	495	147
rect	494	147	495	148
rect	494	148	495	149
rect	494	149	495	150
rect	494	150	495	151
rect	494	151	495	152
rect	494	152	495	153
rect	494	153	495	154
rect	494	154	495	155
rect	494	155	495	156
rect	494	156	495	157
rect	494	157	495	158
rect	494	158	495	159
rect	494	159	495	160
rect	494	160	495	161
rect	494	161	495	162
rect	494	162	495	163
rect	494	163	495	164
rect	494	164	495	165
rect	494	165	495	166
rect	494	166	495	167
rect	494	167	495	168
rect	494	168	495	169
rect	494	169	495	170
rect	494	170	495	171
rect	494	171	495	172
rect	494	172	495	173
rect	494	173	495	174
rect	494	174	495	175
rect	494	175	495	176
rect	494	176	495	177
rect	494	177	495	178
rect	494	178	495	179
rect	494	179	495	180
rect	494	180	495	181
rect	494	181	495	182
rect	494	182	495	183
rect	494	183	495	184
rect	494	184	495	185
rect	494	185	495	186
rect	494	186	495	187
rect	494	187	495	188
rect	494	188	495	189
rect	494	189	495	190
rect	494	190	495	191
rect	494	191	495	192
rect	494	192	495	193
rect	494	193	495	194
rect	494	194	495	195
rect	494	195	495	196
rect	494	196	495	197
rect	494	197	495	198
rect	494	198	495	199
rect	494	199	495	200
rect	494	200	495	201
rect	494	201	495	202
rect	494	202	495	203
rect	494	203	495	204
rect	494	204	495	205
rect	494	205	495	206
rect	494	206	495	207
rect	494	207	495	208
rect	494	208	495	209
rect	494	209	495	210
rect	494	210	495	211
rect	494	211	495	212
rect	494	212	495	213
rect	494	213	495	214
rect	494	214	495	215
rect	494	215	495	216
rect	494	216	495	217
rect	494	217	495	218
rect	494	218	495	219
rect	494	219	495	220
rect	494	220	495	221
rect	494	221	495	222
rect	494	222	495	223
rect	494	223	495	224
rect	494	224	495	225
rect	494	225	495	226
rect	494	226	495	227
rect	494	227	495	228
rect	494	228	495	229
rect	494	229	495	230
rect	494	230	495	231
rect	494	231	495	232
rect	494	232	495	233
rect	494	233	495	234
rect	494	234	495	235
rect	494	235	495	236
rect	494	236	495	237
rect	494	237	495	238
rect	494	238	495	239
rect	494	239	495	240
rect	494	240	495	241
rect	494	241	495	242
rect	494	242	495	243
rect	494	243	495	244
rect	494	244	495	245
rect	494	245	495	246
rect	494	246	495	247
rect	494	247	495	248
rect	494	248	495	249
rect	494	249	495	250
rect	494	250	495	251
rect	494	251	495	252
rect	494	252	495	253
rect	494	253	495	254
rect	494	254	495	255
rect	494	255	495	256
rect	494	256	495	257
rect	494	257	495	258
rect	494	258	495	259
rect	494	259	495	260
rect	494	260	495	261
rect	494	261	495	262
rect	494	262	495	263
rect	494	263	495	264
rect	494	264	495	265
rect	494	265	495	266
rect	494	266	495	267
rect	494	267	495	268
rect	494	268	495	269
rect	494	269	495	270
rect	494	270	495	271
rect	494	271	495	272
rect	494	272	495	273
rect	494	273	495	274
rect	494	274	495	275
rect	494	275	495	276
rect	494	276	495	277
rect	494	277	495	278
rect	494	278	495	279
rect	494	279	495	280
rect	494	280	495	281
rect	494	281	495	282
rect	494	282	495	283
rect	494	283	495	284
rect	494	284	495	285
rect	494	285	495	286
rect	494	286	495	287
rect	494	287	495	288
rect	494	288	495	289
rect	494	289	495	290
rect	494	290	495	291
rect	494	291	495	292
rect	494	292	495	293
rect	494	293	495	294
rect	494	294	495	295
rect	494	295	495	296
rect	494	296	495	297
rect	494	297	495	298
rect	494	298	495	299
rect	494	299	495	300
rect	494	300	495	301
rect	494	301	495	302
rect	494	302	495	303
rect	494	303	495	304
rect	494	304	495	305
rect	494	305	495	306
rect	494	306	495	307
rect	494	307	495	308
rect	494	308	495	309
rect	494	309	495	310
rect	494	310	495	311
rect	494	311	495	312
rect	494	312	495	313
rect	494	313	495	314
rect	494	314	495	315
rect	494	315	495	316
rect	494	316	495	317
rect	494	317	495	318
rect	494	318	495	319
rect	494	319	495	320
rect	494	320	495	321
rect	524	0	525	1
rect	524	1	525	2
rect	524	2	525	3
rect	524	3	525	4
rect	524	4	525	5
rect	524	5	525	6
rect	524	6	525	7
rect	524	7	525	8
rect	524	8	525	9
rect	524	9	525	10
rect	524	10	525	11
rect	524	11	525	12
rect	524	12	525	13
rect	524	13	525	14
rect	524	14	525	15
rect	524	15	525	16
rect	524	16	525	17
rect	524	17	525	18
rect	524	18	525	19
rect	524	19	525	20
rect	524	20	525	21
rect	524	21	525	22
rect	524	22	525	23
rect	524	23	525	24
rect	524	24	525	25
rect	524	25	525	26
rect	524	26	525	27
rect	524	27	525	28
rect	524	28	525	29
rect	524	29	525	30
rect	524	30	525	31
rect	524	31	525	32
rect	524	32	525	33
rect	524	33	525	34
rect	524	34	525	35
rect	524	35	525	36
rect	524	36	525	37
rect	524	37	525	38
rect	524	38	525	39
rect	524	39	525	40
rect	524	40	525	41
rect	524	41	525	42
rect	524	42	525	43
rect	524	43	525	44
rect	524	44	525	45
rect	524	45	525	46
rect	524	46	525	47
rect	524	47	525	48
rect	524	48	525	49
rect	524	49	525	50
rect	524	50	525	51
rect	524	51	525	52
rect	524	52	525	53
rect	524	53	525	54
rect	524	54	525	55
rect	524	55	525	56
rect	524	56	525	57
rect	524	57	525	58
rect	524	58	525	59
rect	524	59	525	60
rect	524	60	525	61
rect	524	61	525	62
rect	524	62	525	63
rect	524	63	525	64
rect	524	64	525	65
rect	524	65	525	66
rect	524	66	525	67
rect	524	67	525	68
rect	524	68	525	69
rect	524	69	525	70
rect	524	70	525	71
rect	524	71	525	72
rect	524	72	525	73
rect	524	73	525	74
rect	524	74	525	75
rect	524	75	525	76
rect	524	76	525	77
rect	524	77	525	78
rect	524	78	525	79
rect	524	79	525	80
rect	524	80	525	81
rect	524	81	525	82
rect	524	82	525	83
rect	524	83	525	84
rect	524	84	525	85
rect	524	85	525	86
rect	524	86	525	87
rect	524	87	525	88
rect	524	88	525	89
rect	524	89	525	90
rect	524	90	525	91
rect	524	91	525	92
rect	524	92	525	93
rect	524	93	525	94
rect	524	94	525	95
rect	524	95	525	96
rect	524	96	525	97
rect	524	97	525	98
rect	524	98	525	99
rect	524	99	525	100
rect	524	100	525	101
rect	524	101	525	102
rect	524	102	525	103
rect	524	103	525	104
rect	524	104	525	105
rect	524	105	525	106
rect	524	106	525	107
rect	524	107	525	108
rect	524	108	525	109
rect	524	109	525	110
rect	524	110	525	111
rect	524	111	525	112
rect	524	112	525	113
rect	524	113	525	114
rect	524	114	525	115
rect	524	115	525	116
rect	524	116	525	117
rect	524	117	525	118
rect	524	118	525	119
rect	524	119	525	120
rect	524	120	525	121
rect	524	121	525	122
rect	524	122	525	123
rect	524	123	525	124
rect	524	124	525	125
rect	524	125	525	126
rect	524	126	525	127
rect	524	127	525	128
rect	524	128	525	129
rect	524	129	525	130
rect	524	130	525	131
rect	524	131	525	132
rect	524	132	525	133
rect	524	133	525	134
rect	524	134	525	135
rect	524	135	525	136
rect	524	136	525	137
rect	524	137	525	138
rect	524	138	525	139
rect	524	139	525	140
rect	524	140	525	141
rect	524	141	525	142
rect	524	142	525	143
rect	524	143	525	144
rect	524	144	525	145
rect	524	145	525	146
rect	524	146	525	147
rect	524	147	525	148
rect	524	148	525	149
rect	524	149	525	150
rect	524	150	525	151
rect	524	151	525	152
rect	524	152	525	153
rect	524	153	525	154
rect	524	154	525	155
rect	524	155	525	156
rect	524	156	525	157
rect	524	157	525	158
rect	524	158	525	159
rect	524	159	525	160
rect	524	160	525	161
rect	524	161	525	162
rect	524	162	525	163
rect	524	163	525	164
rect	524	164	525	165
rect	524	165	525	166
rect	524	166	525	167
rect	524	167	525	168
rect	524	168	525	169
rect	524	169	525	170
rect	524	170	525	171
rect	524	171	525	172
rect	524	172	525	173
rect	524	173	525	174
rect	524	174	525	175
rect	524	175	525	176
rect	524	176	525	177
rect	524	177	525	178
rect	524	178	525	179
rect	524	179	525	180
rect	524	180	525	181
rect	524	181	525	182
rect	524	182	525	183
rect	524	183	525	184
rect	524	184	525	185
rect	524	185	525	186
rect	524	186	525	187
rect	524	187	525	188
rect	524	188	525	189
rect	524	189	525	190
rect	524	190	525	191
rect	524	191	525	192
rect	524	192	525	193
rect	524	193	525	194
rect	524	194	525	195
rect	524	195	525	196
rect	524	196	525	197
rect	524	197	525	198
rect	524	198	525	199
rect	524	199	525	200
rect	524	200	525	201
rect	524	201	525	202
rect	524	202	525	203
rect	524	203	525	204
rect	524	204	525	205
rect	524	205	525	206
rect	524	206	525	207
rect	524	207	525	208
rect	524	208	525	209
rect	524	209	525	210
rect	524	210	525	211
rect	524	211	525	212
rect	524	212	525	213
rect	524	213	525	214
rect	524	214	525	215
rect	524	215	525	216
rect	524	216	525	217
rect	524	217	525	218
rect	524	218	525	219
rect	524	219	525	220
rect	524	220	525	221
rect	524	221	525	222
rect	524	222	525	223
rect	524	223	525	224
rect	524	224	525	225
rect	524	225	525	226
rect	524	226	525	227
rect	524	227	525	228
rect	524	228	525	229
rect	524	229	525	230
rect	524	230	525	231
rect	524	231	525	232
rect	524	232	525	233
rect	524	233	525	234
rect	524	234	525	235
rect	524	235	525	236
rect	524	236	525	237
rect	524	237	525	238
rect	524	238	525	239
rect	524	239	525	240
rect	524	240	525	241
rect	524	241	525	242
rect	524	242	525	243
rect	524	243	525	244
rect	524	244	525	245
rect	524	245	525	246
rect	524	246	525	247
rect	524	247	525	248
rect	524	248	525	249
rect	524	249	525	250
rect	524	250	525	251
rect	524	251	525	252
rect	524	252	525	253
rect	524	253	525	254
rect	524	254	525	255
rect	524	255	525	256
rect	524	256	525	257
rect	524	257	525	258
rect	524	258	525	259
rect	524	259	525	260
rect	524	260	525	261
rect	524	261	525	262
rect	524	262	525	263
rect	524	263	525	264
rect	524	264	525	265
rect	524	265	525	266
rect	524	266	525	267
rect	524	267	525	268
rect	524	268	525	269
rect	524	269	525	270
rect	524	270	525	271
rect	524	271	525	272
rect	524	272	525	273
rect	524	273	525	274
rect	524	274	525	275
rect	524	275	525	276
rect	524	276	525	277
rect	524	277	525	278
rect	524	278	525	279
rect	524	279	525	280
rect	524	280	525	281
rect	524	281	525	282
rect	524	282	525	283
rect	524	283	525	284
rect	524	284	525	285
rect	524	285	525	286
rect	524	286	525	287
rect	524	287	525	288
rect	525	0	526	1
rect	525	1	526	2
rect	525	2	526	3
rect	525	3	526	4
rect	525	4	526	5
rect	525	5	526	6
rect	525	6	526	7
rect	525	7	526	8
rect	525	8	526	9
rect	525	9	526	10
rect	525	10	526	11
rect	525	11	526	12
rect	525	12	526	13
rect	525	13	526	14
rect	525	14	526	15
rect	525	15	526	16
rect	525	16	526	17
rect	525	17	526	18
rect	525	18	526	19
rect	525	19	526	20
rect	525	20	526	21
rect	525	21	526	22
rect	525	22	526	23
rect	525	23	526	24
rect	525	24	526	25
rect	525	25	526	26
rect	525	26	526	27
rect	525	27	526	28
rect	525	28	526	29
rect	525	29	526	30
rect	525	30	526	31
rect	525	31	526	32
rect	525	32	526	33
rect	525	33	526	34
rect	525	34	526	35
rect	525	35	526	36
rect	525	36	526	37
rect	525	37	526	38
rect	525	38	526	39
rect	525	39	526	40
rect	525	40	526	41
rect	525	41	526	42
rect	525	42	526	43
rect	525	43	526	44
rect	525	44	526	45
rect	525	45	526	46
rect	525	46	526	47
rect	525	47	526	48
rect	525	48	526	49
rect	525	49	526	50
rect	525	50	526	51
rect	525	51	526	52
rect	525	52	526	53
rect	525	53	526	54
rect	525	54	526	55
rect	525	55	526	56
rect	525	56	526	57
rect	525	57	526	58
rect	525	58	526	59
rect	525	59	526	60
rect	525	60	526	61
rect	525	61	526	62
rect	525	62	526	63
rect	525	63	526	64
rect	525	64	526	65
rect	525	65	526	66
rect	525	66	526	67
rect	525	67	526	68
rect	525	68	526	69
rect	525	69	526	70
rect	525	70	526	71
rect	525	71	526	72
rect	525	72	526	73
rect	525	73	526	74
rect	525	74	526	75
rect	525	75	526	76
rect	525	76	526	77
rect	525	77	526	78
rect	525	78	526	79
rect	525	79	526	80
rect	525	80	526	81
rect	525	81	526	82
rect	525	82	526	83
rect	525	83	526	84
rect	525	84	526	85
rect	525	85	526	86
rect	525	86	526	87
rect	525	87	526	88
rect	525	88	526	89
rect	525	89	526	90
rect	525	90	526	91
rect	525	91	526	92
rect	525	92	526	93
rect	525	93	526	94
rect	525	94	526	95
rect	525	95	526	96
rect	525	96	526	97
rect	525	97	526	98
rect	525	98	526	99
rect	525	99	526	100
rect	525	100	526	101
rect	525	101	526	102
rect	525	102	526	103
rect	525	103	526	104
rect	525	104	526	105
rect	525	105	526	106
rect	525	106	526	107
rect	525	107	526	108
rect	525	108	526	109
rect	525	109	526	110
rect	525	110	526	111
rect	525	111	526	112
rect	525	112	526	113
rect	525	113	526	114
rect	525	114	526	115
rect	525	115	526	116
rect	525	116	526	117
rect	525	117	526	118
rect	525	118	526	119
rect	525	119	526	120
rect	525	120	526	121
rect	525	121	526	122
rect	525	122	526	123
rect	525	123	526	124
rect	525	124	526	125
rect	525	125	526	126
rect	525	126	526	127
rect	525	127	526	128
rect	525	128	526	129
rect	525	129	526	130
rect	525	130	526	131
rect	525	131	526	132
rect	525	132	526	133
rect	525	133	526	134
rect	525	134	526	135
rect	525	135	526	136
rect	525	136	526	137
rect	525	137	526	138
rect	525	138	526	139
rect	525	139	526	140
rect	525	140	526	141
rect	525	141	526	142
rect	525	142	526	143
rect	525	143	526	144
rect	525	144	526	145
rect	525	145	526	146
rect	525	146	526	147
rect	525	147	526	148
rect	525	148	526	149
rect	525	149	526	150
rect	525	150	526	151
rect	525	151	526	152
rect	525	152	526	153
rect	525	153	526	154
rect	525	154	526	155
rect	525	155	526	156
rect	525	156	526	157
rect	525	157	526	158
rect	525	158	526	159
rect	525	159	526	160
rect	525	160	526	161
rect	525	161	526	162
rect	525	162	526	163
rect	525	163	526	164
rect	525	164	526	165
rect	525	165	526	166
rect	525	166	526	167
rect	525	167	526	168
rect	525	168	526	169
rect	525	169	526	170
rect	525	170	526	171
rect	525	171	526	172
rect	525	172	526	173
rect	525	173	526	174
rect	525	174	526	175
rect	525	175	526	176
rect	525	176	526	177
rect	525	177	526	178
rect	525	178	526	179
rect	525	179	526	180
rect	525	180	526	181
rect	525	181	526	182
rect	525	182	526	183
rect	525	183	526	184
rect	525	184	526	185
rect	525	185	526	186
rect	525	186	526	187
rect	525	187	526	188
rect	525	188	526	189
rect	525	189	526	190
rect	525	190	526	191
rect	525	191	526	192
rect	525	192	526	193
rect	525	193	526	194
rect	525	194	526	195
rect	525	195	526	196
rect	525	196	526	197
rect	525	197	526	198
rect	525	198	526	199
rect	525	199	526	200
rect	525	200	526	201
rect	525	201	526	202
rect	525	202	526	203
rect	525	203	526	204
rect	525	204	526	205
rect	525	205	526	206
rect	525	206	526	207
rect	525	207	526	208
rect	525	208	526	209
rect	525	209	526	210
rect	525	210	526	211
rect	525	211	526	212
rect	525	212	526	213
rect	525	213	526	214
rect	525	214	526	215
rect	525	215	526	216
rect	525	216	526	217
rect	525	217	526	218
rect	525	218	526	219
rect	525	219	526	220
rect	525	220	526	221
rect	525	221	526	222
rect	525	222	526	223
rect	525	223	526	224
rect	525	224	526	225
rect	525	225	526	226
rect	525	226	526	227
rect	525	227	526	228
rect	525	228	526	229
rect	525	229	526	230
rect	525	230	526	231
rect	525	231	526	232
rect	525	232	526	233
rect	525	233	526	234
rect	525	234	526	235
rect	525	235	526	236
rect	525	236	526	237
rect	525	237	526	238
rect	525	238	526	239
rect	525	239	526	240
rect	525	240	526	241
rect	525	241	526	242
rect	525	242	526	243
rect	525	243	526	244
rect	525	244	526	245
rect	525	245	526	246
rect	525	246	526	247
rect	525	247	526	248
rect	525	248	526	249
rect	525	249	526	250
rect	525	250	526	251
rect	525	251	526	252
rect	525	252	526	253
rect	525	253	526	254
rect	525	254	526	255
rect	525	255	526	256
rect	525	256	526	257
rect	525	257	526	258
rect	525	258	526	259
rect	525	259	526	260
rect	525	260	526	261
rect	525	261	526	262
rect	525	262	526	263
rect	525	263	526	264
rect	525	264	526	265
rect	525	265	526	266
rect	525	266	526	267
rect	525	267	526	268
rect	525	268	526	269
rect	525	269	526	270
rect	525	270	526	271
rect	525	271	526	272
rect	525	272	526	273
rect	525	273	526	274
rect	525	274	526	275
rect	525	275	526	276
rect	525	276	526	277
rect	525	277	526	278
rect	525	278	526	279
rect	525	279	526	280
rect	525	280	526	281
rect	525	281	526	282
rect	525	282	526	283
rect	525	283	526	284
rect	525	284	526	285
rect	525	285	526	286
rect	525	286	526	287
rect	525	287	526	288
rect	526	0	527	1
rect	526	1	527	2
rect	526	2	527	3
rect	526	3	527	4
rect	526	4	527	5
rect	526	5	527	6
rect	526	6	527	7
rect	526	7	527	8
rect	526	8	527	9
rect	526	9	527	10
rect	526	10	527	11
rect	526	11	527	12
rect	526	12	527	13
rect	526	13	527	14
rect	526	14	527	15
rect	526	15	527	16
rect	526	16	527	17
rect	526	17	527	18
rect	526	18	527	19
rect	526	19	527	20
rect	526	20	527	21
rect	526	21	527	22
rect	526	22	527	23
rect	526	23	527	24
rect	526	24	527	25
rect	526	25	527	26
rect	526	26	527	27
rect	526	27	527	28
rect	526	28	527	29
rect	526	29	527	30
rect	526	30	527	31
rect	526	31	527	32
rect	526	32	527	33
rect	526	33	527	34
rect	526	34	527	35
rect	526	35	527	36
rect	526	36	527	37
rect	526	37	527	38
rect	526	38	527	39
rect	526	39	527	40
rect	526	40	527	41
rect	526	41	527	42
rect	526	42	527	43
rect	526	43	527	44
rect	526	44	527	45
rect	526	45	527	46
rect	526	46	527	47
rect	526	47	527	48
rect	526	48	527	49
rect	526	49	527	50
rect	526	50	527	51
rect	526	51	527	52
rect	526	52	527	53
rect	526	53	527	54
rect	526	54	527	55
rect	526	55	527	56
rect	526	56	527	57
rect	526	57	527	58
rect	526	58	527	59
rect	526	59	527	60
rect	526	60	527	61
rect	526	61	527	62
rect	526	62	527	63
rect	526	63	527	64
rect	526	64	527	65
rect	526	65	527	66
rect	526	66	527	67
rect	526	67	527	68
rect	526	68	527	69
rect	526	69	527	70
rect	526	70	527	71
rect	526	71	527	72
rect	526	72	527	73
rect	526	73	527	74
rect	526	74	527	75
rect	526	75	527	76
rect	526	76	527	77
rect	526	77	527	78
rect	526	78	527	79
rect	526	79	527	80
rect	526	80	527	81
rect	526	81	527	82
rect	526	82	527	83
rect	526	83	527	84
rect	526	84	527	85
rect	526	85	527	86
rect	526	86	527	87
rect	526	87	527	88
rect	526	88	527	89
rect	526	89	527	90
rect	526	90	527	91
rect	526	91	527	92
rect	526	92	527	93
rect	526	93	527	94
rect	526	94	527	95
rect	526	95	527	96
rect	526	96	527	97
rect	526	97	527	98
rect	526	98	527	99
rect	526	99	527	100
rect	526	100	527	101
rect	526	101	527	102
rect	526	102	527	103
rect	526	103	527	104
rect	526	104	527	105
rect	526	105	527	106
rect	526	106	527	107
rect	526	107	527	108
rect	526	108	527	109
rect	526	109	527	110
rect	526	110	527	111
rect	526	111	527	112
rect	526	112	527	113
rect	526	113	527	114
rect	526	114	527	115
rect	526	115	527	116
rect	526	116	527	117
rect	526	117	527	118
rect	526	118	527	119
rect	526	119	527	120
rect	526	120	527	121
rect	526	121	527	122
rect	526	122	527	123
rect	526	123	527	124
rect	526	124	527	125
rect	526	125	527	126
rect	526	126	527	127
rect	526	127	527	128
rect	526	128	527	129
rect	526	129	527	130
rect	526	130	527	131
rect	526	131	527	132
rect	526	132	527	133
rect	526	133	527	134
rect	526	134	527	135
rect	526	135	527	136
rect	526	136	527	137
rect	526	137	527	138
rect	526	138	527	139
rect	526	139	527	140
rect	526	140	527	141
rect	526	141	527	142
rect	526	142	527	143
rect	526	143	527	144
rect	526	144	527	145
rect	526	145	527	146
rect	526	146	527	147
rect	526	147	527	148
rect	526	148	527	149
rect	526	149	527	150
rect	526	150	527	151
rect	526	151	527	152
rect	526	152	527	153
rect	526	153	527	154
rect	526	154	527	155
rect	526	155	527	156
rect	526	156	527	157
rect	526	157	527	158
rect	526	158	527	159
rect	526	159	527	160
rect	526	160	527	161
rect	526	161	527	162
rect	526	162	527	163
rect	526	163	527	164
rect	526	164	527	165
rect	526	165	527	166
rect	526	166	527	167
rect	526	167	527	168
rect	526	168	527	169
rect	526	169	527	170
rect	526	170	527	171
rect	526	171	527	172
rect	526	172	527	173
rect	526	173	527	174
rect	526	174	527	175
rect	526	175	527	176
rect	526	176	527	177
rect	526	177	527	178
rect	526	178	527	179
rect	526	179	527	180
rect	526	180	527	181
rect	526	181	527	182
rect	526	182	527	183
rect	526	183	527	184
rect	526	184	527	185
rect	526	185	527	186
rect	526	186	527	187
rect	526	187	527	188
rect	526	188	527	189
rect	526	189	527	190
rect	526	190	527	191
rect	526	191	527	192
rect	526	192	527	193
rect	526	193	527	194
rect	526	194	527	195
rect	526	195	527	196
rect	526	196	527	197
rect	526	197	527	198
rect	526	198	527	199
rect	526	199	527	200
rect	526	200	527	201
rect	526	201	527	202
rect	526	202	527	203
rect	526	203	527	204
rect	526	204	527	205
rect	526	205	527	206
rect	526	206	527	207
rect	526	207	527	208
rect	526	208	527	209
rect	526	209	527	210
rect	526	210	527	211
rect	526	211	527	212
rect	526	212	527	213
rect	526	213	527	214
rect	526	214	527	215
rect	526	215	527	216
rect	526	216	527	217
rect	526	217	527	218
rect	526	218	527	219
rect	526	219	527	220
rect	526	220	527	221
rect	526	221	527	222
rect	526	222	527	223
rect	526	223	527	224
rect	526	224	527	225
rect	526	225	527	226
rect	526	226	527	227
rect	526	227	527	228
rect	526	228	527	229
rect	526	229	527	230
rect	526	230	527	231
rect	526	231	527	232
rect	526	232	527	233
rect	526	233	527	234
rect	526	234	527	235
rect	526	235	527	236
rect	526	236	527	237
rect	526	237	527	238
rect	526	238	527	239
rect	526	239	527	240
rect	526	240	527	241
rect	526	241	527	242
rect	526	242	527	243
rect	526	243	527	244
rect	526	244	527	245
rect	526	245	527	246
rect	526	246	527	247
rect	526	247	527	248
rect	526	248	527	249
rect	526	249	527	250
rect	526	250	527	251
rect	526	251	527	252
rect	526	252	527	253
rect	526	253	527	254
rect	526	254	527	255
rect	526	255	527	256
rect	526	256	527	257
rect	526	257	527	258
rect	526	258	527	259
rect	526	259	527	260
rect	526	260	527	261
rect	526	261	527	262
rect	526	262	527	263
rect	526	263	527	264
rect	526	264	527	265
rect	526	265	527	266
rect	526	266	527	267
rect	526	267	527	268
rect	526	268	527	269
rect	526	269	527	270
rect	526	270	527	271
rect	526	271	527	272
rect	526	272	527	273
rect	526	273	527	274
rect	526	274	527	275
rect	526	275	527	276
rect	526	276	527	277
rect	526	277	527	278
rect	526	278	527	279
rect	526	279	527	280
rect	526	280	527	281
rect	526	281	527	282
rect	526	282	527	283
rect	526	283	527	284
rect	526	284	527	285
rect	526	285	527	286
rect	526	286	527	287
rect	526	287	527	288
rect	527	0	528	1
rect	527	1	528	2
rect	527	2	528	3
rect	527	3	528	4
rect	527	4	528	5
rect	527	5	528	6
rect	527	6	528	7
rect	527	7	528	8
rect	527	8	528	9
rect	527	9	528	10
rect	527	10	528	11
rect	527	11	528	12
rect	527	12	528	13
rect	527	13	528	14
rect	527	14	528	15
rect	527	15	528	16
rect	527	16	528	17
rect	527	17	528	18
rect	527	18	528	19
rect	527	19	528	20
rect	527	20	528	21
rect	527	21	528	22
rect	527	22	528	23
rect	527	23	528	24
rect	527	24	528	25
rect	527	25	528	26
rect	527	26	528	27
rect	527	27	528	28
rect	527	28	528	29
rect	527	29	528	30
rect	527	30	528	31
rect	527	31	528	32
rect	527	32	528	33
rect	527	33	528	34
rect	527	34	528	35
rect	527	35	528	36
rect	527	36	528	37
rect	527	37	528	38
rect	527	38	528	39
rect	527	39	528	40
rect	527	40	528	41
rect	527	41	528	42
rect	527	42	528	43
rect	527	43	528	44
rect	527	44	528	45
rect	527	45	528	46
rect	527	46	528	47
rect	527	47	528	48
rect	527	48	528	49
rect	527	49	528	50
rect	527	50	528	51
rect	527	51	528	52
rect	527	52	528	53
rect	527	53	528	54
rect	527	54	528	55
rect	527	55	528	56
rect	527	56	528	57
rect	527	57	528	58
rect	527	58	528	59
rect	527	59	528	60
rect	527	60	528	61
rect	527	61	528	62
rect	527	62	528	63
rect	527	63	528	64
rect	527	64	528	65
rect	527	65	528	66
rect	527	66	528	67
rect	527	67	528	68
rect	527	68	528	69
rect	527	69	528	70
rect	527	70	528	71
rect	527	71	528	72
rect	527	72	528	73
rect	527	73	528	74
rect	527	74	528	75
rect	527	75	528	76
rect	527	76	528	77
rect	527	77	528	78
rect	527	78	528	79
rect	527	79	528	80
rect	527	80	528	81
rect	527	81	528	82
rect	527	82	528	83
rect	527	83	528	84
rect	527	84	528	85
rect	527	85	528	86
rect	527	86	528	87
rect	527	87	528	88
rect	527	88	528	89
rect	527	89	528	90
rect	527	90	528	91
rect	527	91	528	92
rect	527	92	528	93
rect	527	93	528	94
rect	527	94	528	95
rect	527	95	528	96
rect	527	96	528	97
rect	527	97	528	98
rect	527	98	528	99
rect	527	99	528	100
rect	527	100	528	101
rect	527	101	528	102
rect	527	102	528	103
rect	527	103	528	104
rect	527	104	528	105
rect	527	105	528	106
rect	527	106	528	107
rect	527	107	528	108
rect	527	108	528	109
rect	527	109	528	110
rect	527	110	528	111
rect	527	111	528	112
rect	527	112	528	113
rect	527	113	528	114
rect	527	114	528	115
rect	527	115	528	116
rect	527	116	528	117
rect	527	117	528	118
rect	527	118	528	119
rect	527	119	528	120
rect	527	120	528	121
rect	527	121	528	122
rect	527	122	528	123
rect	527	123	528	124
rect	527	124	528	125
rect	527	125	528	126
rect	527	126	528	127
rect	527	127	528	128
rect	527	128	528	129
rect	527	129	528	130
rect	527	130	528	131
rect	527	131	528	132
rect	527	132	528	133
rect	527	133	528	134
rect	527	134	528	135
rect	527	135	528	136
rect	527	136	528	137
rect	527	137	528	138
rect	527	138	528	139
rect	527	139	528	140
rect	527	140	528	141
rect	527	141	528	142
rect	527	142	528	143
rect	527	143	528	144
rect	527	144	528	145
rect	527	145	528	146
rect	527	146	528	147
rect	527	147	528	148
rect	527	148	528	149
rect	527	149	528	150
rect	527	150	528	151
rect	527	151	528	152
rect	527	152	528	153
rect	527	153	528	154
rect	527	154	528	155
rect	527	155	528	156
rect	527	156	528	157
rect	527	157	528	158
rect	527	158	528	159
rect	527	159	528	160
rect	527	160	528	161
rect	527	161	528	162
rect	527	162	528	163
rect	527	163	528	164
rect	527	164	528	165
rect	527	165	528	166
rect	527	166	528	167
rect	527	167	528	168
rect	527	168	528	169
rect	527	169	528	170
rect	527	170	528	171
rect	527	171	528	172
rect	527	172	528	173
rect	527	173	528	174
rect	527	174	528	175
rect	527	175	528	176
rect	527	176	528	177
rect	527	177	528	178
rect	527	178	528	179
rect	527	179	528	180
rect	527	180	528	181
rect	527	181	528	182
rect	527	182	528	183
rect	527	183	528	184
rect	527	184	528	185
rect	527	185	528	186
rect	527	186	528	187
rect	527	187	528	188
rect	527	188	528	189
rect	527	189	528	190
rect	527	190	528	191
rect	527	191	528	192
rect	527	192	528	193
rect	527	193	528	194
rect	527	194	528	195
rect	527	195	528	196
rect	527	196	528	197
rect	527	197	528	198
rect	527	198	528	199
rect	527	199	528	200
rect	527	200	528	201
rect	527	201	528	202
rect	527	202	528	203
rect	527	203	528	204
rect	527	204	528	205
rect	527	205	528	206
rect	527	206	528	207
rect	527	207	528	208
rect	527	208	528	209
rect	527	209	528	210
rect	527	210	528	211
rect	527	211	528	212
rect	527	212	528	213
rect	527	213	528	214
rect	527	214	528	215
rect	527	215	528	216
rect	527	216	528	217
rect	527	217	528	218
rect	527	218	528	219
rect	527	219	528	220
rect	527	220	528	221
rect	527	221	528	222
rect	527	222	528	223
rect	527	223	528	224
rect	527	224	528	225
rect	527	225	528	226
rect	527	226	528	227
rect	527	227	528	228
rect	527	228	528	229
rect	527	229	528	230
rect	527	230	528	231
rect	527	231	528	232
rect	527	232	528	233
rect	527	233	528	234
rect	527	234	528	235
rect	527	235	528	236
rect	527	236	528	237
rect	527	237	528	238
rect	527	238	528	239
rect	527	239	528	240
rect	527	240	528	241
rect	527	241	528	242
rect	527	242	528	243
rect	527	243	528	244
rect	527	244	528	245
rect	527	245	528	246
rect	527	246	528	247
rect	527	247	528	248
rect	527	248	528	249
rect	527	249	528	250
rect	527	250	528	251
rect	527	251	528	252
rect	527	252	528	253
rect	527	253	528	254
rect	527	254	528	255
rect	527	255	528	256
rect	527	256	528	257
rect	527	257	528	258
rect	527	258	528	259
rect	527	259	528	260
rect	527	260	528	261
rect	527	261	528	262
rect	527	262	528	263
rect	527	263	528	264
rect	527	264	528	265
rect	527	265	528	266
rect	527	266	528	267
rect	527	267	528	268
rect	527	268	528	269
rect	527	269	528	270
rect	527	270	528	271
rect	527	271	528	272
rect	527	272	528	273
rect	527	273	528	274
rect	527	274	528	275
rect	527	275	528	276
rect	527	276	528	277
rect	527	277	528	278
rect	527	278	528	279
rect	527	279	528	280
rect	527	280	528	281
rect	527	281	528	282
rect	527	282	528	283
rect	527	283	528	284
rect	527	284	528	285
rect	527	285	528	286
rect	527	286	528	287
rect	527	287	528	288
rect	528	0	529	1
rect	528	1	529	2
rect	528	2	529	3
rect	528	3	529	4
rect	528	4	529	5
rect	528	5	529	6
rect	528	6	529	7
rect	528	7	529	8
rect	528	8	529	9
rect	528	9	529	10
rect	528	10	529	11
rect	528	11	529	12
rect	528	12	529	13
rect	528	13	529	14
rect	528	14	529	15
rect	528	15	529	16
rect	528	16	529	17
rect	528	17	529	18
rect	528	18	529	19
rect	528	19	529	20
rect	528	20	529	21
rect	528	21	529	22
rect	528	22	529	23
rect	528	23	529	24
rect	528	24	529	25
rect	528	25	529	26
rect	528	26	529	27
rect	528	27	529	28
rect	528	28	529	29
rect	528	29	529	30
rect	528	30	529	31
rect	528	31	529	32
rect	528	32	529	33
rect	528	33	529	34
rect	528	34	529	35
rect	528	35	529	36
rect	528	36	529	37
rect	528	37	529	38
rect	528	38	529	39
rect	528	39	529	40
rect	528	40	529	41
rect	528	41	529	42
rect	528	42	529	43
rect	528	43	529	44
rect	528	44	529	45
rect	528	45	529	46
rect	528	46	529	47
rect	528	47	529	48
rect	528	48	529	49
rect	528	49	529	50
rect	528	50	529	51
rect	528	51	529	52
rect	528	52	529	53
rect	528	53	529	54
rect	528	54	529	55
rect	528	55	529	56
rect	528	56	529	57
rect	528	57	529	58
rect	528	58	529	59
rect	528	59	529	60
rect	528	60	529	61
rect	528	61	529	62
rect	528	62	529	63
rect	528	63	529	64
rect	528	64	529	65
rect	528	65	529	66
rect	528	66	529	67
rect	528	67	529	68
rect	528	68	529	69
rect	528	69	529	70
rect	528	70	529	71
rect	528	71	529	72
rect	528	72	529	73
rect	528	73	529	74
rect	528	74	529	75
rect	528	75	529	76
rect	528	76	529	77
rect	528	77	529	78
rect	528	78	529	79
rect	528	79	529	80
rect	528	80	529	81
rect	528	81	529	82
rect	528	82	529	83
rect	528	83	529	84
rect	528	84	529	85
rect	528	85	529	86
rect	528	86	529	87
rect	528	87	529	88
rect	528	88	529	89
rect	528	89	529	90
rect	528	90	529	91
rect	528	91	529	92
rect	528	92	529	93
rect	528	93	529	94
rect	528	94	529	95
rect	528	95	529	96
rect	528	96	529	97
rect	528	97	529	98
rect	528	98	529	99
rect	528	99	529	100
rect	528	100	529	101
rect	528	101	529	102
rect	528	102	529	103
rect	528	103	529	104
rect	528	104	529	105
rect	528	105	529	106
rect	528	106	529	107
rect	528	107	529	108
rect	528	108	529	109
rect	528	109	529	110
rect	528	110	529	111
rect	528	111	529	112
rect	528	112	529	113
rect	528	113	529	114
rect	528	114	529	115
rect	528	115	529	116
rect	528	116	529	117
rect	528	117	529	118
rect	528	118	529	119
rect	528	119	529	120
rect	528	120	529	121
rect	528	121	529	122
rect	528	122	529	123
rect	528	123	529	124
rect	528	124	529	125
rect	528	125	529	126
rect	528	126	529	127
rect	528	127	529	128
rect	528	128	529	129
rect	528	129	529	130
rect	528	130	529	131
rect	528	131	529	132
rect	528	132	529	133
rect	528	133	529	134
rect	528	134	529	135
rect	528	135	529	136
rect	528	136	529	137
rect	528	137	529	138
rect	528	138	529	139
rect	528	139	529	140
rect	528	140	529	141
rect	528	141	529	142
rect	528	142	529	143
rect	528	143	529	144
rect	528	144	529	145
rect	528	145	529	146
rect	528	146	529	147
rect	528	147	529	148
rect	528	148	529	149
rect	528	149	529	150
rect	528	150	529	151
rect	528	151	529	152
rect	528	152	529	153
rect	528	153	529	154
rect	528	154	529	155
rect	528	155	529	156
rect	528	156	529	157
rect	528	157	529	158
rect	528	158	529	159
rect	528	159	529	160
rect	528	160	529	161
rect	528	161	529	162
rect	528	162	529	163
rect	528	163	529	164
rect	528	164	529	165
rect	528	165	529	166
rect	528	166	529	167
rect	528	167	529	168
rect	528	168	529	169
rect	528	169	529	170
rect	528	170	529	171
rect	528	171	529	172
rect	528	172	529	173
rect	528	173	529	174
rect	528	174	529	175
rect	528	175	529	176
rect	528	176	529	177
rect	528	177	529	178
rect	528	178	529	179
rect	528	179	529	180
rect	528	180	529	181
rect	528	181	529	182
rect	528	182	529	183
rect	528	183	529	184
rect	528	184	529	185
rect	528	185	529	186
rect	528	186	529	187
rect	528	187	529	188
rect	528	188	529	189
rect	528	189	529	190
rect	528	190	529	191
rect	528	191	529	192
rect	528	192	529	193
rect	528	193	529	194
rect	528	194	529	195
rect	528	195	529	196
rect	528	196	529	197
rect	528	197	529	198
rect	528	198	529	199
rect	528	199	529	200
rect	528	200	529	201
rect	528	201	529	202
rect	528	202	529	203
rect	528	203	529	204
rect	528	204	529	205
rect	528	205	529	206
rect	528	206	529	207
rect	528	207	529	208
rect	528	208	529	209
rect	528	209	529	210
rect	528	210	529	211
rect	528	211	529	212
rect	528	212	529	213
rect	528	213	529	214
rect	528	214	529	215
rect	528	215	529	216
rect	528	216	529	217
rect	528	217	529	218
rect	528	218	529	219
rect	528	219	529	220
rect	528	220	529	221
rect	528	221	529	222
rect	528	222	529	223
rect	528	223	529	224
rect	528	224	529	225
rect	528	225	529	226
rect	528	226	529	227
rect	528	227	529	228
rect	528	228	529	229
rect	528	229	529	230
rect	528	230	529	231
rect	528	231	529	232
rect	528	232	529	233
rect	528	233	529	234
rect	528	234	529	235
rect	528	235	529	236
rect	528	236	529	237
rect	528	237	529	238
rect	528	238	529	239
rect	528	239	529	240
rect	528	240	529	241
rect	528	241	529	242
rect	528	242	529	243
rect	528	243	529	244
rect	528	244	529	245
rect	528	245	529	246
rect	528	246	529	247
rect	528	247	529	248
rect	528	248	529	249
rect	528	249	529	250
rect	528	250	529	251
rect	528	251	529	252
rect	528	252	529	253
rect	528	253	529	254
rect	528	254	529	255
rect	528	255	529	256
rect	528	256	529	257
rect	528	257	529	258
rect	528	258	529	259
rect	528	259	529	260
rect	528	260	529	261
rect	528	261	529	262
rect	528	262	529	263
rect	528	263	529	264
rect	528	264	529	265
rect	528	265	529	266
rect	528	266	529	267
rect	528	267	529	268
rect	528	268	529	269
rect	528	269	529	270
rect	528	270	529	271
rect	528	271	529	272
rect	528	272	529	273
rect	528	273	529	274
rect	528	274	529	275
rect	528	275	529	276
rect	528	276	529	277
rect	528	277	529	278
rect	528	278	529	279
rect	528	279	529	280
rect	528	280	529	281
rect	528	281	529	282
rect	528	282	529	283
rect	528	283	529	284
rect	528	284	529	285
rect	528	285	529	286
rect	528	286	529	287
rect	528	287	529	288
rect	529	0	530	1
rect	529	1	530	2
rect	529	2	530	3
rect	529	3	530	4
rect	529	4	530	5
rect	529	5	530	6
rect	529	6	530	7
rect	529	7	530	8
rect	529	8	530	9
rect	529	9	530	10
rect	529	10	530	11
rect	529	11	530	12
rect	529	12	530	13
rect	529	13	530	14
rect	529	14	530	15
rect	529	15	530	16
rect	529	16	530	17
rect	529	17	530	18
rect	529	18	530	19
rect	529	19	530	20
rect	529	20	530	21
rect	529	21	530	22
rect	529	22	530	23
rect	529	23	530	24
rect	529	24	530	25
rect	529	25	530	26
rect	529	26	530	27
rect	529	27	530	28
rect	529	28	530	29
rect	529	29	530	30
rect	529	30	530	31
rect	529	31	530	32
rect	529	32	530	33
rect	529	33	530	34
rect	529	34	530	35
rect	529	35	530	36
rect	529	36	530	37
rect	529	37	530	38
rect	529	38	530	39
rect	529	39	530	40
rect	529	40	530	41
rect	529	41	530	42
rect	529	42	530	43
rect	529	43	530	44
rect	529	44	530	45
rect	529	45	530	46
rect	529	46	530	47
rect	529	47	530	48
rect	529	48	530	49
rect	529	49	530	50
rect	529	50	530	51
rect	529	51	530	52
rect	529	52	530	53
rect	529	53	530	54
rect	529	54	530	55
rect	529	55	530	56
rect	529	56	530	57
rect	529	57	530	58
rect	529	58	530	59
rect	529	59	530	60
rect	529	60	530	61
rect	529	61	530	62
rect	529	62	530	63
rect	529	63	530	64
rect	529	64	530	65
rect	529	65	530	66
rect	529	66	530	67
rect	529	67	530	68
rect	529	68	530	69
rect	529	69	530	70
rect	529	70	530	71
rect	529	71	530	72
rect	529	72	530	73
rect	529	73	530	74
rect	529	74	530	75
rect	529	75	530	76
rect	529	76	530	77
rect	529	77	530	78
rect	529	78	530	79
rect	529	79	530	80
rect	529	80	530	81
rect	529	81	530	82
rect	529	82	530	83
rect	529	83	530	84
rect	529	84	530	85
rect	529	85	530	86
rect	529	86	530	87
rect	529	87	530	88
rect	529	88	530	89
rect	529	89	530	90
rect	529	90	530	91
rect	529	91	530	92
rect	529	92	530	93
rect	529	93	530	94
rect	529	94	530	95
rect	529	95	530	96
rect	529	96	530	97
rect	529	97	530	98
rect	529	98	530	99
rect	529	99	530	100
rect	529	100	530	101
rect	529	101	530	102
rect	529	102	530	103
rect	529	103	530	104
rect	529	104	530	105
rect	529	105	530	106
rect	529	106	530	107
rect	529	107	530	108
rect	529	108	530	109
rect	529	109	530	110
rect	529	110	530	111
rect	529	111	530	112
rect	529	112	530	113
rect	529	113	530	114
rect	529	114	530	115
rect	529	115	530	116
rect	529	116	530	117
rect	529	117	530	118
rect	529	118	530	119
rect	529	119	530	120
rect	529	120	530	121
rect	529	121	530	122
rect	529	122	530	123
rect	529	123	530	124
rect	529	124	530	125
rect	529	125	530	126
rect	529	126	530	127
rect	529	127	530	128
rect	529	128	530	129
rect	529	129	530	130
rect	529	130	530	131
rect	529	131	530	132
rect	529	132	530	133
rect	529	133	530	134
rect	529	134	530	135
rect	529	135	530	136
rect	529	136	530	137
rect	529	137	530	138
rect	529	138	530	139
rect	529	139	530	140
rect	529	140	530	141
rect	529	141	530	142
rect	529	142	530	143
rect	529	143	530	144
rect	529	144	530	145
rect	529	145	530	146
rect	529	146	530	147
rect	529	147	530	148
rect	529	148	530	149
rect	529	149	530	150
rect	529	150	530	151
rect	529	151	530	152
rect	529	152	530	153
rect	529	153	530	154
rect	529	154	530	155
rect	529	155	530	156
rect	529	156	530	157
rect	529	157	530	158
rect	529	158	530	159
rect	529	159	530	160
rect	529	160	530	161
rect	529	161	530	162
rect	529	162	530	163
rect	529	163	530	164
rect	529	164	530	165
rect	529	165	530	166
rect	529	166	530	167
rect	529	167	530	168
rect	529	168	530	169
rect	529	169	530	170
rect	529	170	530	171
rect	529	171	530	172
rect	529	172	530	173
rect	529	173	530	174
rect	529	174	530	175
rect	529	175	530	176
rect	529	176	530	177
rect	529	177	530	178
rect	529	178	530	179
rect	529	179	530	180
rect	529	180	530	181
rect	529	181	530	182
rect	529	182	530	183
rect	529	183	530	184
rect	529	184	530	185
rect	529	185	530	186
rect	529	186	530	187
rect	529	187	530	188
rect	529	188	530	189
rect	529	189	530	190
rect	529	190	530	191
rect	529	191	530	192
rect	529	192	530	193
rect	529	193	530	194
rect	529	194	530	195
rect	529	195	530	196
rect	529	196	530	197
rect	529	197	530	198
rect	529	198	530	199
rect	529	199	530	200
rect	529	200	530	201
rect	529	201	530	202
rect	529	202	530	203
rect	529	203	530	204
rect	529	204	530	205
rect	529	205	530	206
rect	529	206	530	207
rect	529	207	530	208
rect	529	208	530	209
rect	529	209	530	210
rect	529	210	530	211
rect	529	211	530	212
rect	529	212	530	213
rect	529	213	530	214
rect	529	214	530	215
rect	529	215	530	216
rect	529	216	530	217
rect	529	217	530	218
rect	529	218	530	219
rect	529	219	530	220
rect	529	220	530	221
rect	529	221	530	222
rect	529	222	530	223
rect	529	223	530	224
rect	529	224	530	225
rect	529	225	530	226
rect	529	226	530	227
rect	529	227	530	228
rect	529	228	530	229
rect	529	229	530	230
rect	529	230	530	231
rect	529	231	530	232
rect	529	232	530	233
rect	529	233	530	234
rect	529	234	530	235
rect	529	235	530	236
rect	529	236	530	237
rect	529	237	530	238
rect	529	238	530	239
rect	529	239	530	240
rect	529	240	530	241
rect	529	241	530	242
rect	529	242	530	243
rect	529	243	530	244
rect	529	244	530	245
rect	529	245	530	246
rect	529	246	530	247
rect	529	247	530	248
rect	529	248	530	249
rect	529	249	530	250
rect	529	250	530	251
rect	529	251	530	252
rect	529	252	530	253
rect	529	253	530	254
rect	529	254	530	255
rect	529	255	530	256
rect	529	256	530	257
rect	529	257	530	258
rect	529	258	530	259
rect	529	259	530	260
rect	529	260	530	261
rect	529	261	530	262
rect	529	262	530	263
rect	529	263	530	264
rect	529	264	530	265
rect	529	265	530	266
rect	529	266	530	267
rect	529	267	530	268
rect	529	268	530	269
rect	529	269	530	270
rect	529	270	530	271
rect	529	271	530	272
rect	529	272	530	273
rect	529	273	530	274
rect	529	274	530	275
rect	529	275	530	276
rect	529	276	530	277
rect	529	277	530	278
rect	529	278	530	279
rect	529	279	530	280
rect	529	280	530	281
rect	529	281	530	282
rect	529	282	530	283
rect	529	283	530	284
rect	529	284	530	285
rect	529	285	530	286
rect	529	286	530	287
rect	529	287	530	288
rect	547	0	548	1
rect	547	1	548	2
rect	547	2	548	3
rect	547	3	548	4
rect	547	4	548	5
rect	547	5	548	6
rect	547	6	548	7
rect	547	7	548	8
rect	547	8	548	9
rect	547	9	548	10
rect	547	10	548	11
rect	547	11	548	12
rect	547	12	548	13
rect	547	13	548	14
rect	547	14	548	15
rect	547	15	548	16
rect	547	16	548	17
rect	547	17	548	18
rect	547	18	548	19
rect	547	19	548	20
rect	547	20	548	21
rect	547	21	548	22
rect	547	22	548	23
rect	547	23	548	24
rect	547	24	548	25
rect	547	25	548	26
rect	547	26	548	27
rect	547	27	548	28
rect	547	28	548	29
rect	547	29	548	30
rect	547	30	548	31
rect	547	31	548	32
rect	547	32	548	33
rect	547	33	548	34
rect	547	34	548	35
rect	547	35	548	36
rect	547	36	548	37
rect	547	37	548	38
rect	547	38	548	39
rect	547	39	548	40
rect	547	40	548	41
rect	547	41	548	42
rect	547	42	548	43
rect	547	43	548	44
rect	547	44	548	45
rect	547	45	548	46
rect	547	46	548	47
rect	547	47	548	48
rect	547	48	548	49
rect	547	49	548	50
rect	547	50	548	51
rect	547	51	548	52
rect	547	52	548	53
rect	547	53	548	54
rect	547	54	548	55
rect	547	55	548	56
rect	547	56	548	57
rect	547	57	548	58
rect	547	58	548	59
rect	547	59	548	60
rect	547	60	548	61
rect	547	61	548	62
rect	547	62	548	63
rect	547	63	548	64
rect	547	64	548	65
rect	547	65	548	66
rect	547	66	548	67
rect	547	67	548	68
rect	547	68	548	69
rect	547	69	548	70
rect	547	70	548	71
rect	547	71	548	72
rect	547	72	548	73
rect	547	73	548	74
rect	547	74	548	75
rect	547	75	548	76
rect	547	76	548	77
rect	547	77	548	78
rect	547	78	548	79
rect	547	79	548	80
rect	547	80	548	81
rect	547	81	548	82
rect	547	82	548	83
rect	547	83	548	84
rect	547	84	548	85
rect	547	85	548	86
rect	547	86	548	87
rect	547	87	548	88
rect	547	88	548	89
rect	547	89	548	90
rect	547	90	548	91
rect	547	91	548	92
rect	547	92	548	93
rect	547	93	548	94
rect	547	94	548	95
rect	547	95	548	96
rect	547	96	548	97
rect	547	97	548	98
rect	547	98	548	99
rect	547	99	548	100
rect	547	100	548	101
rect	547	101	548	102
rect	547	102	548	103
rect	547	103	548	104
rect	547	104	548	105
rect	547	105	548	106
rect	547	106	548	107
rect	547	107	548	108
rect	547	108	548	109
rect	547	109	548	110
rect	547	110	548	111
rect	547	111	548	112
rect	547	112	548	113
rect	547	113	548	114
rect	547	114	548	115
rect	547	115	548	116
rect	547	116	548	117
rect	547	117	548	118
rect	547	118	548	119
rect	547	119	548	120
rect	547	120	548	121
rect	547	121	548	122
rect	547	122	548	123
rect	547	123	548	124
rect	547	124	548	125
rect	547	125	548	126
rect	547	126	548	127
rect	547	127	548	128
rect	547	128	548	129
rect	547	129	548	130
rect	547	130	548	131
rect	547	131	548	132
rect	547	132	548	133
rect	547	133	548	134
rect	547	134	548	135
rect	547	135	548	136
rect	547	136	548	137
rect	547	137	548	138
rect	547	138	548	139
rect	547	139	548	140
rect	547	140	548	141
rect	547	141	548	142
rect	547	142	548	143
rect	547	143	548	144
rect	547	144	548	145
rect	547	145	548	146
rect	547	146	548	147
rect	547	147	548	148
rect	547	148	548	149
rect	547	149	548	150
rect	547	150	548	151
rect	547	151	548	152
rect	547	152	548	153
rect	547	153	548	154
rect	547	154	548	155
rect	547	155	548	156
rect	547	156	548	157
rect	547	157	548	158
rect	547	158	548	159
rect	547	159	548	160
rect	547	160	548	161
rect	547	161	548	162
rect	547	162	548	163
rect	547	163	548	164
rect	547	164	548	165
rect	547	165	548	166
rect	547	166	548	167
rect	547	167	548	168
rect	547	168	548	169
rect	547	169	548	170
rect	547	170	548	171
rect	547	171	548	172
rect	547	172	548	173
rect	547	173	548	174
rect	547	174	548	175
rect	547	175	548	176
rect	547	176	548	177
rect	547	177	548	178
rect	547	178	548	179
rect	547	179	548	180
rect	547	180	548	181
rect	547	181	548	182
rect	547	182	548	183
rect	547	183	548	184
rect	547	184	548	185
rect	547	185	548	186
rect	547	186	548	187
rect	547	187	548	188
rect	547	188	548	189
rect	547	189	548	190
rect	547	190	548	191
rect	547	191	548	192
rect	547	192	548	193
rect	547	193	548	194
rect	547	194	548	195
rect	547	195	548	196
rect	547	196	548	197
rect	547	197	548	198
rect	547	198	548	199
rect	547	199	548	200
rect	547	200	548	201
rect	547	201	548	202
rect	547	202	548	203
rect	547	203	548	204
rect	547	204	548	205
rect	547	205	548	206
rect	547	206	548	207
rect	547	207	548	208
rect	547	208	548	209
rect	547	209	548	210
rect	547	210	548	211
rect	547	211	548	212
rect	547	212	548	213
rect	547	213	548	214
rect	547	214	548	215
rect	547	215	548	216
rect	547	216	548	217
rect	547	217	548	218
rect	547	218	548	219
rect	547	219	548	220
rect	547	220	548	221
rect	547	221	548	222
rect	547	222	548	223
rect	547	223	548	224
rect	547	224	548	225
rect	547	225	548	226
rect	547	226	548	227
rect	547	227	548	228
rect	547	228	548	229
rect	547	229	548	230
rect	547	230	548	231
rect	547	231	548	232
rect	547	232	548	233
rect	547	233	548	234
rect	547	234	548	235
rect	547	235	548	236
rect	547	236	548	237
rect	547	237	548	238
rect	547	238	548	239
rect	547	239	548	240
rect	547	240	548	241
rect	547	241	548	242
rect	547	242	548	243
rect	547	243	548	244
rect	547	244	548	245
rect	547	245	548	246
rect	547	246	548	247
rect	547	247	548	248
rect	547	248	548	249
rect	547	249	548	250
rect	547	250	548	251
rect	547	251	548	252
rect	547	252	548	253
rect	547	253	548	254
rect	547	254	548	255
rect	547	255	548	256
rect	547	256	548	257
rect	547	257	548	258
rect	547	258	548	259
rect	547	259	548	260
rect	547	260	548	261
rect	547	261	548	262
rect	547	262	548	263
rect	547	263	548	264
rect	547	264	548	265
rect	547	265	548	266
rect	547	266	548	267
rect	547	267	548	268
rect	547	268	548	269
rect	547	269	548	270
rect	547	270	548	271
rect	547	271	548	272
rect	547	272	548	273
rect	547	273	548	274
rect	547	274	548	275
rect	547	275	548	276
rect	547	276	548	277
rect	547	277	548	278
rect	547	278	548	279
rect	547	279	548	280
rect	547	280	548	281
rect	547	281	548	282
rect	547	282	548	283
rect	547	283	548	284
rect	547	284	548	285
rect	548	0	549	1
rect	548	1	549	2
rect	548	2	549	3
rect	548	3	549	4
rect	548	4	549	5
rect	548	5	549	6
rect	548	6	549	7
rect	548	7	549	8
rect	548	8	549	9
rect	548	9	549	10
rect	548	10	549	11
rect	548	11	549	12
rect	548	12	549	13
rect	548	13	549	14
rect	548	14	549	15
rect	548	15	549	16
rect	548	16	549	17
rect	548	17	549	18
rect	548	18	549	19
rect	548	19	549	20
rect	548	20	549	21
rect	548	21	549	22
rect	548	22	549	23
rect	548	23	549	24
rect	548	24	549	25
rect	548	25	549	26
rect	548	26	549	27
rect	548	27	549	28
rect	548	28	549	29
rect	548	29	549	30
rect	548	30	549	31
rect	548	31	549	32
rect	548	32	549	33
rect	548	33	549	34
rect	548	34	549	35
rect	548	35	549	36
rect	548	36	549	37
rect	548	37	549	38
rect	548	38	549	39
rect	548	39	549	40
rect	548	40	549	41
rect	548	41	549	42
rect	548	42	549	43
rect	548	43	549	44
rect	548	44	549	45
rect	548	45	549	46
rect	548	46	549	47
rect	548	47	549	48
rect	548	48	549	49
rect	548	49	549	50
rect	548	50	549	51
rect	548	51	549	52
rect	548	52	549	53
rect	548	53	549	54
rect	548	54	549	55
rect	548	55	549	56
rect	548	56	549	57
rect	548	57	549	58
rect	548	58	549	59
rect	548	59	549	60
rect	548	60	549	61
rect	548	61	549	62
rect	548	62	549	63
rect	548	63	549	64
rect	548	64	549	65
rect	548	65	549	66
rect	548	66	549	67
rect	548	67	549	68
rect	548	68	549	69
rect	548	69	549	70
rect	548	70	549	71
rect	548	71	549	72
rect	548	72	549	73
rect	548	73	549	74
rect	548	74	549	75
rect	548	75	549	76
rect	548	76	549	77
rect	548	77	549	78
rect	548	78	549	79
rect	548	79	549	80
rect	548	80	549	81
rect	548	81	549	82
rect	548	82	549	83
rect	548	83	549	84
rect	548	84	549	85
rect	548	85	549	86
rect	548	86	549	87
rect	548	87	549	88
rect	548	88	549	89
rect	548	89	549	90
rect	548	90	549	91
rect	548	91	549	92
rect	548	92	549	93
rect	548	93	549	94
rect	548	94	549	95
rect	548	95	549	96
rect	548	96	549	97
rect	548	97	549	98
rect	548	98	549	99
rect	548	99	549	100
rect	548	100	549	101
rect	548	101	549	102
rect	548	102	549	103
rect	548	103	549	104
rect	548	104	549	105
rect	548	105	549	106
rect	548	106	549	107
rect	548	107	549	108
rect	548	108	549	109
rect	548	109	549	110
rect	548	110	549	111
rect	548	111	549	112
rect	548	112	549	113
rect	548	113	549	114
rect	548	114	549	115
rect	548	115	549	116
rect	548	116	549	117
rect	548	117	549	118
rect	548	118	549	119
rect	548	119	549	120
rect	548	120	549	121
rect	548	121	549	122
rect	548	122	549	123
rect	548	123	549	124
rect	548	124	549	125
rect	548	125	549	126
rect	548	126	549	127
rect	548	127	549	128
rect	548	128	549	129
rect	548	129	549	130
rect	548	130	549	131
rect	548	131	549	132
rect	548	132	549	133
rect	548	133	549	134
rect	548	134	549	135
rect	548	135	549	136
rect	548	136	549	137
rect	548	137	549	138
rect	548	138	549	139
rect	548	139	549	140
rect	548	140	549	141
rect	548	141	549	142
rect	548	142	549	143
rect	548	143	549	144
rect	548	144	549	145
rect	548	145	549	146
rect	548	146	549	147
rect	548	147	549	148
rect	548	148	549	149
rect	548	149	549	150
rect	548	150	549	151
rect	548	151	549	152
rect	548	152	549	153
rect	548	153	549	154
rect	548	154	549	155
rect	548	155	549	156
rect	548	156	549	157
rect	548	157	549	158
rect	548	158	549	159
rect	548	159	549	160
rect	548	160	549	161
rect	548	161	549	162
rect	548	162	549	163
rect	548	163	549	164
rect	548	164	549	165
rect	548	165	549	166
rect	548	166	549	167
rect	548	167	549	168
rect	548	168	549	169
rect	548	169	549	170
rect	548	170	549	171
rect	548	171	549	172
rect	548	172	549	173
rect	548	173	549	174
rect	548	174	549	175
rect	548	175	549	176
rect	548	176	549	177
rect	548	177	549	178
rect	548	178	549	179
rect	548	179	549	180
rect	548	180	549	181
rect	548	181	549	182
rect	548	182	549	183
rect	548	183	549	184
rect	548	184	549	185
rect	548	185	549	186
rect	548	186	549	187
rect	548	187	549	188
rect	548	188	549	189
rect	548	189	549	190
rect	548	190	549	191
rect	548	191	549	192
rect	548	192	549	193
rect	548	193	549	194
rect	548	194	549	195
rect	548	195	549	196
rect	548	196	549	197
rect	548	197	549	198
rect	548	198	549	199
rect	548	199	549	200
rect	548	200	549	201
rect	548	201	549	202
rect	548	202	549	203
rect	548	203	549	204
rect	548	204	549	205
rect	548	205	549	206
rect	548	206	549	207
rect	548	207	549	208
rect	548	208	549	209
rect	548	209	549	210
rect	548	210	549	211
rect	548	211	549	212
rect	548	212	549	213
rect	548	213	549	214
rect	548	214	549	215
rect	548	215	549	216
rect	548	216	549	217
rect	548	217	549	218
rect	548	218	549	219
rect	548	219	549	220
rect	548	220	549	221
rect	548	221	549	222
rect	548	222	549	223
rect	548	223	549	224
rect	548	224	549	225
rect	548	225	549	226
rect	548	226	549	227
rect	548	227	549	228
rect	548	228	549	229
rect	548	229	549	230
rect	548	230	549	231
rect	548	231	549	232
rect	548	232	549	233
rect	548	233	549	234
rect	548	234	549	235
rect	548	235	549	236
rect	548	236	549	237
rect	548	237	549	238
rect	548	238	549	239
rect	548	239	549	240
rect	548	240	549	241
rect	548	241	549	242
rect	548	242	549	243
rect	548	243	549	244
rect	548	244	549	245
rect	548	245	549	246
rect	548	246	549	247
rect	548	247	549	248
rect	548	248	549	249
rect	548	249	549	250
rect	548	250	549	251
rect	548	251	549	252
rect	548	252	549	253
rect	548	253	549	254
rect	548	254	549	255
rect	548	255	549	256
rect	548	256	549	257
rect	548	257	549	258
rect	548	258	549	259
rect	548	259	549	260
rect	548	260	549	261
rect	548	261	549	262
rect	548	262	549	263
rect	548	263	549	264
rect	548	264	549	265
rect	548	265	549	266
rect	548	266	549	267
rect	548	267	549	268
rect	548	268	549	269
rect	548	269	549	270
rect	548	270	549	271
rect	548	271	549	272
rect	548	272	549	273
rect	548	273	549	274
rect	548	274	549	275
rect	548	275	549	276
rect	548	276	549	277
rect	548	277	549	278
rect	548	278	549	279
rect	548	279	549	280
rect	548	280	549	281
rect	548	281	549	282
rect	548	282	549	283
rect	548	283	549	284
rect	548	284	549	285
rect	549	0	550	1
rect	549	1	550	2
rect	549	2	550	3
rect	549	3	550	4
rect	549	4	550	5
rect	549	5	550	6
rect	549	6	550	7
rect	549	7	550	8
rect	549	8	550	9
rect	549	9	550	10
rect	549	10	550	11
rect	549	11	550	12
rect	549	12	550	13
rect	549	13	550	14
rect	549	14	550	15
rect	549	15	550	16
rect	549	16	550	17
rect	549	17	550	18
rect	549	18	550	19
rect	549	19	550	20
rect	549	20	550	21
rect	549	21	550	22
rect	549	22	550	23
rect	549	23	550	24
rect	549	24	550	25
rect	549	25	550	26
rect	549	26	550	27
rect	549	27	550	28
rect	549	28	550	29
rect	549	29	550	30
rect	549	30	550	31
rect	549	31	550	32
rect	549	32	550	33
rect	549	33	550	34
rect	549	34	550	35
rect	549	35	550	36
rect	549	36	550	37
rect	549	37	550	38
rect	549	38	550	39
rect	549	39	550	40
rect	549	40	550	41
rect	549	41	550	42
rect	549	42	550	43
rect	549	43	550	44
rect	549	44	550	45
rect	549	45	550	46
rect	549	46	550	47
rect	549	47	550	48
rect	549	48	550	49
rect	549	49	550	50
rect	549	50	550	51
rect	549	51	550	52
rect	549	52	550	53
rect	549	53	550	54
rect	549	54	550	55
rect	549	55	550	56
rect	549	56	550	57
rect	549	57	550	58
rect	549	58	550	59
rect	549	59	550	60
rect	549	60	550	61
rect	549	61	550	62
rect	549	62	550	63
rect	549	63	550	64
rect	549	64	550	65
rect	549	65	550	66
rect	549	66	550	67
rect	549	67	550	68
rect	549	68	550	69
rect	549	69	550	70
rect	549	70	550	71
rect	549	71	550	72
rect	549	72	550	73
rect	549	73	550	74
rect	549	74	550	75
rect	549	75	550	76
rect	549	76	550	77
rect	549	77	550	78
rect	549	78	550	79
rect	549	79	550	80
rect	549	80	550	81
rect	549	81	550	82
rect	549	82	550	83
rect	549	83	550	84
rect	549	84	550	85
rect	549	85	550	86
rect	549	86	550	87
rect	549	87	550	88
rect	549	88	550	89
rect	549	89	550	90
rect	549	90	550	91
rect	549	91	550	92
rect	549	92	550	93
rect	549	93	550	94
rect	549	94	550	95
rect	549	95	550	96
rect	549	96	550	97
rect	549	97	550	98
rect	549	98	550	99
rect	549	99	550	100
rect	549	100	550	101
rect	549	101	550	102
rect	549	102	550	103
rect	549	103	550	104
rect	549	104	550	105
rect	549	105	550	106
rect	549	106	550	107
rect	549	107	550	108
rect	549	108	550	109
rect	549	109	550	110
rect	549	110	550	111
rect	549	111	550	112
rect	549	112	550	113
rect	549	113	550	114
rect	549	114	550	115
rect	549	115	550	116
rect	549	116	550	117
rect	549	117	550	118
rect	549	118	550	119
rect	549	119	550	120
rect	549	120	550	121
rect	549	121	550	122
rect	549	122	550	123
rect	549	123	550	124
rect	549	124	550	125
rect	549	125	550	126
rect	549	126	550	127
rect	549	127	550	128
rect	549	128	550	129
rect	549	129	550	130
rect	549	130	550	131
rect	549	131	550	132
rect	549	132	550	133
rect	549	133	550	134
rect	549	134	550	135
rect	549	135	550	136
rect	549	136	550	137
rect	549	137	550	138
rect	549	138	550	139
rect	549	139	550	140
rect	549	140	550	141
rect	549	141	550	142
rect	549	142	550	143
rect	549	143	550	144
rect	549	144	550	145
rect	549	145	550	146
rect	549	146	550	147
rect	549	147	550	148
rect	549	148	550	149
rect	549	149	550	150
rect	549	150	550	151
rect	549	151	550	152
rect	549	152	550	153
rect	549	153	550	154
rect	549	154	550	155
rect	549	155	550	156
rect	549	156	550	157
rect	549	157	550	158
rect	549	158	550	159
rect	549	159	550	160
rect	549	160	550	161
rect	549	161	550	162
rect	549	162	550	163
rect	549	163	550	164
rect	549	164	550	165
rect	549	165	550	166
rect	549	166	550	167
rect	549	167	550	168
rect	549	168	550	169
rect	549	169	550	170
rect	549	170	550	171
rect	549	171	550	172
rect	549	172	550	173
rect	549	173	550	174
rect	549	174	550	175
rect	549	175	550	176
rect	549	176	550	177
rect	549	177	550	178
rect	549	178	550	179
rect	549	179	550	180
rect	549	180	550	181
rect	549	181	550	182
rect	549	182	550	183
rect	549	183	550	184
rect	549	184	550	185
rect	549	185	550	186
rect	549	186	550	187
rect	549	187	550	188
rect	549	188	550	189
rect	549	189	550	190
rect	549	190	550	191
rect	549	191	550	192
rect	549	192	550	193
rect	549	193	550	194
rect	549	194	550	195
rect	549	195	550	196
rect	549	196	550	197
rect	549	197	550	198
rect	549	198	550	199
rect	549	199	550	200
rect	549	200	550	201
rect	549	201	550	202
rect	549	202	550	203
rect	549	203	550	204
rect	549	204	550	205
rect	549	205	550	206
rect	549	206	550	207
rect	549	207	550	208
rect	549	208	550	209
rect	549	209	550	210
rect	549	210	550	211
rect	549	211	550	212
rect	549	212	550	213
rect	549	213	550	214
rect	549	214	550	215
rect	549	215	550	216
rect	549	216	550	217
rect	549	217	550	218
rect	549	218	550	219
rect	549	219	550	220
rect	549	220	550	221
rect	549	221	550	222
rect	549	222	550	223
rect	549	223	550	224
rect	549	224	550	225
rect	549	225	550	226
rect	549	226	550	227
rect	549	227	550	228
rect	549	228	550	229
rect	549	229	550	230
rect	549	230	550	231
rect	549	231	550	232
rect	549	232	550	233
rect	549	233	550	234
rect	549	234	550	235
rect	549	235	550	236
rect	549	236	550	237
rect	549	237	550	238
rect	549	238	550	239
rect	549	239	550	240
rect	549	240	550	241
rect	549	241	550	242
rect	549	242	550	243
rect	549	243	550	244
rect	549	244	550	245
rect	549	245	550	246
rect	549	246	550	247
rect	549	247	550	248
rect	549	248	550	249
rect	549	249	550	250
rect	549	250	550	251
rect	549	251	550	252
rect	549	252	550	253
rect	549	253	550	254
rect	549	254	550	255
rect	549	255	550	256
rect	549	256	550	257
rect	549	257	550	258
rect	549	258	550	259
rect	549	259	550	260
rect	549	260	550	261
rect	549	261	550	262
rect	549	262	550	263
rect	549	263	550	264
rect	549	264	550	265
rect	549	265	550	266
rect	549	266	550	267
rect	549	267	550	268
rect	549	268	550	269
rect	549	269	550	270
rect	549	270	550	271
rect	549	271	550	272
rect	549	272	550	273
rect	549	273	550	274
rect	549	274	550	275
rect	549	275	550	276
rect	549	276	550	277
rect	549	277	550	278
rect	549	278	550	279
rect	549	279	550	280
rect	549	280	550	281
rect	549	281	550	282
rect	549	282	550	283
rect	549	283	550	284
rect	549	284	550	285
rect	550	0	551	1
rect	550	1	551	2
rect	550	2	551	3
rect	550	3	551	4
rect	550	4	551	5
rect	550	5	551	6
rect	550	6	551	7
rect	550	7	551	8
rect	550	8	551	9
rect	550	9	551	10
rect	550	10	551	11
rect	550	11	551	12
rect	550	12	551	13
rect	550	13	551	14
rect	550	14	551	15
rect	550	15	551	16
rect	550	16	551	17
rect	550	17	551	18
rect	550	18	551	19
rect	550	19	551	20
rect	550	20	551	21
rect	550	21	551	22
rect	550	22	551	23
rect	550	23	551	24
rect	550	24	551	25
rect	550	25	551	26
rect	550	26	551	27
rect	550	27	551	28
rect	550	28	551	29
rect	550	29	551	30
rect	550	30	551	31
rect	550	31	551	32
rect	550	32	551	33
rect	550	33	551	34
rect	550	34	551	35
rect	550	35	551	36
rect	550	36	551	37
rect	550	37	551	38
rect	550	38	551	39
rect	550	39	551	40
rect	550	40	551	41
rect	550	41	551	42
rect	550	42	551	43
rect	550	43	551	44
rect	550	44	551	45
rect	550	45	551	46
rect	550	46	551	47
rect	550	47	551	48
rect	550	48	551	49
rect	550	49	551	50
rect	550	50	551	51
rect	550	51	551	52
rect	550	52	551	53
rect	550	53	551	54
rect	550	54	551	55
rect	550	55	551	56
rect	550	56	551	57
rect	550	57	551	58
rect	550	58	551	59
rect	550	59	551	60
rect	550	60	551	61
rect	550	61	551	62
rect	550	62	551	63
rect	550	63	551	64
rect	550	64	551	65
rect	550	65	551	66
rect	550	66	551	67
rect	550	67	551	68
rect	550	68	551	69
rect	550	69	551	70
rect	550	70	551	71
rect	550	71	551	72
rect	550	72	551	73
rect	550	73	551	74
rect	550	74	551	75
rect	550	75	551	76
rect	550	76	551	77
rect	550	77	551	78
rect	550	78	551	79
rect	550	79	551	80
rect	550	80	551	81
rect	550	81	551	82
rect	550	82	551	83
rect	550	83	551	84
rect	550	84	551	85
rect	550	85	551	86
rect	550	86	551	87
rect	550	87	551	88
rect	550	88	551	89
rect	550	89	551	90
rect	550	90	551	91
rect	550	91	551	92
rect	550	92	551	93
rect	550	93	551	94
rect	550	94	551	95
rect	550	95	551	96
rect	550	96	551	97
rect	550	97	551	98
rect	550	98	551	99
rect	550	99	551	100
rect	550	100	551	101
rect	550	101	551	102
rect	550	102	551	103
rect	550	103	551	104
rect	550	104	551	105
rect	550	105	551	106
rect	550	106	551	107
rect	550	107	551	108
rect	550	108	551	109
rect	550	109	551	110
rect	550	110	551	111
rect	550	111	551	112
rect	550	112	551	113
rect	550	113	551	114
rect	550	114	551	115
rect	550	115	551	116
rect	550	116	551	117
rect	550	117	551	118
rect	550	118	551	119
rect	550	119	551	120
rect	550	120	551	121
rect	550	121	551	122
rect	550	122	551	123
rect	550	123	551	124
rect	550	124	551	125
rect	550	125	551	126
rect	550	126	551	127
rect	550	127	551	128
rect	550	128	551	129
rect	550	129	551	130
rect	550	130	551	131
rect	550	131	551	132
rect	550	132	551	133
rect	550	133	551	134
rect	550	134	551	135
rect	550	135	551	136
rect	550	136	551	137
rect	550	137	551	138
rect	550	138	551	139
rect	550	139	551	140
rect	550	140	551	141
rect	550	141	551	142
rect	550	142	551	143
rect	550	143	551	144
rect	550	144	551	145
rect	550	145	551	146
rect	550	146	551	147
rect	550	147	551	148
rect	550	148	551	149
rect	550	149	551	150
rect	550	150	551	151
rect	550	151	551	152
rect	550	152	551	153
rect	550	153	551	154
rect	550	154	551	155
rect	550	155	551	156
rect	550	156	551	157
rect	550	157	551	158
rect	550	158	551	159
rect	550	159	551	160
rect	550	160	551	161
rect	550	161	551	162
rect	550	162	551	163
rect	550	163	551	164
rect	550	164	551	165
rect	550	165	551	166
rect	550	166	551	167
rect	550	167	551	168
rect	550	168	551	169
rect	550	169	551	170
rect	550	170	551	171
rect	550	171	551	172
rect	550	172	551	173
rect	550	173	551	174
rect	550	174	551	175
rect	550	175	551	176
rect	550	176	551	177
rect	550	177	551	178
rect	550	178	551	179
rect	550	179	551	180
rect	550	180	551	181
rect	550	181	551	182
rect	550	182	551	183
rect	550	183	551	184
rect	550	184	551	185
rect	550	185	551	186
rect	550	186	551	187
rect	550	187	551	188
rect	550	188	551	189
rect	550	189	551	190
rect	550	190	551	191
rect	550	191	551	192
rect	550	192	551	193
rect	550	193	551	194
rect	550	194	551	195
rect	550	195	551	196
rect	550	196	551	197
rect	550	197	551	198
rect	550	198	551	199
rect	550	199	551	200
rect	550	200	551	201
rect	550	201	551	202
rect	550	202	551	203
rect	550	203	551	204
rect	550	204	551	205
rect	550	205	551	206
rect	550	206	551	207
rect	550	207	551	208
rect	550	208	551	209
rect	550	209	551	210
rect	550	210	551	211
rect	550	211	551	212
rect	550	212	551	213
rect	550	213	551	214
rect	550	214	551	215
rect	550	215	551	216
rect	550	216	551	217
rect	550	217	551	218
rect	550	218	551	219
rect	550	219	551	220
rect	550	220	551	221
rect	550	221	551	222
rect	550	222	551	223
rect	550	223	551	224
rect	550	224	551	225
rect	550	225	551	226
rect	550	226	551	227
rect	550	227	551	228
rect	550	228	551	229
rect	550	229	551	230
rect	550	230	551	231
rect	550	231	551	232
rect	550	232	551	233
rect	550	233	551	234
rect	550	234	551	235
rect	550	235	551	236
rect	550	236	551	237
rect	550	237	551	238
rect	550	238	551	239
rect	550	239	551	240
rect	550	240	551	241
rect	550	241	551	242
rect	550	242	551	243
rect	550	243	551	244
rect	550	244	551	245
rect	550	245	551	246
rect	550	246	551	247
rect	550	247	551	248
rect	550	248	551	249
rect	550	249	551	250
rect	550	250	551	251
rect	550	251	551	252
rect	550	252	551	253
rect	550	253	551	254
rect	550	254	551	255
rect	550	255	551	256
rect	550	256	551	257
rect	550	257	551	258
rect	550	258	551	259
rect	550	259	551	260
rect	550	260	551	261
rect	550	261	551	262
rect	550	262	551	263
rect	550	263	551	264
rect	550	264	551	265
rect	550	265	551	266
rect	550	266	551	267
rect	550	267	551	268
rect	550	268	551	269
rect	550	269	551	270
rect	550	270	551	271
rect	550	271	551	272
rect	550	272	551	273
rect	550	273	551	274
rect	550	274	551	275
rect	550	275	551	276
rect	550	276	551	277
rect	550	277	551	278
rect	550	278	551	279
rect	550	279	551	280
rect	550	280	551	281
rect	550	281	551	282
rect	550	282	551	283
rect	550	283	551	284
rect	550	284	551	285
rect	551	0	552	1
rect	551	1	552	2
rect	551	2	552	3
rect	551	3	552	4
rect	551	4	552	5
rect	551	5	552	6
rect	551	6	552	7
rect	551	7	552	8
rect	551	8	552	9
rect	551	9	552	10
rect	551	10	552	11
rect	551	11	552	12
rect	551	12	552	13
rect	551	13	552	14
rect	551	14	552	15
rect	551	15	552	16
rect	551	16	552	17
rect	551	17	552	18
rect	551	18	552	19
rect	551	19	552	20
rect	551	20	552	21
rect	551	21	552	22
rect	551	22	552	23
rect	551	23	552	24
rect	551	24	552	25
rect	551	25	552	26
rect	551	26	552	27
rect	551	27	552	28
rect	551	28	552	29
rect	551	29	552	30
rect	551	30	552	31
rect	551	31	552	32
rect	551	32	552	33
rect	551	33	552	34
rect	551	34	552	35
rect	551	35	552	36
rect	551	36	552	37
rect	551	37	552	38
rect	551	38	552	39
rect	551	39	552	40
rect	551	40	552	41
rect	551	41	552	42
rect	551	42	552	43
rect	551	43	552	44
rect	551	44	552	45
rect	551	45	552	46
rect	551	46	552	47
rect	551	47	552	48
rect	551	48	552	49
rect	551	49	552	50
rect	551	50	552	51
rect	551	51	552	52
rect	551	52	552	53
rect	551	53	552	54
rect	551	54	552	55
rect	551	55	552	56
rect	551	56	552	57
rect	551	57	552	58
rect	551	58	552	59
rect	551	59	552	60
rect	551	60	552	61
rect	551	61	552	62
rect	551	62	552	63
rect	551	63	552	64
rect	551	64	552	65
rect	551	65	552	66
rect	551	66	552	67
rect	551	67	552	68
rect	551	68	552	69
rect	551	69	552	70
rect	551	70	552	71
rect	551	71	552	72
rect	551	72	552	73
rect	551	73	552	74
rect	551	74	552	75
rect	551	75	552	76
rect	551	76	552	77
rect	551	77	552	78
rect	551	78	552	79
rect	551	79	552	80
rect	551	80	552	81
rect	551	81	552	82
rect	551	82	552	83
rect	551	83	552	84
rect	551	84	552	85
rect	551	85	552	86
rect	551	86	552	87
rect	551	87	552	88
rect	551	88	552	89
rect	551	89	552	90
rect	551	90	552	91
rect	551	91	552	92
rect	551	92	552	93
rect	551	93	552	94
rect	551	94	552	95
rect	551	95	552	96
rect	551	96	552	97
rect	551	97	552	98
rect	551	98	552	99
rect	551	99	552	100
rect	551	100	552	101
rect	551	101	552	102
rect	551	102	552	103
rect	551	103	552	104
rect	551	104	552	105
rect	551	105	552	106
rect	551	106	552	107
rect	551	107	552	108
rect	551	108	552	109
rect	551	109	552	110
rect	551	110	552	111
rect	551	111	552	112
rect	551	112	552	113
rect	551	113	552	114
rect	551	114	552	115
rect	551	115	552	116
rect	551	116	552	117
rect	551	117	552	118
rect	551	118	552	119
rect	551	119	552	120
rect	551	120	552	121
rect	551	121	552	122
rect	551	122	552	123
rect	551	123	552	124
rect	551	124	552	125
rect	551	125	552	126
rect	551	126	552	127
rect	551	127	552	128
rect	551	128	552	129
rect	551	129	552	130
rect	551	130	552	131
rect	551	131	552	132
rect	551	132	552	133
rect	551	133	552	134
rect	551	134	552	135
rect	551	135	552	136
rect	551	136	552	137
rect	551	137	552	138
rect	551	138	552	139
rect	551	139	552	140
rect	551	140	552	141
rect	551	141	552	142
rect	551	142	552	143
rect	551	143	552	144
rect	551	144	552	145
rect	551	145	552	146
rect	551	146	552	147
rect	551	147	552	148
rect	551	148	552	149
rect	551	149	552	150
rect	551	150	552	151
rect	551	151	552	152
rect	551	152	552	153
rect	551	153	552	154
rect	551	154	552	155
rect	551	155	552	156
rect	551	156	552	157
rect	551	157	552	158
rect	551	158	552	159
rect	551	159	552	160
rect	551	160	552	161
rect	551	161	552	162
rect	551	162	552	163
rect	551	163	552	164
rect	551	164	552	165
rect	551	165	552	166
rect	551	166	552	167
rect	551	167	552	168
rect	551	168	552	169
rect	551	169	552	170
rect	551	170	552	171
rect	551	171	552	172
rect	551	172	552	173
rect	551	173	552	174
rect	551	174	552	175
rect	551	175	552	176
rect	551	176	552	177
rect	551	177	552	178
rect	551	178	552	179
rect	551	179	552	180
rect	551	180	552	181
rect	551	181	552	182
rect	551	182	552	183
rect	551	183	552	184
rect	551	184	552	185
rect	551	185	552	186
rect	551	186	552	187
rect	551	187	552	188
rect	551	188	552	189
rect	551	189	552	190
rect	551	190	552	191
rect	551	191	552	192
rect	551	192	552	193
rect	551	193	552	194
rect	551	194	552	195
rect	551	195	552	196
rect	551	196	552	197
rect	551	197	552	198
rect	551	198	552	199
rect	551	199	552	200
rect	551	200	552	201
rect	551	201	552	202
rect	551	202	552	203
rect	551	203	552	204
rect	551	204	552	205
rect	551	205	552	206
rect	551	206	552	207
rect	551	207	552	208
rect	551	208	552	209
rect	551	209	552	210
rect	551	210	552	211
rect	551	211	552	212
rect	551	212	552	213
rect	551	213	552	214
rect	551	214	552	215
rect	551	215	552	216
rect	551	216	552	217
rect	551	217	552	218
rect	551	218	552	219
rect	551	219	552	220
rect	551	220	552	221
rect	551	221	552	222
rect	551	222	552	223
rect	551	223	552	224
rect	551	224	552	225
rect	551	225	552	226
rect	551	226	552	227
rect	551	227	552	228
rect	551	228	552	229
rect	551	229	552	230
rect	551	230	552	231
rect	551	231	552	232
rect	551	232	552	233
rect	551	233	552	234
rect	551	234	552	235
rect	551	235	552	236
rect	551	236	552	237
rect	551	237	552	238
rect	551	238	552	239
rect	551	239	552	240
rect	551	240	552	241
rect	551	241	552	242
rect	551	242	552	243
rect	551	243	552	244
rect	551	244	552	245
rect	551	245	552	246
rect	551	246	552	247
rect	551	247	552	248
rect	551	248	552	249
rect	551	249	552	250
rect	551	250	552	251
rect	551	251	552	252
rect	551	252	552	253
rect	551	253	552	254
rect	551	254	552	255
rect	551	255	552	256
rect	551	256	552	257
rect	551	257	552	258
rect	551	258	552	259
rect	551	259	552	260
rect	551	260	552	261
rect	551	261	552	262
rect	551	262	552	263
rect	551	263	552	264
rect	551	264	552	265
rect	551	265	552	266
rect	551	266	552	267
rect	551	267	552	268
rect	551	268	552	269
rect	551	269	552	270
rect	551	270	552	271
rect	551	271	552	272
rect	551	272	552	273
rect	551	273	552	274
rect	551	274	552	275
rect	551	275	552	276
rect	551	276	552	277
rect	551	277	552	278
rect	551	278	552	279
rect	551	279	552	280
rect	551	280	552	281
rect	551	281	552	282
rect	551	282	552	283
rect	551	283	552	284
rect	551	284	552	285
rect	552	0	553	1
rect	552	1	553	2
rect	552	2	553	3
rect	552	3	553	4
rect	552	4	553	5
rect	552	5	553	6
rect	552	6	553	7
rect	552	7	553	8
rect	552	8	553	9
rect	552	9	553	10
rect	552	10	553	11
rect	552	11	553	12
rect	552	12	553	13
rect	552	13	553	14
rect	552	14	553	15
rect	552	15	553	16
rect	552	16	553	17
rect	552	17	553	18
rect	552	18	553	19
rect	552	19	553	20
rect	552	20	553	21
rect	552	21	553	22
rect	552	22	553	23
rect	552	23	553	24
rect	552	24	553	25
rect	552	25	553	26
rect	552	26	553	27
rect	552	27	553	28
rect	552	28	553	29
rect	552	29	553	30
rect	552	30	553	31
rect	552	31	553	32
rect	552	32	553	33
rect	552	33	553	34
rect	552	34	553	35
rect	552	35	553	36
rect	552	36	553	37
rect	552	37	553	38
rect	552	38	553	39
rect	552	39	553	40
rect	552	40	553	41
rect	552	41	553	42
rect	552	42	553	43
rect	552	43	553	44
rect	552	44	553	45
rect	552	45	553	46
rect	552	46	553	47
rect	552	47	553	48
rect	552	48	553	49
rect	552	49	553	50
rect	552	50	553	51
rect	552	51	553	52
rect	552	52	553	53
rect	552	53	553	54
rect	552	54	553	55
rect	552	55	553	56
rect	552	56	553	57
rect	552	57	553	58
rect	552	58	553	59
rect	552	59	553	60
rect	552	60	553	61
rect	552	61	553	62
rect	552	62	553	63
rect	552	63	553	64
rect	552	64	553	65
rect	552	65	553	66
rect	552	66	553	67
rect	552	67	553	68
rect	552	68	553	69
rect	552	69	553	70
rect	552	70	553	71
rect	552	71	553	72
rect	552	72	553	73
rect	552	73	553	74
rect	552	74	553	75
rect	552	75	553	76
rect	552	76	553	77
rect	552	77	553	78
rect	552	78	553	79
rect	552	79	553	80
rect	552	80	553	81
rect	552	81	553	82
rect	552	82	553	83
rect	552	83	553	84
rect	552	84	553	85
rect	552	85	553	86
rect	552	86	553	87
rect	552	87	553	88
rect	552	88	553	89
rect	552	89	553	90
rect	552	90	553	91
rect	552	91	553	92
rect	552	92	553	93
rect	552	93	553	94
rect	552	94	553	95
rect	552	95	553	96
rect	552	96	553	97
rect	552	97	553	98
rect	552	98	553	99
rect	552	99	553	100
rect	552	100	553	101
rect	552	101	553	102
rect	552	102	553	103
rect	552	103	553	104
rect	552	104	553	105
rect	552	105	553	106
rect	552	106	553	107
rect	552	107	553	108
rect	552	108	553	109
rect	552	109	553	110
rect	552	110	553	111
rect	552	111	553	112
rect	552	112	553	113
rect	552	113	553	114
rect	552	114	553	115
rect	552	115	553	116
rect	552	116	553	117
rect	552	117	553	118
rect	552	118	553	119
rect	552	119	553	120
rect	552	120	553	121
rect	552	121	553	122
rect	552	122	553	123
rect	552	123	553	124
rect	552	124	553	125
rect	552	125	553	126
rect	552	126	553	127
rect	552	127	553	128
rect	552	128	553	129
rect	552	129	553	130
rect	552	130	553	131
rect	552	131	553	132
rect	552	132	553	133
rect	552	133	553	134
rect	552	134	553	135
rect	552	135	553	136
rect	552	136	553	137
rect	552	137	553	138
rect	552	138	553	139
rect	552	139	553	140
rect	552	140	553	141
rect	552	141	553	142
rect	552	142	553	143
rect	552	143	553	144
rect	552	144	553	145
rect	552	145	553	146
rect	552	146	553	147
rect	552	147	553	148
rect	552	148	553	149
rect	552	149	553	150
rect	552	150	553	151
rect	552	151	553	152
rect	552	152	553	153
rect	552	153	553	154
rect	552	154	553	155
rect	552	155	553	156
rect	552	156	553	157
rect	552	157	553	158
rect	552	158	553	159
rect	552	159	553	160
rect	552	160	553	161
rect	552	161	553	162
rect	552	162	553	163
rect	552	163	553	164
rect	552	164	553	165
rect	552	165	553	166
rect	552	166	553	167
rect	552	167	553	168
rect	552	168	553	169
rect	552	169	553	170
rect	552	170	553	171
rect	552	171	553	172
rect	552	172	553	173
rect	552	173	553	174
rect	552	174	553	175
rect	552	175	553	176
rect	552	176	553	177
rect	552	177	553	178
rect	552	178	553	179
rect	552	179	553	180
rect	552	180	553	181
rect	552	181	553	182
rect	552	182	553	183
rect	552	183	553	184
rect	552	184	553	185
rect	552	185	553	186
rect	552	186	553	187
rect	552	187	553	188
rect	552	188	553	189
rect	552	189	553	190
rect	552	190	553	191
rect	552	191	553	192
rect	552	192	553	193
rect	552	193	553	194
rect	552	194	553	195
rect	552	195	553	196
rect	552	196	553	197
rect	552	197	553	198
rect	552	198	553	199
rect	552	199	553	200
rect	552	200	553	201
rect	552	201	553	202
rect	552	202	553	203
rect	552	203	553	204
rect	552	204	553	205
rect	552	205	553	206
rect	552	206	553	207
rect	552	207	553	208
rect	552	208	553	209
rect	552	209	553	210
rect	552	210	553	211
rect	552	211	553	212
rect	552	212	553	213
rect	552	213	553	214
rect	552	214	553	215
rect	552	215	553	216
rect	552	216	553	217
rect	552	217	553	218
rect	552	218	553	219
rect	552	219	553	220
rect	552	220	553	221
rect	552	221	553	222
rect	552	222	553	223
rect	552	223	553	224
rect	552	224	553	225
rect	552	225	553	226
rect	552	226	553	227
rect	552	227	553	228
rect	552	228	553	229
rect	552	229	553	230
rect	552	230	553	231
rect	552	231	553	232
rect	552	232	553	233
rect	552	233	553	234
rect	552	234	553	235
rect	552	235	553	236
rect	552	236	553	237
rect	552	237	553	238
rect	552	238	553	239
rect	552	239	553	240
rect	552	240	553	241
rect	552	241	553	242
rect	552	242	553	243
rect	552	243	553	244
rect	552	244	553	245
rect	552	245	553	246
rect	552	246	553	247
rect	552	247	553	248
rect	552	248	553	249
rect	552	249	553	250
rect	552	250	553	251
rect	552	251	553	252
rect	552	252	553	253
rect	552	253	553	254
rect	552	254	553	255
rect	552	255	553	256
rect	552	256	553	257
rect	552	257	553	258
rect	552	258	553	259
rect	552	259	553	260
rect	552	260	553	261
rect	552	261	553	262
rect	552	262	553	263
rect	552	263	553	264
rect	552	264	553	265
rect	552	265	553	266
rect	552	266	553	267
rect	552	267	553	268
rect	552	268	553	269
rect	552	269	553	270
rect	552	270	553	271
rect	552	271	553	272
rect	552	272	553	273
rect	552	273	553	274
rect	552	274	553	275
rect	552	275	553	276
rect	552	276	553	277
rect	552	277	553	278
rect	552	278	553	279
rect	552	279	553	280
rect	552	280	553	281
rect	552	281	553	282
rect	552	282	553	283
rect	552	283	553	284
rect	552	284	553	285
rect	570	0	571	1
rect	570	1	571	2
rect	570	2	571	3
rect	570	3	571	4
rect	570	4	571	5
rect	570	5	571	6
rect	570	6	571	7
rect	570	7	571	8
rect	570	8	571	9
rect	570	9	571	10
rect	570	10	571	11
rect	570	11	571	12
rect	570	12	571	13
rect	570	13	571	14
rect	570	14	571	15
rect	570	15	571	16
rect	570	16	571	17
rect	570	17	571	18
rect	570	18	571	19
rect	570	19	571	20
rect	570	20	571	21
rect	570	21	571	22
rect	570	22	571	23
rect	570	23	571	24
rect	570	24	571	25
rect	570	25	571	26
rect	570	26	571	27
rect	570	27	571	28
rect	570	28	571	29
rect	570	29	571	30
rect	570	30	571	31
rect	570	31	571	32
rect	570	32	571	33
rect	570	33	571	34
rect	570	34	571	35
rect	570	35	571	36
rect	570	36	571	37
rect	570	37	571	38
rect	570	38	571	39
rect	570	39	571	40
rect	570	40	571	41
rect	570	41	571	42
rect	570	42	571	43
rect	570	43	571	44
rect	570	44	571	45
rect	570	45	571	46
rect	570	46	571	47
rect	570	47	571	48
rect	570	48	571	49
rect	570	49	571	50
rect	570	50	571	51
rect	570	51	571	52
rect	570	52	571	53
rect	570	53	571	54
rect	570	54	571	55
rect	570	55	571	56
rect	570	56	571	57
rect	570	57	571	58
rect	570	58	571	59
rect	570	59	571	60
rect	570	60	571	61
rect	570	61	571	62
rect	570	62	571	63
rect	570	63	571	64
rect	570	64	571	65
rect	570	65	571	66
rect	570	66	571	67
rect	570	67	571	68
rect	570	68	571	69
rect	570	69	571	70
rect	570	70	571	71
rect	570	71	571	72
rect	570	72	571	73
rect	570	73	571	74
rect	570	74	571	75
rect	570	75	571	76
rect	570	76	571	77
rect	570	77	571	78
rect	570	78	571	79
rect	570	79	571	80
rect	570	80	571	81
rect	570	81	571	82
rect	570	82	571	83
rect	570	83	571	84
rect	570	84	571	85
rect	570	85	571	86
rect	570	86	571	87
rect	570	87	571	88
rect	570	88	571	89
rect	570	89	571	90
rect	570	90	571	91
rect	570	91	571	92
rect	570	92	571	93
rect	570	93	571	94
rect	570	94	571	95
rect	570	95	571	96
rect	570	96	571	97
rect	570	97	571	98
rect	570	98	571	99
rect	570	99	571	100
rect	570	100	571	101
rect	570	101	571	102
rect	570	102	571	103
rect	570	103	571	104
rect	570	104	571	105
rect	570	105	571	106
rect	570	106	571	107
rect	570	107	571	108
rect	570	108	571	109
rect	570	109	571	110
rect	570	110	571	111
rect	570	111	571	112
rect	570	112	571	113
rect	570	113	571	114
rect	570	114	571	115
rect	570	115	571	116
rect	570	116	571	117
rect	570	117	571	118
rect	570	118	571	119
rect	570	119	571	120
rect	570	120	571	121
rect	570	121	571	122
rect	570	122	571	123
rect	570	123	571	124
rect	570	124	571	125
rect	570	125	571	126
rect	570	126	571	127
rect	570	127	571	128
rect	570	128	571	129
rect	570	129	571	130
rect	570	130	571	131
rect	570	131	571	132
rect	570	132	571	133
rect	570	133	571	134
rect	570	134	571	135
rect	570	135	571	136
rect	570	136	571	137
rect	570	137	571	138
rect	570	138	571	139
rect	570	139	571	140
rect	570	140	571	141
rect	570	141	571	142
rect	570	142	571	143
rect	570	143	571	144
rect	570	144	571	145
rect	570	145	571	146
rect	570	146	571	147
rect	570	147	571	148
rect	570	148	571	149
rect	570	149	571	150
rect	570	150	571	151
rect	570	151	571	152
rect	570	152	571	153
rect	570	153	571	154
rect	570	154	571	155
rect	570	155	571	156
rect	570	156	571	157
rect	570	157	571	158
rect	570	158	571	159
rect	570	159	571	160
rect	570	160	571	161
rect	570	161	571	162
rect	570	162	571	163
rect	570	163	571	164
rect	570	164	571	165
rect	570	165	571	166
rect	570	166	571	167
rect	570	167	571	168
rect	570	168	571	169
rect	570	169	571	170
rect	570	170	571	171
rect	570	171	571	172
rect	570	172	571	173
rect	570	173	571	174
rect	570	174	571	175
rect	570	175	571	176
rect	570	176	571	177
rect	570	177	571	178
rect	570	178	571	179
rect	570	179	571	180
rect	570	180	571	181
rect	570	181	571	182
rect	570	182	571	183
rect	570	183	571	184
rect	570	184	571	185
rect	570	185	571	186
rect	570	186	571	187
rect	570	187	571	188
rect	570	188	571	189
rect	570	189	571	190
rect	570	190	571	191
rect	570	191	571	192
rect	570	192	571	193
rect	570	193	571	194
rect	570	194	571	195
rect	570	195	571	196
rect	570	196	571	197
rect	570	197	571	198
rect	570	198	571	199
rect	570	199	571	200
rect	570	200	571	201
rect	570	201	571	202
rect	570	202	571	203
rect	570	203	571	204
rect	570	204	571	205
rect	570	205	571	206
rect	570	206	571	207
rect	570	207	571	208
rect	570	208	571	209
rect	570	209	571	210
rect	570	210	571	211
rect	570	211	571	212
rect	570	212	571	213
rect	570	213	571	214
rect	570	214	571	215
rect	570	215	571	216
rect	570	216	571	217
rect	570	217	571	218
rect	570	218	571	219
rect	570	219	571	220
rect	570	220	571	221
rect	570	221	571	222
rect	570	222	571	223
rect	570	223	571	224
rect	570	224	571	225
rect	570	225	571	226
rect	570	226	571	227
rect	570	227	571	228
rect	570	228	571	229
rect	570	229	571	230
rect	570	230	571	231
rect	570	231	571	232
rect	570	232	571	233
rect	570	233	571	234
rect	570	234	571	235
rect	570	235	571	236
rect	570	236	571	237
rect	570	237	571	238
rect	570	238	571	239
rect	570	239	571	240
rect	570	240	571	241
rect	570	241	571	242
rect	570	242	571	243
rect	570	243	571	244
rect	570	244	571	245
rect	570	245	571	246
rect	570	246	571	247
rect	570	247	571	248
rect	570	248	571	249
rect	570	249	571	250
rect	570	250	571	251
rect	570	251	571	252
rect	570	252	571	253
rect	570	253	571	254
rect	570	254	571	255
rect	570	255	571	256
rect	570	256	571	257
rect	570	257	571	258
rect	570	258	571	259
rect	570	259	571	260
rect	570	260	571	261
rect	570	261	571	262
rect	570	262	571	263
rect	570	263	571	264
rect	570	264	571	265
rect	570	265	571	266
rect	570	266	571	267
rect	570	267	571	268
rect	570	268	571	269
rect	570	269	571	270
rect	571	0	572	1
rect	571	1	572	2
rect	571	2	572	3
rect	571	3	572	4
rect	571	4	572	5
rect	571	5	572	6
rect	571	6	572	7
rect	571	7	572	8
rect	571	8	572	9
rect	571	9	572	10
rect	571	10	572	11
rect	571	11	572	12
rect	571	12	572	13
rect	571	13	572	14
rect	571	14	572	15
rect	571	15	572	16
rect	571	16	572	17
rect	571	17	572	18
rect	571	18	572	19
rect	571	19	572	20
rect	571	20	572	21
rect	571	21	572	22
rect	571	22	572	23
rect	571	23	572	24
rect	571	24	572	25
rect	571	25	572	26
rect	571	26	572	27
rect	571	27	572	28
rect	571	28	572	29
rect	571	29	572	30
rect	571	30	572	31
rect	571	31	572	32
rect	571	32	572	33
rect	571	33	572	34
rect	571	34	572	35
rect	571	35	572	36
rect	571	36	572	37
rect	571	37	572	38
rect	571	38	572	39
rect	571	39	572	40
rect	571	40	572	41
rect	571	41	572	42
rect	571	42	572	43
rect	571	43	572	44
rect	571	44	572	45
rect	571	45	572	46
rect	571	46	572	47
rect	571	47	572	48
rect	571	48	572	49
rect	571	49	572	50
rect	571	50	572	51
rect	571	51	572	52
rect	571	52	572	53
rect	571	53	572	54
rect	571	54	572	55
rect	571	55	572	56
rect	571	56	572	57
rect	571	57	572	58
rect	571	58	572	59
rect	571	59	572	60
rect	571	60	572	61
rect	571	61	572	62
rect	571	62	572	63
rect	571	63	572	64
rect	571	64	572	65
rect	571	65	572	66
rect	571	66	572	67
rect	571	67	572	68
rect	571	68	572	69
rect	571	69	572	70
rect	571	70	572	71
rect	571	71	572	72
rect	571	72	572	73
rect	571	73	572	74
rect	571	74	572	75
rect	571	75	572	76
rect	571	76	572	77
rect	571	77	572	78
rect	571	78	572	79
rect	571	79	572	80
rect	571	80	572	81
rect	571	81	572	82
rect	571	82	572	83
rect	571	83	572	84
rect	571	84	572	85
rect	571	85	572	86
rect	571	86	572	87
rect	571	87	572	88
rect	571	88	572	89
rect	571	89	572	90
rect	571	90	572	91
rect	571	91	572	92
rect	571	92	572	93
rect	571	93	572	94
rect	571	94	572	95
rect	571	95	572	96
rect	571	96	572	97
rect	571	97	572	98
rect	571	98	572	99
rect	571	99	572	100
rect	571	100	572	101
rect	571	101	572	102
rect	571	102	572	103
rect	571	103	572	104
rect	571	104	572	105
rect	571	105	572	106
rect	571	106	572	107
rect	571	107	572	108
rect	571	108	572	109
rect	571	109	572	110
rect	571	110	572	111
rect	571	111	572	112
rect	571	112	572	113
rect	571	113	572	114
rect	571	114	572	115
rect	571	115	572	116
rect	571	116	572	117
rect	571	117	572	118
rect	571	118	572	119
rect	571	119	572	120
rect	571	120	572	121
rect	571	121	572	122
rect	571	122	572	123
rect	571	123	572	124
rect	571	124	572	125
rect	571	125	572	126
rect	571	126	572	127
rect	571	127	572	128
rect	571	128	572	129
rect	571	129	572	130
rect	571	130	572	131
rect	571	131	572	132
rect	571	132	572	133
rect	571	133	572	134
rect	571	134	572	135
rect	571	135	572	136
rect	571	136	572	137
rect	571	137	572	138
rect	571	138	572	139
rect	571	139	572	140
rect	571	140	572	141
rect	571	141	572	142
rect	571	142	572	143
rect	571	143	572	144
rect	571	144	572	145
rect	571	145	572	146
rect	571	146	572	147
rect	571	147	572	148
rect	571	148	572	149
rect	571	149	572	150
rect	571	150	572	151
rect	571	151	572	152
rect	571	152	572	153
rect	571	153	572	154
rect	571	154	572	155
rect	571	155	572	156
rect	571	156	572	157
rect	571	157	572	158
rect	571	158	572	159
rect	571	159	572	160
rect	571	160	572	161
rect	571	161	572	162
rect	571	162	572	163
rect	571	163	572	164
rect	571	164	572	165
rect	571	165	572	166
rect	571	166	572	167
rect	571	167	572	168
rect	571	168	572	169
rect	571	169	572	170
rect	571	170	572	171
rect	571	171	572	172
rect	571	172	572	173
rect	571	173	572	174
rect	571	174	572	175
rect	571	175	572	176
rect	571	176	572	177
rect	571	177	572	178
rect	571	178	572	179
rect	571	179	572	180
rect	571	180	572	181
rect	571	181	572	182
rect	571	182	572	183
rect	571	183	572	184
rect	571	184	572	185
rect	571	185	572	186
rect	571	186	572	187
rect	571	187	572	188
rect	571	188	572	189
rect	571	189	572	190
rect	571	190	572	191
rect	571	191	572	192
rect	571	192	572	193
rect	571	193	572	194
rect	571	194	572	195
rect	571	195	572	196
rect	571	196	572	197
rect	571	197	572	198
rect	571	198	572	199
rect	571	199	572	200
rect	571	200	572	201
rect	571	201	572	202
rect	571	202	572	203
rect	571	203	572	204
rect	571	204	572	205
rect	571	205	572	206
rect	571	206	572	207
rect	571	207	572	208
rect	571	208	572	209
rect	571	209	572	210
rect	571	210	572	211
rect	571	211	572	212
rect	571	212	572	213
rect	571	213	572	214
rect	571	214	572	215
rect	571	215	572	216
rect	571	216	572	217
rect	571	217	572	218
rect	571	218	572	219
rect	571	219	572	220
rect	571	220	572	221
rect	571	221	572	222
rect	571	222	572	223
rect	571	223	572	224
rect	571	224	572	225
rect	571	225	572	226
rect	571	226	572	227
rect	571	227	572	228
rect	571	228	572	229
rect	571	229	572	230
rect	571	230	572	231
rect	571	231	572	232
rect	571	232	572	233
rect	571	233	572	234
rect	571	234	572	235
rect	571	235	572	236
rect	571	236	572	237
rect	571	237	572	238
rect	571	238	572	239
rect	571	239	572	240
rect	571	240	572	241
rect	571	241	572	242
rect	571	242	572	243
rect	571	243	572	244
rect	571	244	572	245
rect	571	245	572	246
rect	571	246	572	247
rect	571	247	572	248
rect	571	248	572	249
rect	571	249	572	250
rect	571	250	572	251
rect	571	251	572	252
rect	571	252	572	253
rect	571	253	572	254
rect	571	254	572	255
rect	571	255	572	256
rect	571	256	572	257
rect	571	257	572	258
rect	571	258	572	259
rect	571	259	572	260
rect	571	260	572	261
rect	571	261	572	262
rect	571	262	572	263
rect	571	263	572	264
rect	571	264	572	265
rect	571	265	572	266
rect	571	266	572	267
rect	571	267	572	268
rect	571	268	572	269
rect	571	269	572	270
rect	572	0	573	1
rect	572	1	573	2
rect	572	2	573	3
rect	572	3	573	4
rect	572	4	573	5
rect	572	5	573	6
rect	572	6	573	7
rect	572	7	573	8
rect	572	8	573	9
rect	572	9	573	10
rect	572	10	573	11
rect	572	11	573	12
rect	572	12	573	13
rect	572	13	573	14
rect	572	14	573	15
rect	572	15	573	16
rect	572	16	573	17
rect	572	17	573	18
rect	572	18	573	19
rect	572	19	573	20
rect	572	20	573	21
rect	572	21	573	22
rect	572	22	573	23
rect	572	23	573	24
rect	572	24	573	25
rect	572	25	573	26
rect	572	26	573	27
rect	572	27	573	28
rect	572	28	573	29
rect	572	29	573	30
rect	572	30	573	31
rect	572	31	573	32
rect	572	32	573	33
rect	572	33	573	34
rect	572	34	573	35
rect	572	35	573	36
rect	572	36	573	37
rect	572	37	573	38
rect	572	38	573	39
rect	572	39	573	40
rect	572	40	573	41
rect	572	41	573	42
rect	572	42	573	43
rect	572	43	573	44
rect	572	44	573	45
rect	572	45	573	46
rect	572	46	573	47
rect	572	47	573	48
rect	572	48	573	49
rect	572	49	573	50
rect	572	50	573	51
rect	572	51	573	52
rect	572	52	573	53
rect	572	53	573	54
rect	572	54	573	55
rect	572	55	573	56
rect	572	56	573	57
rect	572	57	573	58
rect	572	58	573	59
rect	572	59	573	60
rect	572	60	573	61
rect	572	61	573	62
rect	572	62	573	63
rect	572	63	573	64
rect	572	64	573	65
rect	572	65	573	66
rect	572	66	573	67
rect	572	67	573	68
rect	572	68	573	69
rect	572	69	573	70
rect	572	70	573	71
rect	572	71	573	72
rect	572	72	573	73
rect	572	73	573	74
rect	572	74	573	75
rect	572	75	573	76
rect	572	76	573	77
rect	572	77	573	78
rect	572	78	573	79
rect	572	79	573	80
rect	572	80	573	81
rect	572	81	573	82
rect	572	82	573	83
rect	572	83	573	84
rect	572	84	573	85
rect	572	85	573	86
rect	572	86	573	87
rect	572	87	573	88
rect	572	88	573	89
rect	572	89	573	90
rect	572	90	573	91
rect	572	91	573	92
rect	572	92	573	93
rect	572	93	573	94
rect	572	94	573	95
rect	572	95	573	96
rect	572	96	573	97
rect	572	97	573	98
rect	572	98	573	99
rect	572	99	573	100
rect	572	100	573	101
rect	572	101	573	102
rect	572	102	573	103
rect	572	103	573	104
rect	572	104	573	105
rect	572	105	573	106
rect	572	106	573	107
rect	572	107	573	108
rect	572	108	573	109
rect	572	109	573	110
rect	572	110	573	111
rect	572	111	573	112
rect	572	112	573	113
rect	572	113	573	114
rect	572	114	573	115
rect	572	115	573	116
rect	572	116	573	117
rect	572	117	573	118
rect	572	118	573	119
rect	572	119	573	120
rect	572	120	573	121
rect	572	121	573	122
rect	572	122	573	123
rect	572	123	573	124
rect	572	124	573	125
rect	572	125	573	126
rect	572	126	573	127
rect	572	127	573	128
rect	572	128	573	129
rect	572	129	573	130
rect	572	130	573	131
rect	572	131	573	132
rect	572	132	573	133
rect	572	133	573	134
rect	572	134	573	135
rect	572	135	573	136
rect	572	136	573	137
rect	572	137	573	138
rect	572	138	573	139
rect	572	139	573	140
rect	572	140	573	141
rect	572	141	573	142
rect	572	142	573	143
rect	572	143	573	144
rect	572	144	573	145
rect	572	145	573	146
rect	572	146	573	147
rect	572	147	573	148
rect	572	148	573	149
rect	572	149	573	150
rect	572	150	573	151
rect	572	151	573	152
rect	572	152	573	153
rect	572	153	573	154
rect	572	154	573	155
rect	572	155	573	156
rect	572	156	573	157
rect	572	157	573	158
rect	572	158	573	159
rect	572	159	573	160
rect	572	160	573	161
rect	572	161	573	162
rect	572	162	573	163
rect	572	163	573	164
rect	572	164	573	165
rect	572	165	573	166
rect	572	166	573	167
rect	572	167	573	168
rect	572	168	573	169
rect	572	169	573	170
rect	572	170	573	171
rect	572	171	573	172
rect	572	172	573	173
rect	572	173	573	174
rect	572	174	573	175
rect	572	175	573	176
rect	572	176	573	177
rect	572	177	573	178
rect	572	178	573	179
rect	572	179	573	180
rect	572	180	573	181
rect	572	181	573	182
rect	572	182	573	183
rect	572	183	573	184
rect	572	184	573	185
rect	572	185	573	186
rect	572	186	573	187
rect	572	187	573	188
rect	572	188	573	189
rect	572	189	573	190
rect	572	190	573	191
rect	572	191	573	192
rect	572	192	573	193
rect	572	193	573	194
rect	572	194	573	195
rect	572	195	573	196
rect	572	196	573	197
rect	572	197	573	198
rect	572	198	573	199
rect	572	199	573	200
rect	572	200	573	201
rect	572	201	573	202
rect	572	202	573	203
rect	572	203	573	204
rect	572	204	573	205
rect	572	205	573	206
rect	572	206	573	207
rect	572	207	573	208
rect	572	208	573	209
rect	572	209	573	210
rect	572	210	573	211
rect	572	211	573	212
rect	572	212	573	213
rect	572	213	573	214
rect	572	214	573	215
rect	572	215	573	216
rect	572	216	573	217
rect	572	217	573	218
rect	572	218	573	219
rect	572	219	573	220
rect	572	220	573	221
rect	572	221	573	222
rect	572	222	573	223
rect	572	223	573	224
rect	572	224	573	225
rect	572	225	573	226
rect	572	226	573	227
rect	572	227	573	228
rect	572	228	573	229
rect	572	229	573	230
rect	572	230	573	231
rect	572	231	573	232
rect	572	232	573	233
rect	572	233	573	234
rect	572	234	573	235
rect	572	235	573	236
rect	572	236	573	237
rect	572	237	573	238
rect	572	238	573	239
rect	572	239	573	240
rect	572	240	573	241
rect	572	241	573	242
rect	572	242	573	243
rect	572	243	573	244
rect	572	244	573	245
rect	572	245	573	246
rect	572	246	573	247
rect	572	247	573	248
rect	572	248	573	249
rect	572	249	573	250
rect	572	250	573	251
rect	572	251	573	252
rect	572	252	573	253
rect	572	253	573	254
rect	572	254	573	255
rect	572	255	573	256
rect	572	256	573	257
rect	572	257	573	258
rect	572	258	573	259
rect	572	259	573	260
rect	572	260	573	261
rect	572	261	573	262
rect	572	262	573	263
rect	572	263	573	264
rect	572	264	573	265
rect	572	265	573	266
rect	572	266	573	267
rect	572	267	573	268
rect	572	268	573	269
rect	572	269	573	270
rect	573	0	574	1
rect	573	1	574	2
rect	573	2	574	3
rect	573	3	574	4
rect	573	4	574	5
rect	573	5	574	6
rect	573	6	574	7
rect	573	7	574	8
rect	573	8	574	9
rect	573	9	574	10
rect	573	10	574	11
rect	573	11	574	12
rect	573	12	574	13
rect	573	13	574	14
rect	573	14	574	15
rect	573	15	574	16
rect	573	16	574	17
rect	573	17	574	18
rect	573	18	574	19
rect	573	19	574	20
rect	573	20	574	21
rect	573	21	574	22
rect	573	22	574	23
rect	573	23	574	24
rect	573	24	574	25
rect	573	25	574	26
rect	573	26	574	27
rect	573	27	574	28
rect	573	28	574	29
rect	573	29	574	30
rect	573	30	574	31
rect	573	31	574	32
rect	573	32	574	33
rect	573	33	574	34
rect	573	34	574	35
rect	573	35	574	36
rect	573	36	574	37
rect	573	37	574	38
rect	573	38	574	39
rect	573	39	574	40
rect	573	40	574	41
rect	573	41	574	42
rect	573	42	574	43
rect	573	43	574	44
rect	573	44	574	45
rect	573	45	574	46
rect	573	46	574	47
rect	573	47	574	48
rect	573	48	574	49
rect	573	49	574	50
rect	573	50	574	51
rect	573	51	574	52
rect	573	52	574	53
rect	573	53	574	54
rect	573	54	574	55
rect	573	55	574	56
rect	573	56	574	57
rect	573	57	574	58
rect	573	58	574	59
rect	573	59	574	60
rect	573	60	574	61
rect	573	61	574	62
rect	573	62	574	63
rect	573	63	574	64
rect	573	64	574	65
rect	573	65	574	66
rect	573	66	574	67
rect	573	67	574	68
rect	573	68	574	69
rect	573	69	574	70
rect	573	70	574	71
rect	573	71	574	72
rect	573	72	574	73
rect	573	73	574	74
rect	573	74	574	75
rect	573	75	574	76
rect	573	76	574	77
rect	573	77	574	78
rect	573	78	574	79
rect	573	79	574	80
rect	573	80	574	81
rect	573	81	574	82
rect	573	82	574	83
rect	573	83	574	84
rect	573	84	574	85
rect	573	85	574	86
rect	573	86	574	87
rect	573	87	574	88
rect	573	88	574	89
rect	573	89	574	90
rect	573	90	574	91
rect	573	91	574	92
rect	573	92	574	93
rect	573	93	574	94
rect	573	94	574	95
rect	573	95	574	96
rect	573	96	574	97
rect	573	97	574	98
rect	573	98	574	99
rect	573	99	574	100
rect	573	100	574	101
rect	573	101	574	102
rect	573	102	574	103
rect	573	103	574	104
rect	573	104	574	105
rect	573	105	574	106
rect	573	106	574	107
rect	573	107	574	108
rect	573	108	574	109
rect	573	109	574	110
rect	573	110	574	111
rect	573	111	574	112
rect	573	112	574	113
rect	573	113	574	114
rect	573	114	574	115
rect	573	115	574	116
rect	573	116	574	117
rect	573	117	574	118
rect	573	118	574	119
rect	573	119	574	120
rect	573	120	574	121
rect	573	121	574	122
rect	573	122	574	123
rect	573	123	574	124
rect	573	124	574	125
rect	573	125	574	126
rect	573	126	574	127
rect	573	127	574	128
rect	573	128	574	129
rect	573	129	574	130
rect	573	130	574	131
rect	573	131	574	132
rect	573	132	574	133
rect	573	133	574	134
rect	573	134	574	135
rect	573	135	574	136
rect	573	136	574	137
rect	573	137	574	138
rect	573	138	574	139
rect	573	139	574	140
rect	573	140	574	141
rect	573	141	574	142
rect	573	142	574	143
rect	573	143	574	144
rect	573	144	574	145
rect	573	145	574	146
rect	573	146	574	147
rect	573	147	574	148
rect	573	148	574	149
rect	573	149	574	150
rect	573	150	574	151
rect	573	151	574	152
rect	573	152	574	153
rect	573	153	574	154
rect	573	154	574	155
rect	573	155	574	156
rect	573	156	574	157
rect	573	157	574	158
rect	573	158	574	159
rect	573	159	574	160
rect	573	160	574	161
rect	573	161	574	162
rect	573	162	574	163
rect	573	163	574	164
rect	573	164	574	165
rect	573	165	574	166
rect	573	166	574	167
rect	573	167	574	168
rect	573	168	574	169
rect	573	169	574	170
rect	573	170	574	171
rect	573	171	574	172
rect	573	172	574	173
rect	573	173	574	174
rect	573	174	574	175
rect	573	175	574	176
rect	573	176	574	177
rect	573	177	574	178
rect	573	178	574	179
rect	573	179	574	180
rect	573	180	574	181
rect	573	181	574	182
rect	573	182	574	183
rect	573	183	574	184
rect	573	184	574	185
rect	573	185	574	186
rect	573	186	574	187
rect	573	187	574	188
rect	573	188	574	189
rect	573	189	574	190
rect	573	190	574	191
rect	573	191	574	192
rect	573	192	574	193
rect	573	193	574	194
rect	573	194	574	195
rect	573	195	574	196
rect	573	196	574	197
rect	573	197	574	198
rect	573	198	574	199
rect	573	199	574	200
rect	573	200	574	201
rect	573	201	574	202
rect	573	202	574	203
rect	573	203	574	204
rect	573	204	574	205
rect	573	205	574	206
rect	573	206	574	207
rect	573	207	574	208
rect	573	208	574	209
rect	573	209	574	210
rect	573	210	574	211
rect	573	211	574	212
rect	573	212	574	213
rect	573	213	574	214
rect	573	214	574	215
rect	573	215	574	216
rect	573	216	574	217
rect	573	217	574	218
rect	573	218	574	219
rect	573	219	574	220
rect	573	220	574	221
rect	573	221	574	222
rect	573	222	574	223
rect	573	223	574	224
rect	573	224	574	225
rect	573	225	574	226
rect	573	226	574	227
rect	573	227	574	228
rect	573	228	574	229
rect	573	229	574	230
rect	573	230	574	231
rect	573	231	574	232
rect	573	232	574	233
rect	573	233	574	234
rect	573	234	574	235
rect	573	235	574	236
rect	573	236	574	237
rect	573	237	574	238
rect	573	238	574	239
rect	573	239	574	240
rect	573	240	574	241
rect	573	241	574	242
rect	573	242	574	243
rect	573	243	574	244
rect	573	244	574	245
rect	573	245	574	246
rect	573	246	574	247
rect	573	247	574	248
rect	573	248	574	249
rect	573	249	574	250
rect	573	250	574	251
rect	573	251	574	252
rect	573	252	574	253
rect	573	253	574	254
rect	573	254	574	255
rect	573	255	574	256
rect	573	256	574	257
rect	573	257	574	258
rect	573	258	574	259
rect	573	259	574	260
rect	573	260	574	261
rect	573	261	574	262
rect	573	262	574	263
rect	573	263	574	264
rect	573	264	574	265
rect	573	265	574	266
rect	573	266	574	267
rect	573	267	574	268
rect	573	268	574	269
rect	573	269	574	270
rect	574	0	575	1
rect	574	1	575	2
rect	574	2	575	3
rect	574	3	575	4
rect	574	4	575	5
rect	574	5	575	6
rect	574	6	575	7
rect	574	7	575	8
rect	574	8	575	9
rect	574	9	575	10
rect	574	10	575	11
rect	574	11	575	12
rect	574	12	575	13
rect	574	13	575	14
rect	574	14	575	15
rect	574	15	575	16
rect	574	16	575	17
rect	574	17	575	18
rect	574	18	575	19
rect	574	19	575	20
rect	574	20	575	21
rect	574	21	575	22
rect	574	22	575	23
rect	574	23	575	24
rect	574	24	575	25
rect	574	25	575	26
rect	574	26	575	27
rect	574	27	575	28
rect	574	28	575	29
rect	574	29	575	30
rect	574	30	575	31
rect	574	31	575	32
rect	574	32	575	33
rect	574	33	575	34
rect	574	34	575	35
rect	574	35	575	36
rect	574	36	575	37
rect	574	37	575	38
rect	574	38	575	39
rect	574	39	575	40
rect	574	40	575	41
rect	574	41	575	42
rect	574	42	575	43
rect	574	43	575	44
rect	574	44	575	45
rect	574	45	575	46
rect	574	46	575	47
rect	574	47	575	48
rect	574	48	575	49
rect	574	49	575	50
rect	574	50	575	51
rect	574	51	575	52
rect	574	52	575	53
rect	574	53	575	54
rect	574	54	575	55
rect	574	55	575	56
rect	574	56	575	57
rect	574	57	575	58
rect	574	58	575	59
rect	574	59	575	60
rect	574	60	575	61
rect	574	61	575	62
rect	574	62	575	63
rect	574	63	575	64
rect	574	64	575	65
rect	574	65	575	66
rect	574	66	575	67
rect	574	67	575	68
rect	574	68	575	69
rect	574	69	575	70
rect	574	70	575	71
rect	574	71	575	72
rect	574	72	575	73
rect	574	73	575	74
rect	574	74	575	75
rect	574	75	575	76
rect	574	76	575	77
rect	574	77	575	78
rect	574	78	575	79
rect	574	79	575	80
rect	574	80	575	81
rect	574	81	575	82
rect	574	82	575	83
rect	574	83	575	84
rect	574	84	575	85
rect	574	85	575	86
rect	574	86	575	87
rect	574	87	575	88
rect	574	88	575	89
rect	574	89	575	90
rect	574	90	575	91
rect	574	91	575	92
rect	574	92	575	93
rect	574	93	575	94
rect	574	94	575	95
rect	574	95	575	96
rect	574	96	575	97
rect	574	97	575	98
rect	574	98	575	99
rect	574	99	575	100
rect	574	100	575	101
rect	574	101	575	102
rect	574	102	575	103
rect	574	103	575	104
rect	574	104	575	105
rect	574	105	575	106
rect	574	106	575	107
rect	574	107	575	108
rect	574	108	575	109
rect	574	109	575	110
rect	574	110	575	111
rect	574	111	575	112
rect	574	112	575	113
rect	574	113	575	114
rect	574	114	575	115
rect	574	115	575	116
rect	574	116	575	117
rect	574	117	575	118
rect	574	118	575	119
rect	574	119	575	120
rect	574	120	575	121
rect	574	121	575	122
rect	574	122	575	123
rect	574	123	575	124
rect	574	124	575	125
rect	574	125	575	126
rect	574	126	575	127
rect	574	127	575	128
rect	574	128	575	129
rect	574	129	575	130
rect	574	130	575	131
rect	574	131	575	132
rect	574	132	575	133
rect	574	133	575	134
rect	574	134	575	135
rect	574	135	575	136
rect	574	136	575	137
rect	574	137	575	138
rect	574	138	575	139
rect	574	139	575	140
rect	574	140	575	141
rect	574	141	575	142
rect	574	142	575	143
rect	574	143	575	144
rect	574	144	575	145
rect	574	145	575	146
rect	574	146	575	147
rect	574	147	575	148
rect	574	148	575	149
rect	574	149	575	150
rect	574	150	575	151
rect	574	151	575	152
rect	574	152	575	153
rect	574	153	575	154
rect	574	154	575	155
rect	574	155	575	156
rect	574	156	575	157
rect	574	157	575	158
rect	574	158	575	159
rect	574	159	575	160
rect	574	160	575	161
rect	574	161	575	162
rect	574	162	575	163
rect	574	163	575	164
rect	574	164	575	165
rect	574	165	575	166
rect	574	166	575	167
rect	574	167	575	168
rect	574	168	575	169
rect	574	169	575	170
rect	574	170	575	171
rect	574	171	575	172
rect	574	172	575	173
rect	574	173	575	174
rect	574	174	575	175
rect	574	175	575	176
rect	574	176	575	177
rect	574	177	575	178
rect	574	178	575	179
rect	574	179	575	180
rect	574	180	575	181
rect	574	181	575	182
rect	574	182	575	183
rect	574	183	575	184
rect	574	184	575	185
rect	574	185	575	186
rect	574	186	575	187
rect	574	187	575	188
rect	574	188	575	189
rect	574	189	575	190
rect	574	190	575	191
rect	574	191	575	192
rect	574	192	575	193
rect	574	193	575	194
rect	574	194	575	195
rect	574	195	575	196
rect	574	196	575	197
rect	574	197	575	198
rect	574	198	575	199
rect	574	199	575	200
rect	574	200	575	201
rect	574	201	575	202
rect	574	202	575	203
rect	574	203	575	204
rect	574	204	575	205
rect	574	205	575	206
rect	574	206	575	207
rect	574	207	575	208
rect	574	208	575	209
rect	574	209	575	210
rect	574	210	575	211
rect	574	211	575	212
rect	574	212	575	213
rect	574	213	575	214
rect	574	214	575	215
rect	574	215	575	216
rect	574	216	575	217
rect	574	217	575	218
rect	574	218	575	219
rect	574	219	575	220
rect	574	220	575	221
rect	574	221	575	222
rect	574	222	575	223
rect	574	223	575	224
rect	574	224	575	225
rect	574	225	575	226
rect	574	226	575	227
rect	574	227	575	228
rect	574	228	575	229
rect	574	229	575	230
rect	574	230	575	231
rect	574	231	575	232
rect	574	232	575	233
rect	574	233	575	234
rect	574	234	575	235
rect	574	235	575	236
rect	574	236	575	237
rect	574	237	575	238
rect	574	238	575	239
rect	574	239	575	240
rect	574	240	575	241
rect	574	241	575	242
rect	574	242	575	243
rect	574	243	575	244
rect	574	244	575	245
rect	574	245	575	246
rect	574	246	575	247
rect	574	247	575	248
rect	574	248	575	249
rect	574	249	575	250
rect	574	250	575	251
rect	574	251	575	252
rect	574	252	575	253
rect	574	253	575	254
rect	574	254	575	255
rect	574	255	575	256
rect	574	256	575	257
rect	574	257	575	258
rect	574	258	575	259
rect	574	259	575	260
rect	574	260	575	261
rect	574	261	575	262
rect	574	262	575	263
rect	574	263	575	264
rect	574	264	575	265
rect	574	265	575	266
rect	574	266	575	267
rect	574	267	575	268
rect	574	268	575	269
rect	574	269	575	270
rect	575	0	576	1
rect	575	1	576	2
rect	575	2	576	3
rect	575	3	576	4
rect	575	4	576	5
rect	575	5	576	6
rect	575	6	576	7
rect	575	7	576	8
rect	575	8	576	9
rect	575	9	576	10
rect	575	10	576	11
rect	575	11	576	12
rect	575	12	576	13
rect	575	13	576	14
rect	575	14	576	15
rect	575	15	576	16
rect	575	16	576	17
rect	575	17	576	18
rect	575	18	576	19
rect	575	19	576	20
rect	575	20	576	21
rect	575	21	576	22
rect	575	22	576	23
rect	575	23	576	24
rect	575	24	576	25
rect	575	25	576	26
rect	575	26	576	27
rect	575	27	576	28
rect	575	28	576	29
rect	575	29	576	30
rect	575	30	576	31
rect	575	31	576	32
rect	575	32	576	33
rect	575	33	576	34
rect	575	34	576	35
rect	575	35	576	36
rect	575	36	576	37
rect	575	37	576	38
rect	575	38	576	39
rect	575	39	576	40
rect	575	40	576	41
rect	575	41	576	42
rect	575	42	576	43
rect	575	43	576	44
rect	575	44	576	45
rect	575	45	576	46
rect	575	46	576	47
rect	575	47	576	48
rect	575	48	576	49
rect	575	49	576	50
rect	575	50	576	51
rect	575	51	576	52
rect	575	52	576	53
rect	575	53	576	54
rect	575	54	576	55
rect	575	55	576	56
rect	575	56	576	57
rect	575	57	576	58
rect	575	58	576	59
rect	575	59	576	60
rect	575	60	576	61
rect	575	61	576	62
rect	575	62	576	63
rect	575	63	576	64
rect	575	64	576	65
rect	575	65	576	66
rect	575	66	576	67
rect	575	67	576	68
rect	575	68	576	69
rect	575	69	576	70
rect	575	70	576	71
rect	575	71	576	72
rect	575	72	576	73
rect	575	73	576	74
rect	575	74	576	75
rect	575	75	576	76
rect	575	76	576	77
rect	575	77	576	78
rect	575	78	576	79
rect	575	79	576	80
rect	575	80	576	81
rect	575	81	576	82
rect	575	82	576	83
rect	575	83	576	84
rect	575	84	576	85
rect	575	85	576	86
rect	575	86	576	87
rect	575	87	576	88
rect	575	88	576	89
rect	575	89	576	90
rect	575	90	576	91
rect	575	91	576	92
rect	575	92	576	93
rect	575	93	576	94
rect	575	94	576	95
rect	575	95	576	96
rect	575	96	576	97
rect	575	97	576	98
rect	575	98	576	99
rect	575	99	576	100
rect	575	100	576	101
rect	575	101	576	102
rect	575	102	576	103
rect	575	103	576	104
rect	575	104	576	105
rect	575	105	576	106
rect	575	106	576	107
rect	575	107	576	108
rect	575	108	576	109
rect	575	109	576	110
rect	575	110	576	111
rect	575	111	576	112
rect	575	112	576	113
rect	575	113	576	114
rect	575	114	576	115
rect	575	115	576	116
rect	575	116	576	117
rect	575	117	576	118
rect	575	118	576	119
rect	575	119	576	120
rect	575	120	576	121
rect	575	121	576	122
rect	575	122	576	123
rect	575	123	576	124
rect	575	124	576	125
rect	575	125	576	126
rect	575	126	576	127
rect	575	127	576	128
rect	575	128	576	129
rect	575	129	576	130
rect	575	130	576	131
rect	575	131	576	132
rect	575	132	576	133
rect	575	133	576	134
rect	575	134	576	135
rect	575	135	576	136
rect	575	136	576	137
rect	575	137	576	138
rect	575	138	576	139
rect	575	139	576	140
rect	575	140	576	141
rect	575	141	576	142
rect	575	142	576	143
rect	575	143	576	144
rect	575	144	576	145
rect	575	145	576	146
rect	575	146	576	147
rect	575	147	576	148
rect	575	148	576	149
rect	575	149	576	150
rect	575	150	576	151
rect	575	151	576	152
rect	575	152	576	153
rect	575	153	576	154
rect	575	154	576	155
rect	575	155	576	156
rect	575	156	576	157
rect	575	157	576	158
rect	575	158	576	159
rect	575	159	576	160
rect	575	160	576	161
rect	575	161	576	162
rect	575	162	576	163
rect	575	163	576	164
rect	575	164	576	165
rect	575	165	576	166
rect	575	166	576	167
rect	575	167	576	168
rect	575	168	576	169
rect	575	169	576	170
rect	575	170	576	171
rect	575	171	576	172
rect	575	172	576	173
rect	575	173	576	174
rect	575	174	576	175
rect	575	175	576	176
rect	575	176	576	177
rect	575	177	576	178
rect	575	178	576	179
rect	575	179	576	180
rect	575	180	576	181
rect	575	181	576	182
rect	575	182	576	183
rect	575	183	576	184
rect	575	184	576	185
rect	575	185	576	186
rect	575	186	576	187
rect	575	187	576	188
rect	575	188	576	189
rect	575	189	576	190
rect	575	190	576	191
rect	575	191	576	192
rect	575	192	576	193
rect	575	193	576	194
rect	575	194	576	195
rect	575	195	576	196
rect	575	196	576	197
rect	575	197	576	198
rect	575	198	576	199
rect	575	199	576	200
rect	575	200	576	201
rect	575	201	576	202
rect	575	202	576	203
rect	575	203	576	204
rect	575	204	576	205
rect	575	205	576	206
rect	575	206	576	207
rect	575	207	576	208
rect	575	208	576	209
rect	575	209	576	210
rect	575	210	576	211
rect	575	211	576	212
rect	575	212	576	213
rect	575	213	576	214
rect	575	214	576	215
rect	575	215	576	216
rect	575	216	576	217
rect	575	217	576	218
rect	575	218	576	219
rect	575	219	576	220
rect	575	220	576	221
rect	575	221	576	222
rect	575	222	576	223
rect	575	223	576	224
rect	575	224	576	225
rect	575	225	576	226
rect	575	226	576	227
rect	575	227	576	228
rect	575	228	576	229
rect	575	229	576	230
rect	575	230	576	231
rect	575	231	576	232
rect	575	232	576	233
rect	575	233	576	234
rect	575	234	576	235
rect	575	235	576	236
rect	575	236	576	237
rect	575	237	576	238
rect	575	238	576	239
rect	575	239	576	240
rect	575	240	576	241
rect	575	241	576	242
rect	575	242	576	243
rect	575	243	576	244
rect	575	244	576	245
rect	575	245	576	246
rect	575	246	576	247
rect	575	247	576	248
rect	575	248	576	249
rect	575	249	576	250
rect	575	250	576	251
rect	575	251	576	252
rect	575	252	576	253
rect	575	253	576	254
rect	575	254	576	255
rect	575	255	576	256
rect	575	256	576	257
rect	575	257	576	258
rect	575	258	576	259
rect	575	259	576	260
rect	575	260	576	261
rect	575	261	576	262
rect	575	262	576	263
rect	575	263	576	264
rect	575	264	576	265
rect	575	265	576	266
rect	575	266	576	267
rect	575	267	576	268
rect	575	268	576	269
rect	575	269	576	270
rect	597	0	598	1
rect	597	1	598	2
rect	597	2	598	3
rect	597	3	598	4
rect	597	4	598	5
rect	597	5	598	6
rect	597	6	598	7
rect	597	7	598	8
rect	597	8	598	9
rect	597	9	598	10
rect	597	10	598	11
rect	597	11	598	12
rect	597	12	598	13
rect	597	13	598	14
rect	597	14	598	15
rect	597	15	598	16
rect	597	16	598	17
rect	597	17	598	18
rect	597	18	598	19
rect	597	19	598	20
rect	597	20	598	21
rect	597	21	598	22
rect	597	22	598	23
rect	597	23	598	24
rect	597	24	598	25
rect	597	25	598	26
rect	597	26	598	27
rect	597	27	598	28
rect	597	28	598	29
rect	597	29	598	30
rect	597	30	598	31
rect	597	31	598	32
rect	597	32	598	33
rect	597	33	598	34
rect	597	34	598	35
rect	597	35	598	36
rect	597	36	598	37
rect	597	37	598	38
rect	597	38	598	39
rect	597	39	598	40
rect	597	40	598	41
rect	597	41	598	42
rect	597	42	598	43
rect	597	43	598	44
rect	597	44	598	45
rect	597	45	598	46
rect	597	46	598	47
rect	597	47	598	48
rect	597	48	598	49
rect	597	49	598	50
rect	597	50	598	51
rect	597	51	598	52
rect	597	52	598	53
rect	597	53	598	54
rect	597	54	598	55
rect	597	55	598	56
rect	597	56	598	57
rect	597	57	598	58
rect	597	58	598	59
rect	597	59	598	60
rect	597	60	598	61
rect	597	61	598	62
rect	597	62	598	63
rect	597	63	598	64
rect	597	64	598	65
rect	597	65	598	66
rect	597	66	598	67
rect	597	67	598	68
rect	597	68	598	69
rect	597	69	598	70
rect	597	70	598	71
rect	597	71	598	72
rect	597	72	598	73
rect	597	73	598	74
rect	597	74	598	75
rect	597	75	598	76
rect	597	76	598	77
rect	597	77	598	78
rect	597	78	598	79
rect	597	79	598	80
rect	597	80	598	81
rect	597	81	598	82
rect	597	82	598	83
rect	597	83	598	84
rect	597	84	598	85
rect	597	85	598	86
rect	597	86	598	87
rect	597	87	598	88
rect	597	88	598	89
rect	597	89	598	90
rect	597	90	598	91
rect	597	91	598	92
rect	597	92	598	93
rect	597	93	598	94
rect	597	94	598	95
rect	597	95	598	96
rect	597	96	598	97
rect	597	97	598	98
rect	597	98	598	99
rect	597	99	598	100
rect	597	100	598	101
rect	597	101	598	102
rect	597	102	598	103
rect	597	103	598	104
rect	597	104	598	105
rect	597	105	598	106
rect	597	106	598	107
rect	597	107	598	108
rect	597	108	598	109
rect	597	109	598	110
rect	597	110	598	111
rect	597	111	598	112
rect	597	112	598	113
rect	597	113	598	114
rect	597	114	598	115
rect	597	115	598	116
rect	597	116	598	117
rect	597	117	598	118
rect	597	118	598	119
rect	597	119	598	120
rect	597	120	598	121
rect	597	121	598	122
rect	597	122	598	123
rect	597	123	598	124
rect	597	124	598	125
rect	597	125	598	126
rect	597	126	598	127
rect	597	127	598	128
rect	597	128	598	129
rect	597	129	598	130
rect	597	130	598	131
rect	597	131	598	132
rect	597	132	598	133
rect	597	133	598	134
rect	597	134	598	135
rect	597	135	598	136
rect	597	136	598	137
rect	597	137	598	138
rect	597	138	598	139
rect	597	139	598	140
rect	597	140	598	141
rect	597	141	598	142
rect	597	142	598	143
rect	597	143	598	144
rect	597	144	598	145
rect	597	145	598	146
rect	597	146	598	147
rect	597	147	598	148
rect	597	148	598	149
rect	597	149	598	150
rect	597	150	598	151
rect	597	151	598	152
rect	597	152	598	153
rect	597	153	598	154
rect	597	154	598	155
rect	597	155	598	156
rect	597	156	598	157
rect	597	157	598	158
rect	597	158	598	159
rect	597	159	598	160
rect	597	160	598	161
rect	597	161	598	162
rect	597	162	598	163
rect	597	163	598	164
rect	597	164	598	165
rect	597	165	598	166
rect	597	166	598	167
rect	597	167	598	168
rect	597	168	598	169
rect	597	169	598	170
rect	597	170	598	171
rect	597	171	598	172
rect	597	172	598	173
rect	597	173	598	174
rect	597	174	598	175
rect	597	175	598	176
rect	597	176	598	177
rect	597	177	598	178
rect	597	178	598	179
rect	597	179	598	180
rect	597	180	598	181
rect	597	181	598	182
rect	597	182	598	183
rect	597	183	598	184
rect	597	184	598	185
rect	597	185	598	186
rect	597	186	598	187
rect	597	187	598	188
rect	597	188	598	189
rect	597	189	598	190
rect	597	190	598	191
rect	597	191	598	192
rect	597	192	598	193
rect	597	193	598	194
rect	597	194	598	195
rect	597	195	598	196
rect	597	196	598	197
rect	597	197	598	198
rect	597	198	598	199
rect	597	199	598	200
rect	597	200	598	201
rect	597	201	598	202
rect	597	202	598	203
rect	597	203	598	204
rect	597	204	598	205
rect	597	205	598	206
rect	597	206	598	207
rect	597	207	598	208
rect	597	208	598	209
rect	597	209	598	210
rect	597	210	598	211
rect	597	211	598	212
rect	597	212	598	213
rect	597	213	598	214
rect	597	214	598	215
rect	597	215	598	216
rect	597	216	598	217
rect	597	217	598	218
rect	597	218	598	219
rect	597	219	598	220
rect	597	220	598	221
rect	597	221	598	222
rect	597	222	598	223
rect	597	223	598	224
rect	597	224	598	225
rect	597	225	598	226
rect	597	226	598	227
rect	597	227	598	228
rect	597	228	598	229
rect	597	229	598	230
rect	597	230	598	231
rect	597	231	598	232
rect	597	232	598	233
rect	597	233	598	234
rect	597	234	598	235
rect	597	235	598	236
rect	597	236	598	237
rect	597	237	598	238
rect	597	238	598	239
rect	597	239	598	240
rect	597	240	598	241
rect	597	241	598	242
rect	597	242	598	243
rect	597	243	598	244
rect	597	244	598	245
rect	597	245	598	246
rect	597	246	598	247
rect	597	247	598	248
rect	597	248	598	249
rect	597	249	598	250
rect	597	250	598	251
rect	597	251	598	252
rect	598	0	599	1
rect	598	1	599	2
rect	598	2	599	3
rect	598	3	599	4
rect	598	4	599	5
rect	598	5	599	6
rect	598	6	599	7
rect	598	7	599	8
rect	598	8	599	9
rect	598	9	599	10
rect	598	10	599	11
rect	598	11	599	12
rect	598	12	599	13
rect	598	13	599	14
rect	598	14	599	15
rect	598	15	599	16
rect	598	16	599	17
rect	598	17	599	18
rect	598	18	599	19
rect	598	19	599	20
rect	598	20	599	21
rect	598	21	599	22
rect	598	22	599	23
rect	598	23	599	24
rect	598	24	599	25
rect	598	25	599	26
rect	598	26	599	27
rect	598	27	599	28
rect	598	28	599	29
rect	598	29	599	30
rect	598	30	599	31
rect	598	31	599	32
rect	598	32	599	33
rect	598	33	599	34
rect	598	34	599	35
rect	598	35	599	36
rect	598	36	599	37
rect	598	37	599	38
rect	598	38	599	39
rect	598	39	599	40
rect	598	40	599	41
rect	598	41	599	42
rect	598	42	599	43
rect	598	43	599	44
rect	598	44	599	45
rect	598	45	599	46
rect	598	46	599	47
rect	598	47	599	48
rect	598	48	599	49
rect	598	49	599	50
rect	598	50	599	51
rect	598	51	599	52
rect	598	52	599	53
rect	598	53	599	54
rect	598	54	599	55
rect	598	55	599	56
rect	598	56	599	57
rect	598	57	599	58
rect	598	58	599	59
rect	598	59	599	60
rect	598	60	599	61
rect	598	61	599	62
rect	598	62	599	63
rect	598	63	599	64
rect	598	64	599	65
rect	598	65	599	66
rect	598	66	599	67
rect	598	67	599	68
rect	598	68	599	69
rect	598	69	599	70
rect	598	70	599	71
rect	598	71	599	72
rect	598	72	599	73
rect	598	73	599	74
rect	598	74	599	75
rect	598	75	599	76
rect	598	76	599	77
rect	598	77	599	78
rect	598	78	599	79
rect	598	79	599	80
rect	598	80	599	81
rect	598	81	599	82
rect	598	82	599	83
rect	598	83	599	84
rect	598	84	599	85
rect	598	85	599	86
rect	598	86	599	87
rect	598	87	599	88
rect	598	88	599	89
rect	598	89	599	90
rect	598	90	599	91
rect	598	91	599	92
rect	598	92	599	93
rect	598	93	599	94
rect	598	94	599	95
rect	598	95	599	96
rect	598	96	599	97
rect	598	97	599	98
rect	598	98	599	99
rect	598	99	599	100
rect	598	100	599	101
rect	598	101	599	102
rect	598	102	599	103
rect	598	103	599	104
rect	598	104	599	105
rect	598	105	599	106
rect	598	106	599	107
rect	598	107	599	108
rect	598	108	599	109
rect	598	109	599	110
rect	598	110	599	111
rect	598	111	599	112
rect	598	112	599	113
rect	598	113	599	114
rect	598	114	599	115
rect	598	115	599	116
rect	598	116	599	117
rect	598	117	599	118
rect	598	118	599	119
rect	598	119	599	120
rect	598	120	599	121
rect	598	121	599	122
rect	598	122	599	123
rect	598	123	599	124
rect	598	124	599	125
rect	598	125	599	126
rect	598	126	599	127
rect	598	127	599	128
rect	598	128	599	129
rect	598	129	599	130
rect	598	130	599	131
rect	598	131	599	132
rect	598	132	599	133
rect	598	133	599	134
rect	598	134	599	135
rect	598	135	599	136
rect	598	136	599	137
rect	598	137	599	138
rect	598	138	599	139
rect	598	139	599	140
rect	598	140	599	141
rect	598	141	599	142
rect	598	142	599	143
rect	598	143	599	144
rect	598	144	599	145
rect	598	145	599	146
rect	598	146	599	147
rect	598	147	599	148
rect	598	148	599	149
rect	598	149	599	150
rect	598	150	599	151
rect	598	151	599	152
rect	598	152	599	153
rect	598	153	599	154
rect	598	154	599	155
rect	598	155	599	156
rect	598	156	599	157
rect	598	157	599	158
rect	598	158	599	159
rect	598	159	599	160
rect	598	160	599	161
rect	598	161	599	162
rect	598	162	599	163
rect	598	163	599	164
rect	598	164	599	165
rect	598	165	599	166
rect	598	166	599	167
rect	598	167	599	168
rect	598	168	599	169
rect	598	169	599	170
rect	598	170	599	171
rect	598	171	599	172
rect	598	172	599	173
rect	598	173	599	174
rect	598	174	599	175
rect	598	175	599	176
rect	598	176	599	177
rect	598	177	599	178
rect	598	178	599	179
rect	598	179	599	180
rect	598	180	599	181
rect	598	181	599	182
rect	598	182	599	183
rect	598	183	599	184
rect	598	184	599	185
rect	598	185	599	186
rect	598	186	599	187
rect	598	187	599	188
rect	598	188	599	189
rect	598	189	599	190
rect	598	190	599	191
rect	598	191	599	192
rect	598	192	599	193
rect	598	193	599	194
rect	598	194	599	195
rect	598	195	599	196
rect	598	196	599	197
rect	598	197	599	198
rect	598	198	599	199
rect	598	199	599	200
rect	598	200	599	201
rect	598	201	599	202
rect	598	202	599	203
rect	598	203	599	204
rect	598	204	599	205
rect	598	205	599	206
rect	598	206	599	207
rect	598	207	599	208
rect	598	208	599	209
rect	598	209	599	210
rect	598	210	599	211
rect	598	211	599	212
rect	598	212	599	213
rect	598	213	599	214
rect	598	214	599	215
rect	598	215	599	216
rect	598	216	599	217
rect	598	217	599	218
rect	598	218	599	219
rect	598	219	599	220
rect	598	220	599	221
rect	598	221	599	222
rect	598	222	599	223
rect	598	223	599	224
rect	598	224	599	225
rect	598	225	599	226
rect	598	226	599	227
rect	598	227	599	228
rect	598	228	599	229
rect	598	229	599	230
rect	598	230	599	231
rect	598	231	599	232
rect	598	232	599	233
rect	598	233	599	234
rect	598	234	599	235
rect	598	235	599	236
rect	598	236	599	237
rect	598	237	599	238
rect	598	238	599	239
rect	598	239	599	240
rect	598	240	599	241
rect	598	241	599	242
rect	598	242	599	243
rect	598	243	599	244
rect	598	244	599	245
rect	598	245	599	246
rect	598	246	599	247
rect	598	247	599	248
rect	598	248	599	249
rect	598	249	599	250
rect	598	250	599	251
rect	598	251	599	252
rect	599	0	600	1
rect	599	1	600	2
rect	599	2	600	3
rect	599	3	600	4
rect	599	4	600	5
rect	599	5	600	6
rect	599	6	600	7
rect	599	7	600	8
rect	599	8	600	9
rect	599	9	600	10
rect	599	10	600	11
rect	599	11	600	12
rect	599	12	600	13
rect	599	13	600	14
rect	599	14	600	15
rect	599	15	600	16
rect	599	16	600	17
rect	599	17	600	18
rect	599	18	600	19
rect	599	19	600	20
rect	599	20	600	21
rect	599	21	600	22
rect	599	22	600	23
rect	599	23	600	24
rect	599	24	600	25
rect	599	25	600	26
rect	599	26	600	27
rect	599	27	600	28
rect	599	28	600	29
rect	599	29	600	30
rect	599	30	600	31
rect	599	31	600	32
rect	599	32	600	33
rect	599	33	600	34
rect	599	34	600	35
rect	599	35	600	36
rect	599	36	600	37
rect	599	37	600	38
rect	599	38	600	39
rect	599	39	600	40
rect	599	40	600	41
rect	599	41	600	42
rect	599	42	600	43
rect	599	43	600	44
rect	599	44	600	45
rect	599	45	600	46
rect	599	46	600	47
rect	599	47	600	48
rect	599	48	600	49
rect	599	49	600	50
rect	599	50	600	51
rect	599	51	600	52
rect	599	52	600	53
rect	599	53	600	54
rect	599	54	600	55
rect	599	55	600	56
rect	599	56	600	57
rect	599	57	600	58
rect	599	58	600	59
rect	599	59	600	60
rect	599	60	600	61
rect	599	61	600	62
rect	599	62	600	63
rect	599	63	600	64
rect	599	64	600	65
rect	599	65	600	66
rect	599	66	600	67
rect	599	67	600	68
rect	599	68	600	69
rect	599	69	600	70
rect	599	70	600	71
rect	599	71	600	72
rect	599	72	600	73
rect	599	73	600	74
rect	599	74	600	75
rect	599	75	600	76
rect	599	76	600	77
rect	599	77	600	78
rect	599	78	600	79
rect	599	79	600	80
rect	599	80	600	81
rect	599	81	600	82
rect	599	82	600	83
rect	599	83	600	84
rect	599	84	600	85
rect	599	85	600	86
rect	599	86	600	87
rect	599	87	600	88
rect	599	88	600	89
rect	599	89	600	90
rect	599	90	600	91
rect	599	91	600	92
rect	599	92	600	93
rect	599	93	600	94
rect	599	94	600	95
rect	599	95	600	96
rect	599	96	600	97
rect	599	97	600	98
rect	599	98	600	99
rect	599	99	600	100
rect	599	100	600	101
rect	599	101	600	102
rect	599	102	600	103
rect	599	103	600	104
rect	599	104	600	105
rect	599	105	600	106
rect	599	106	600	107
rect	599	107	600	108
rect	599	108	600	109
rect	599	109	600	110
rect	599	110	600	111
rect	599	111	600	112
rect	599	112	600	113
rect	599	113	600	114
rect	599	114	600	115
rect	599	115	600	116
rect	599	116	600	117
rect	599	117	600	118
rect	599	118	600	119
rect	599	119	600	120
rect	599	120	600	121
rect	599	121	600	122
rect	599	122	600	123
rect	599	123	600	124
rect	599	124	600	125
rect	599	125	600	126
rect	599	126	600	127
rect	599	127	600	128
rect	599	128	600	129
rect	599	129	600	130
rect	599	130	600	131
rect	599	131	600	132
rect	599	132	600	133
rect	599	133	600	134
rect	599	134	600	135
rect	599	135	600	136
rect	599	136	600	137
rect	599	137	600	138
rect	599	138	600	139
rect	599	139	600	140
rect	599	140	600	141
rect	599	141	600	142
rect	599	142	600	143
rect	599	143	600	144
rect	599	144	600	145
rect	599	145	600	146
rect	599	146	600	147
rect	599	147	600	148
rect	599	148	600	149
rect	599	149	600	150
rect	599	150	600	151
rect	599	151	600	152
rect	599	152	600	153
rect	599	153	600	154
rect	599	154	600	155
rect	599	155	600	156
rect	599	156	600	157
rect	599	157	600	158
rect	599	158	600	159
rect	599	159	600	160
rect	599	160	600	161
rect	599	161	600	162
rect	599	162	600	163
rect	599	163	600	164
rect	599	164	600	165
rect	599	165	600	166
rect	599	166	600	167
rect	599	167	600	168
rect	599	168	600	169
rect	599	169	600	170
rect	599	170	600	171
rect	599	171	600	172
rect	599	172	600	173
rect	599	173	600	174
rect	599	174	600	175
rect	599	175	600	176
rect	599	176	600	177
rect	599	177	600	178
rect	599	178	600	179
rect	599	179	600	180
rect	599	180	600	181
rect	599	181	600	182
rect	599	182	600	183
rect	599	183	600	184
rect	599	184	600	185
rect	599	185	600	186
rect	599	186	600	187
rect	599	187	600	188
rect	599	188	600	189
rect	599	189	600	190
rect	599	190	600	191
rect	599	191	600	192
rect	599	192	600	193
rect	599	193	600	194
rect	599	194	600	195
rect	599	195	600	196
rect	599	196	600	197
rect	599	197	600	198
rect	599	198	600	199
rect	599	199	600	200
rect	599	200	600	201
rect	599	201	600	202
rect	599	202	600	203
rect	599	203	600	204
rect	599	204	600	205
rect	599	205	600	206
rect	599	206	600	207
rect	599	207	600	208
rect	599	208	600	209
rect	599	209	600	210
rect	599	210	600	211
rect	599	211	600	212
rect	599	212	600	213
rect	599	213	600	214
rect	599	214	600	215
rect	599	215	600	216
rect	599	216	600	217
rect	599	217	600	218
rect	599	218	600	219
rect	599	219	600	220
rect	599	220	600	221
rect	599	221	600	222
rect	599	222	600	223
rect	599	223	600	224
rect	599	224	600	225
rect	599	225	600	226
rect	599	226	600	227
rect	599	227	600	228
rect	599	228	600	229
rect	599	229	600	230
rect	599	230	600	231
rect	599	231	600	232
rect	599	232	600	233
rect	599	233	600	234
rect	599	234	600	235
rect	599	235	600	236
rect	599	236	600	237
rect	599	237	600	238
rect	599	238	600	239
rect	599	239	600	240
rect	599	240	600	241
rect	599	241	600	242
rect	599	242	600	243
rect	599	243	600	244
rect	599	244	600	245
rect	599	245	600	246
rect	599	246	600	247
rect	599	247	600	248
rect	599	248	600	249
rect	599	249	600	250
rect	599	250	600	251
rect	599	251	600	252
rect	600	0	601	1
rect	600	1	601	2
rect	600	2	601	3
rect	600	3	601	4
rect	600	4	601	5
rect	600	5	601	6
rect	600	6	601	7
rect	600	7	601	8
rect	600	8	601	9
rect	600	9	601	10
rect	600	10	601	11
rect	600	11	601	12
rect	600	12	601	13
rect	600	13	601	14
rect	600	14	601	15
rect	600	15	601	16
rect	600	16	601	17
rect	600	17	601	18
rect	600	18	601	19
rect	600	19	601	20
rect	600	20	601	21
rect	600	21	601	22
rect	600	22	601	23
rect	600	23	601	24
rect	600	24	601	25
rect	600	25	601	26
rect	600	26	601	27
rect	600	27	601	28
rect	600	28	601	29
rect	600	29	601	30
rect	600	30	601	31
rect	600	31	601	32
rect	600	32	601	33
rect	600	33	601	34
rect	600	34	601	35
rect	600	35	601	36
rect	600	36	601	37
rect	600	37	601	38
rect	600	38	601	39
rect	600	39	601	40
rect	600	40	601	41
rect	600	41	601	42
rect	600	42	601	43
rect	600	43	601	44
rect	600	44	601	45
rect	600	45	601	46
rect	600	46	601	47
rect	600	47	601	48
rect	600	48	601	49
rect	600	49	601	50
rect	600	50	601	51
rect	600	51	601	52
rect	600	52	601	53
rect	600	53	601	54
rect	600	54	601	55
rect	600	55	601	56
rect	600	56	601	57
rect	600	57	601	58
rect	600	58	601	59
rect	600	59	601	60
rect	600	60	601	61
rect	600	61	601	62
rect	600	62	601	63
rect	600	63	601	64
rect	600	64	601	65
rect	600	65	601	66
rect	600	66	601	67
rect	600	67	601	68
rect	600	68	601	69
rect	600	69	601	70
rect	600	70	601	71
rect	600	71	601	72
rect	600	72	601	73
rect	600	73	601	74
rect	600	74	601	75
rect	600	75	601	76
rect	600	76	601	77
rect	600	77	601	78
rect	600	78	601	79
rect	600	79	601	80
rect	600	80	601	81
rect	600	81	601	82
rect	600	82	601	83
rect	600	83	601	84
rect	600	84	601	85
rect	600	85	601	86
rect	600	86	601	87
rect	600	87	601	88
rect	600	88	601	89
rect	600	89	601	90
rect	600	90	601	91
rect	600	91	601	92
rect	600	92	601	93
rect	600	93	601	94
rect	600	94	601	95
rect	600	95	601	96
rect	600	96	601	97
rect	600	97	601	98
rect	600	98	601	99
rect	600	99	601	100
rect	600	100	601	101
rect	600	101	601	102
rect	600	102	601	103
rect	600	103	601	104
rect	600	104	601	105
rect	600	105	601	106
rect	600	106	601	107
rect	600	107	601	108
rect	600	108	601	109
rect	600	109	601	110
rect	600	110	601	111
rect	600	111	601	112
rect	600	112	601	113
rect	600	113	601	114
rect	600	114	601	115
rect	600	115	601	116
rect	600	116	601	117
rect	600	117	601	118
rect	600	118	601	119
rect	600	119	601	120
rect	600	120	601	121
rect	600	121	601	122
rect	600	122	601	123
rect	600	123	601	124
rect	600	124	601	125
rect	600	125	601	126
rect	600	126	601	127
rect	600	127	601	128
rect	600	128	601	129
rect	600	129	601	130
rect	600	130	601	131
rect	600	131	601	132
rect	600	132	601	133
rect	600	133	601	134
rect	600	134	601	135
rect	600	135	601	136
rect	600	136	601	137
rect	600	137	601	138
rect	600	138	601	139
rect	600	139	601	140
rect	600	140	601	141
rect	600	141	601	142
rect	600	142	601	143
rect	600	143	601	144
rect	600	144	601	145
rect	600	145	601	146
rect	600	146	601	147
rect	600	147	601	148
rect	600	148	601	149
rect	600	149	601	150
rect	600	150	601	151
rect	600	151	601	152
rect	600	152	601	153
rect	600	153	601	154
rect	600	154	601	155
rect	600	155	601	156
rect	600	156	601	157
rect	600	157	601	158
rect	600	158	601	159
rect	600	159	601	160
rect	600	160	601	161
rect	600	161	601	162
rect	600	162	601	163
rect	600	163	601	164
rect	600	164	601	165
rect	600	165	601	166
rect	600	166	601	167
rect	600	167	601	168
rect	600	168	601	169
rect	600	169	601	170
rect	600	170	601	171
rect	600	171	601	172
rect	600	172	601	173
rect	600	173	601	174
rect	600	174	601	175
rect	600	175	601	176
rect	600	176	601	177
rect	600	177	601	178
rect	600	178	601	179
rect	600	179	601	180
rect	600	180	601	181
rect	600	181	601	182
rect	600	182	601	183
rect	600	183	601	184
rect	600	184	601	185
rect	600	185	601	186
rect	600	186	601	187
rect	600	187	601	188
rect	600	188	601	189
rect	600	189	601	190
rect	600	190	601	191
rect	600	191	601	192
rect	600	192	601	193
rect	600	193	601	194
rect	600	194	601	195
rect	600	195	601	196
rect	600	196	601	197
rect	600	197	601	198
rect	600	198	601	199
rect	600	199	601	200
rect	600	200	601	201
rect	600	201	601	202
rect	600	202	601	203
rect	600	203	601	204
rect	600	204	601	205
rect	600	205	601	206
rect	600	206	601	207
rect	600	207	601	208
rect	600	208	601	209
rect	600	209	601	210
rect	600	210	601	211
rect	600	211	601	212
rect	600	212	601	213
rect	600	213	601	214
rect	600	214	601	215
rect	600	215	601	216
rect	600	216	601	217
rect	600	217	601	218
rect	600	218	601	219
rect	600	219	601	220
rect	600	220	601	221
rect	600	221	601	222
rect	600	222	601	223
rect	600	223	601	224
rect	600	224	601	225
rect	600	225	601	226
rect	600	226	601	227
rect	600	227	601	228
rect	600	228	601	229
rect	600	229	601	230
rect	600	230	601	231
rect	600	231	601	232
rect	600	232	601	233
rect	600	233	601	234
rect	600	234	601	235
rect	600	235	601	236
rect	600	236	601	237
rect	600	237	601	238
rect	600	238	601	239
rect	600	239	601	240
rect	600	240	601	241
rect	600	241	601	242
rect	600	242	601	243
rect	600	243	601	244
rect	600	244	601	245
rect	600	245	601	246
rect	600	246	601	247
rect	600	247	601	248
rect	600	248	601	249
rect	600	249	601	250
rect	600	250	601	251
rect	600	251	601	252
rect	601	0	602	1
rect	601	1	602	2
rect	601	2	602	3
rect	601	3	602	4
rect	601	4	602	5
rect	601	5	602	6
rect	601	6	602	7
rect	601	7	602	8
rect	601	8	602	9
rect	601	9	602	10
rect	601	10	602	11
rect	601	11	602	12
rect	601	12	602	13
rect	601	13	602	14
rect	601	14	602	15
rect	601	15	602	16
rect	601	16	602	17
rect	601	17	602	18
rect	601	18	602	19
rect	601	19	602	20
rect	601	20	602	21
rect	601	21	602	22
rect	601	22	602	23
rect	601	23	602	24
rect	601	24	602	25
rect	601	25	602	26
rect	601	26	602	27
rect	601	27	602	28
rect	601	28	602	29
rect	601	29	602	30
rect	601	30	602	31
rect	601	31	602	32
rect	601	32	602	33
rect	601	33	602	34
rect	601	34	602	35
rect	601	35	602	36
rect	601	36	602	37
rect	601	37	602	38
rect	601	38	602	39
rect	601	39	602	40
rect	601	40	602	41
rect	601	41	602	42
rect	601	42	602	43
rect	601	43	602	44
rect	601	44	602	45
rect	601	45	602	46
rect	601	46	602	47
rect	601	47	602	48
rect	601	48	602	49
rect	601	49	602	50
rect	601	50	602	51
rect	601	51	602	52
rect	601	52	602	53
rect	601	53	602	54
rect	601	54	602	55
rect	601	55	602	56
rect	601	56	602	57
rect	601	57	602	58
rect	601	58	602	59
rect	601	59	602	60
rect	601	60	602	61
rect	601	61	602	62
rect	601	62	602	63
rect	601	63	602	64
rect	601	64	602	65
rect	601	65	602	66
rect	601	66	602	67
rect	601	67	602	68
rect	601	68	602	69
rect	601	69	602	70
rect	601	70	602	71
rect	601	71	602	72
rect	601	72	602	73
rect	601	73	602	74
rect	601	74	602	75
rect	601	75	602	76
rect	601	76	602	77
rect	601	77	602	78
rect	601	78	602	79
rect	601	79	602	80
rect	601	80	602	81
rect	601	81	602	82
rect	601	82	602	83
rect	601	83	602	84
rect	601	84	602	85
rect	601	85	602	86
rect	601	86	602	87
rect	601	87	602	88
rect	601	88	602	89
rect	601	89	602	90
rect	601	90	602	91
rect	601	91	602	92
rect	601	92	602	93
rect	601	93	602	94
rect	601	94	602	95
rect	601	95	602	96
rect	601	96	602	97
rect	601	97	602	98
rect	601	98	602	99
rect	601	99	602	100
rect	601	100	602	101
rect	601	101	602	102
rect	601	102	602	103
rect	601	103	602	104
rect	601	104	602	105
rect	601	105	602	106
rect	601	106	602	107
rect	601	107	602	108
rect	601	108	602	109
rect	601	109	602	110
rect	601	110	602	111
rect	601	111	602	112
rect	601	112	602	113
rect	601	113	602	114
rect	601	114	602	115
rect	601	115	602	116
rect	601	116	602	117
rect	601	117	602	118
rect	601	118	602	119
rect	601	119	602	120
rect	601	120	602	121
rect	601	121	602	122
rect	601	122	602	123
rect	601	123	602	124
rect	601	124	602	125
rect	601	125	602	126
rect	601	126	602	127
rect	601	127	602	128
rect	601	128	602	129
rect	601	129	602	130
rect	601	130	602	131
rect	601	131	602	132
rect	601	132	602	133
rect	601	133	602	134
rect	601	134	602	135
rect	601	135	602	136
rect	601	136	602	137
rect	601	137	602	138
rect	601	138	602	139
rect	601	139	602	140
rect	601	140	602	141
rect	601	141	602	142
rect	601	142	602	143
rect	601	143	602	144
rect	601	144	602	145
rect	601	145	602	146
rect	601	146	602	147
rect	601	147	602	148
rect	601	148	602	149
rect	601	149	602	150
rect	601	150	602	151
rect	601	151	602	152
rect	601	152	602	153
rect	601	153	602	154
rect	601	154	602	155
rect	601	155	602	156
rect	601	156	602	157
rect	601	157	602	158
rect	601	158	602	159
rect	601	159	602	160
rect	601	160	602	161
rect	601	161	602	162
rect	601	162	602	163
rect	601	163	602	164
rect	601	164	602	165
rect	601	165	602	166
rect	601	166	602	167
rect	601	167	602	168
rect	601	168	602	169
rect	601	169	602	170
rect	601	170	602	171
rect	601	171	602	172
rect	601	172	602	173
rect	601	173	602	174
rect	601	174	602	175
rect	601	175	602	176
rect	601	176	602	177
rect	601	177	602	178
rect	601	178	602	179
rect	601	179	602	180
rect	601	180	602	181
rect	601	181	602	182
rect	601	182	602	183
rect	601	183	602	184
rect	601	184	602	185
rect	601	185	602	186
rect	601	186	602	187
rect	601	187	602	188
rect	601	188	602	189
rect	601	189	602	190
rect	601	190	602	191
rect	601	191	602	192
rect	601	192	602	193
rect	601	193	602	194
rect	601	194	602	195
rect	601	195	602	196
rect	601	196	602	197
rect	601	197	602	198
rect	601	198	602	199
rect	601	199	602	200
rect	601	200	602	201
rect	601	201	602	202
rect	601	202	602	203
rect	601	203	602	204
rect	601	204	602	205
rect	601	205	602	206
rect	601	206	602	207
rect	601	207	602	208
rect	601	208	602	209
rect	601	209	602	210
rect	601	210	602	211
rect	601	211	602	212
rect	601	212	602	213
rect	601	213	602	214
rect	601	214	602	215
rect	601	215	602	216
rect	601	216	602	217
rect	601	217	602	218
rect	601	218	602	219
rect	601	219	602	220
rect	601	220	602	221
rect	601	221	602	222
rect	601	222	602	223
rect	601	223	602	224
rect	601	224	602	225
rect	601	225	602	226
rect	601	226	602	227
rect	601	227	602	228
rect	601	228	602	229
rect	601	229	602	230
rect	601	230	602	231
rect	601	231	602	232
rect	601	232	602	233
rect	601	233	602	234
rect	601	234	602	235
rect	601	235	602	236
rect	601	236	602	237
rect	601	237	602	238
rect	601	238	602	239
rect	601	239	602	240
rect	601	240	602	241
rect	601	241	602	242
rect	601	242	602	243
rect	601	243	602	244
rect	601	244	602	245
rect	601	245	602	246
rect	601	246	602	247
rect	601	247	602	248
rect	601	248	602	249
rect	601	249	602	250
rect	601	250	602	251
rect	601	251	602	252
rect	602	0	603	1
rect	602	1	603	2
rect	602	2	603	3
rect	602	3	603	4
rect	602	4	603	5
rect	602	5	603	6
rect	602	6	603	7
rect	602	7	603	8
rect	602	8	603	9
rect	602	9	603	10
rect	602	10	603	11
rect	602	11	603	12
rect	602	12	603	13
rect	602	13	603	14
rect	602	14	603	15
rect	602	15	603	16
rect	602	16	603	17
rect	602	17	603	18
rect	602	18	603	19
rect	602	19	603	20
rect	602	20	603	21
rect	602	21	603	22
rect	602	22	603	23
rect	602	23	603	24
rect	602	24	603	25
rect	602	25	603	26
rect	602	26	603	27
rect	602	27	603	28
rect	602	28	603	29
rect	602	29	603	30
rect	602	30	603	31
rect	602	31	603	32
rect	602	32	603	33
rect	602	33	603	34
rect	602	34	603	35
rect	602	35	603	36
rect	602	36	603	37
rect	602	37	603	38
rect	602	38	603	39
rect	602	39	603	40
rect	602	40	603	41
rect	602	41	603	42
rect	602	42	603	43
rect	602	43	603	44
rect	602	44	603	45
rect	602	45	603	46
rect	602	46	603	47
rect	602	47	603	48
rect	602	48	603	49
rect	602	49	603	50
rect	602	50	603	51
rect	602	51	603	52
rect	602	52	603	53
rect	602	53	603	54
rect	602	54	603	55
rect	602	55	603	56
rect	602	56	603	57
rect	602	57	603	58
rect	602	58	603	59
rect	602	59	603	60
rect	602	60	603	61
rect	602	61	603	62
rect	602	62	603	63
rect	602	63	603	64
rect	602	64	603	65
rect	602	65	603	66
rect	602	66	603	67
rect	602	67	603	68
rect	602	68	603	69
rect	602	69	603	70
rect	602	70	603	71
rect	602	71	603	72
rect	602	72	603	73
rect	602	73	603	74
rect	602	74	603	75
rect	602	75	603	76
rect	602	76	603	77
rect	602	77	603	78
rect	602	78	603	79
rect	602	79	603	80
rect	602	80	603	81
rect	602	81	603	82
rect	602	82	603	83
rect	602	83	603	84
rect	602	84	603	85
rect	602	85	603	86
rect	602	86	603	87
rect	602	87	603	88
rect	602	88	603	89
rect	602	89	603	90
rect	602	90	603	91
rect	602	91	603	92
rect	602	92	603	93
rect	602	93	603	94
rect	602	94	603	95
rect	602	95	603	96
rect	602	96	603	97
rect	602	97	603	98
rect	602	98	603	99
rect	602	99	603	100
rect	602	100	603	101
rect	602	101	603	102
rect	602	102	603	103
rect	602	103	603	104
rect	602	104	603	105
rect	602	105	603	106
rect	602	106	603	107
rect	602	107	603	108
rect	602	108	603	109
rect	602	109	603	110
rect	602	110	603	111
rect	602	111	603	112
rect	602	112	603	113
rect	602	113	603	114
rect	602	114	603	115
rect	602	115	603	116
rect	602	116	603	117
rect	602	117	603	118
rect	602	118	603	119
rect	602	119	603	120
rect	602	120	603	121
rect	602	121	603	122
rect	602	122	603	123
rect	602	123	603	124
rect	602	124	603	125
rect	602	125	603	126
rect	602	126	603	127
rect	602	127	603	128
rect	602	128	603	129
rect	602	129	603	130
rect	602	130	603	131
rect	602	131	603	132
rect	602	132	603	133
rect	602	133	603	134
rect	602	134	603	135
rect	602	135	603	136
rect	602	136	603	137
rect	602	137	603	138
rect	602	138	603	139
rect	602	139	603	140
rect	602	140	603	141
rect	602	141	603	142
rect	602	142	603	143
rect	602	143	603	144
rect	602	144	603	145
rect	602	145	603	146
rect	602	146	603	147
rect	602	147	603	148
rect	602	148	603	149
rect	602	149	603	150
rect	602	150	603	151
rect	602	151	603	152
rect	602	152	603	153
rect	602	153	603	154
rect	602	154	603	155
rect	602	155	603	156
rect	602	156	603	157
rect	602	157	603	158
rect	602	158	603	159
rect	602	159	603	160
rect	602	160	603	161
rect	602	161	603	162
rect	602	162	603	163
rect	602	163	603	164
rect	602	164	603	165
rect	602	165	603	166
rect	602	166	603	167
rect	602	167	603	168
rect	602	168	603	169
rect	602	169	603	170
rect	602	170	603	171
rect	602	171	603	172
rect	602	172	603	173
rect	602	173	603	174
rect	602	174	603	175
rect	602	175	603	176
rect	602	176	603	177
rect	602	177	603	178
rect	602	178	603	179
rect	602	179	603	180
rect	602	180	603	181
rect	602	181	603	182
rect	602	182	603	183
rect	602	183	603	184
rect	602	184	603	185
rect	602	185	603	186
rect	602	186	603	187
rect	602	187	603	188
rect	602	188	603	189
rect	602	189	603	190
rect	602	190	603	191
rect	602	191	603	192
rect	602	192	603	193
rect	602	193	603	194
rect	602	194	603	195
rect	602	195	603	196
rect	602	196	603	197
rect	602	197	603	198
rect	602	198	603	199
rect	602	199	603	200
rect	602	200	603	201
rect	602	201	603	202
rect	602	202	603	203
rect	602	203	603	204
rect	602	204	603	205
rect	602	205	603	206
rect	602	206	603	207
rect	602	207	603	208
rect	602	208	603	209
rect	602	209	603	210
rect	602	210	603	211
rect	602	211	603	212
rect	602	212	603	213
rect	602	213	603	214
rect	602	214	603	215
rect	602	215	603	216
rect	602	216	603	217
rect	602	217	603	218
rect	602	218	603	219
rect	602	219	603	220
rect	602	220	603	221
rect	602	221	603	222
rect	602	222	603	223
rect	602	223	603	224
rect	602	224	603	225
rect	602	225	603	226
rect	602	226	603	227
rect	602	227	603	228
rect	602	228	603	229
rect	602	229	603	230
rect	602	230	603	231
rect	602	231	603	232
rect	602	232	603	233
rect	602	233	603	234
rect	602	234	603	235
rect	602	235	603	236
rect	602	236	603	237
rect	602	237	603	238
rect	602	238	603	239
rect	602	239	603	240
rect	602	240	603	241
rect	602	241	603	242
rect	602	242	603	243
rect	602	243	603	244
rect	602	244	603	245
rect	602	245	603	246
rect	602	246	603	247
rect	602	247	603	248
rect	602	248	603	249
rect	602	249	603	250
rect	602	250	603	251
rect	602	251	603	252
rect	612	0	613	1
rect	612	1	613	2
rect	612	2	613	3
rect	612	3	613	4
rect	612	4	613	5
rect	612	5	613	6
rect	612	6	613	7
rect	612	7	613	8
rect	612	8	613	9
rect	612	9	613	10
rect	612	10	613	11
rect	612	11	613	12
rect	612	12	613	13
rect	612	13	613	14
rect	612	14	613	15
rect	612	15	613	16
rect	612	16	613	17
rect	612	17	613	18
rect	612	18	613	19
rect	612	19	613	20
rect	612	20	613	21
rect	612	21	613	22
rect	612	22	613	23
rect	612	23	613	24
rect	612	24	613	25
rect	612	25	613	26
rect	612	26	613	27
rect	612	27	613	28
rect	612	28	613	29
rect	612	29	613	30
rect	612	30	613	31
rect	612	31	613	32
rect	612	32	613	33
rect	612	33	613	34
rect	612	34	613	35
rect	612	35	613	36
rect	612	36	613	37
rect	612	37	613	38
rect	612	38	613	39
rect	612	39	613	40
rect	612	40	613	41
rect	612	41	613	42
rect	612	42	613	43
rect	612	43	613	44
rect	612	44	613	45
rect	612	45	613	46
rect	612	46	613	47
rect	612	47	613	48
rect	612	48	613	49
rect	612	49	613	50
rect	612	50	613	51
rect	612	51	613	52
rect	612	52	613	53
rect	612	53	613	54
rect	612	54	613	55
rect	612	55	613	56
rect	612	56	613	57
rect	612	57	613	58
rect	612	58	613	59
rect	612	59	613	60
rect	612	60	613	61
rect	612	61	613	62
rect	612	62	613	63
rect	612	63	613	64
rect	612	64	613	65
rect	612	65	613	66
rect	612	66	613	67
rect	612	67	613	68
rect	612	68	613	69
rect	612	69	613	70
rect	612	70	613	71
rect	612	71	613	72
rect	612	72	613	73
rect	612	73	613	74
rect	612	74	613	75
rect	612	75	613	76
rect	612	76	613	77
rect	612	77	613	78
rect	612	78	613	79
rect	612	79	613	80
rect	612	80	613	81
rect	612	81	613	82
rect	612	82	613	83
rect	612	83	613	84
rect	612	84	613	85
rect	612	85	613	86
rect	612	86	613	87
rect	612	87	613	88
rect	612	88	613	89
rect	612	89	613	90
rect	612	90	613	91
rect	612	91	613	92
rect	612	92	613	93
rect	612	93	613	94
rect	612	94	613	95
rect	612	95	613	96
rect	612	96	613	97
rect	612	97	613	98
rect	612	98	613	99
rect	612	99	613	100
rect	612	100	613	101
rect	612	101	613	102
rect	612	102	613	103
rect	612	103	613	104
rect	612	104	613	105
rect	612	105	613	106
rect	612	106	613	107
rect	612	107	613	108
rect	612	108	613	109
rect	612	109	613	110
rect	612	110	613	111
rect	612	111	613	112
rect	612	112	613	113
rect	612	113	613	114
rect	612	114	613	115
rect	612	115	613	116
rect	612	116	613	117
rect	612	117	613	118
rect	612	118	613	119
rect	612	119	613	120
rect	612	120	613	121
rect	612	121	613	122
rect	612	122	613	123
rect	612	123	613	124
rect	612	124	613	125
rect	612	125	613	126
rect	612	126	613	127
rect	612	127	613	128
rect	612	128	613	129
rect	612	129	613	130
rect	612	130	613	131
rect	612	131	613	132
rect	612	132	613	133
rect	612	133	613	134
rect	612	134	613	135
rect	612	135	613	136
rect	612	136	613	137
rect	612	137	613	138
rect	612	138	613	139
rect	612	139	613	140
rect	612	140	613	141
rect	612	141	613	142
rect	612	142	613	143
rect	612	143	613	144
rect	612	144	613	145
rect	612	145	613	146
rect	612	146	613	147
rect	612	147	613	148
rect	612	148	613	149
rect	612	149	613	150
rect	612	150	613	151
rect	612	151	613	152
rect	612	152	613	153
rect	612	153	613	154
rect	612	154	613	155
rect	612	155	613	156
rect	612	156	613	157
rect	612	157	613	158
rect	612	158	613	159
rect	612	159	613	160
rect	612	160	613	161
rect	612	161	613	162
rect	612	162	613	163
rect	612	163	613	164
rect	612	164	613	165
rect	612	165	613	166
rect	612	166	613	167
rect	612	167	613	168
rect	612	168	613	169
rect	612	169	613	170
rect	612	170	613	171
rect	612	171	613	172
rect	612	172	613	173
rect	612	173	613	174
rect	612	174	613	175
rect	612	175	613	176
rect	612	176	613	177
rect	612	177	613	178
rect	612	178	613	179
rect	612	179	613	180
rect	612	180	613	181
rect	612	181	613	182
rect	612	182	613	183
rect	612	183	613	184
rect	612	184	613	185
rect	612	185	613	186
rect	612	186	613	187
rect	612	187	613	188
rect	612	188	613	189
rect	612	189	613	190
rect	612	190	613	191
rect	612	191	613	192
rect	612	192	613	193
rect	612	193	613	194
rect	612	194	613	195
rect	612	195	613	196
rect	612	196	613	197
rect	612	197	613	198
rect	612	198	613	199
rect	612	199	613	200
rect	612	200	613	201
rect	612	201	613	202
rect	612	202	613	203
rect	612	203	613	204
rect	612	204	613	205
rect	612	205	613	206
rect	612	206	613	207
rect	612	207	613	208
rect	612	208	613	209
rect	612	209	613	210
rect	612	210	613	211
rect	612	211	613	212
rect	612	212	613	213
rect	612	213	613	214
rect	612	214	613	215
rect	612	215	613	216
rect	612	216	613	217
rect	612	217	613	218
rect	612	218	613	219
rect	612	219	613	220
rect	612	220	613	221
rect	612	221	613	222
rect	612	222	613	223
rect	612	223	613	224
rect	612	224	613	225
rect	612	225	613	226
rect	612	226	613	227
rect	612	227	613	228
rect	612	228	613	229
rect	612	229	613	230
rect	612	230	613	231
rect	612	231	613	232
rect	612	232	613	233
rect	612	233	613	234
rect	612	234	613	235
rect	612	235	613	236
rect	612	236	613	237
rect	612	237	613	238
rect	612	238	613	239
rect	612	239	613	240
rect	613	0	614	1
rect	613	1	614	2
rect	613	2	614	3
rect	613	3	614	4
rect	613	4	614	5
rect	613	5	614	6
rect	613	6	614	7
rect	613	7	614	8
rect	613	8	614	9
rect	613	9	614	10
rect	613	10	614	11
rect	613	11	614	12
rect	613	12	614	13
rect	613	13	614	14
rect	613	14	614	15
rect	613	15	614	16
rect	613	16	614	17
rect	613	17	614	18
rect	613	18	614	19
rect	613	19	614	20
rect	613	20	614	21
rect	613	21	614	22
rect	613	22	614	23
rect	613	23	614	24
rect	613	24	614	25
rect	613	25	614	26
rect	613	26	614	27
rect	613	27	614	28
rect	613	28	614	29
rect	613	29	614	30
rect	613	30	614	31
rect	613	31	614	32
rect	613	32	614	33
rect	613	33	614	34
rect	613	34	614	35
rect	613	35	614	36
rect	613	36	614	37
rect	613	37	614	38
rect	613	38	614	39
rect	613	39	614	40
rect	613	40	614	41
rect	613	41	614	42
rect	613	42	614	43
rect	613	43	614	44
rect	613	44	614	45
rect	613	45	614	46
rect	613	46	614	47
rect	613	47	614	48
rect	613	48	614	49
rect	613	49	614	50
rect	613	50	614	51
rect	613	51	614	52
rect	613	52	614	53
rect	613	53	614	54
rect	613	54	614	55
rect	613	55	614	56
rect	613	56	614	57
rect	613	57	614	58
rect	613	58	614	59
rect	613	59	614	60
rect	613	60	614	61
rect	613	61	614	62
rect	613	62	614	63
rect	613	63	614	64
rect	613	64	614	65
rect	613	65	614	66
rect	613	66	614	67
rect	613	67	614	68
rect	613	68	614	69
rect	613	69	614	70
rect	613	70	614	71
rect	613	71	614	72
rect	613	72	614	73
rect	613	73	614	74
rect	613	74	614	75
rect	613	75	614	76
rect	613	76	614	77
rect	613	77	614	78
rect	613	78	614	79
rect	613	79	614	80
rect	613	80	614	81
rect	613	81	614	82
rect	613	82	614	83
rect	613	83	614	84
rect	613	84	614	85
rect	613	85	614	86
rect	613	86	614	87
rect	613	87	614	88
rect	613	88	614	89
rect	613	89	614	90
rect	613	90	614	91
rect	613	91	614	92
rect	613	92	614	93
rect	613	93	614	94
rect	613	94	614	95
rect	613	95	614	96
rect	613	96	614	97
rect	613	97	614	98
rect	613	98	614	99
rect	613	99	614	100
rect	613	100	614	101
rect	613	101	614	102
rect	613	102	614	103
rect	613	103	614	104
rect	613	104	614	105
rect	613	105	614	106
rect	613	106	614	107
rect	613	107	614	108
rect	613	108	614	109
rect	613	109	614	110
rect	613	110	614	111
rect	613	111	614	112
rect	613	112	614	113
rect	613	113	614	114
rect	613	114	614	115
rect	613	115	614	116
rect	613	116	614	117
rect	613	117	614	118
rect	613	118	614	119
rect	613	119	614	120
rect	613	120	614	121
rect	613	121	614	122
rect	613	122	614	123
rect	613	123	614	124
rect	613	124	614	125
rect	613	125	614	126
rect	613	126	614	127
rect	613	127	614	128
rect	613	128	614	129
rect	613	129	614	130
rect	613	130	614	131
rect	613	131	614	132
rect	613	132	614	133
rect	613	133	614	134
rect	613	134	614	135
rect	613	135	614	136
rect	613	136	614	137
rect	613	137	614	138
rect	613	138	614	139
rect	613	139	614	140
rect	613	140	614	141
rect	613	141	614	142
rect	613	142	614	143
rect	613	143	614	144
rect	613	144	614	145
rect	613	145	614	146
rect	613	146	614	147
rect	613	147	614	148
rect	613	148	614	149
rect	613	149	614	150
rect	613	150	614	151
rect	613	151	614	152
rect	613	152	614	153
rect	613	153	614	154
rect	613	154	614	155
rect	613	155	614	156
rect	613	156	614	157
rect	613	157	614	158
rect	613	158	614	159
rect	613	159	614	160
rect	613	160	614	161
rect	613	161	614	162
rect	613	162	614	163
rect	613	163	614	164
rect	613	164	614	165
rect	613	165	614	166
rect	613	166	614	167
rect	613	167	614	168
rect	613	168	614	169
rect	613	169	614	170
rect	613	170	614	171
rect	613	171	614	172
rect	613	172	614	173
rect	613	173	614	174
rect	613	174	614	175
rect	613	175	614	176
rect	613	176	614	177
rect	613	177	614	178
rect	613	178	614	179
rect	613	179	614	180
rect	613	180	614	181
rect	613	181	614	182
rect	613	182	614	183
rect	613	183	614	184
rect	613	184	614	185
rect	613	185	614	186
rect	613	186	614	187
rect	613	187	614	188
rect	613	188	614	189
rect	613	189	614	190
rect	613	190	614	191
rect	613	191	614	192
rect	613	192	614	193
rect	613	193	614	194
rect	613	194	614	195
rect	613	195	614	196
rect	613	196	614	197
rect	613	197	614	198
rect	613	198	614	199
rect	613	199	614	200
rect	613	200	614	201
rect	613	201	614	202
rect	613	202	614	203
rect	613	203	614	204
rect	613	204	614	205
rect	613	205	614	206
rect	613	206	614	207
rect	613	207	614	208
rect	613	208	614	209
rect	613	209	614	210
rect	613	210	614	211
rect	613	211	614	212
rect	613	212	614	213
rect	613	213	614	214
rect	613	214	614	215
rect	613	215	614	216
rect	613	216	614	217
rect	613	217	614	218
rect	613	218	614	219
rect	613	219	614	220
rect	613	220	614	221
rect	613	221	614	222
rect	613	222	614	223
rect	613	223	614	224
rect	613	224	614	225
rect	613	225	614	226
rect	613	226	614	227
rect	613	227	614	228
rect	613	228	614	229
rect	613	229	614	230
rect	613	230	614	231
rect	613	231	614	232
rect	613	232	614	233
rect	613	233	614	234
rect	613	234	614	235
rect	613	235	614	236
rect	613	236	614	237
rect	613	237	614	238
rect	613	238	614	239
rect	613	239	614	240
rect	614	0	615	1
rect	614	1	615	2
rect	614	2	615	3
rect	614	3	615	4
rect	614	4	615	5
rect	614	5	615	6
rect	614	6	615	7
rect	614	7	615	8
rect	614	8	615	9
rect	614	9	615	10
rect	614	10	615	11
rect	614	11	615	12
rect	614	12	615	13
rect	614	13	615	14
rect	614	14	615	15
rect	614	15	615	16
rect	614	16	615	17
rect	614	17	615	18
rect	614	18	615	19
rect	614	19	615	20
rect	614	20	615	21
rect	614	21	615	22
rect	614	22	615	23
rect	614	23	615	24
rect	614	24	615	25
rect	614	25	615	26
rect	614	26	615	27
rect	614	27	615	28
rect	614	28	615	29
rect	614	29	615	30
rect	614	30	615	31
rect	614	31	615	32
rect	614	32	615	33
rect	614	33	615	34
rect	614	34	615	35
rect	614	35	615	36
rect	614	36	615	37
rect	614	37	615	38
rect	614	38	615	39
rect	614	39	615	40
rect	614	40	615	41
rect	614	41	615	42
rect	614	42	615	43
rect	614	43	615	44
rect	614	44	615	45
rect	614	45	615	46
rect	614	46	615	47
rect	614	47	615	48
rect	614	48	615	49
rect	614	49	615	50
rect	614	50	615	51
rect	614	51	615	52
rect	614	52	615	53
rect	614	53	615	54
rect	614	54	615	55
rect	614	55	615	56
rect	614	56	615	57
rect	614	57	615	58
rect	614	58	615	59
rect	614	59	615	60
rect	614	60	615	61
rect	614	61	615	62
rect	614	62	615	63
rect	614	63	615	64
rect	614	64	615	65
rect	614	65	615	66
rect	614	66	615	67
rect	614	67	615	68
rect	614	68	615	69
rect	614	69	615	70
rect	614	70	615	71
rect	614	71	615	72
rect	614	72	615	73
rect	614	73	615	74
rect	614	74	615	75
rect	614	75	615	76
rect	614	76	615	77
rect	614	77	615	78
rect	614	78	615	79
rect	614	79	615	80
rect	614	80	615	81
rect	614	81	615	82
rect	614	82	615	83
rect	614	83	615	84
rect	614	84	615	85
rect	614	85	615	86
rect	614	86	615	87
rect	614	87	615	88
rect	614	88	615	89
rect	614	89	615	90
rect	614	90	615	91
rect	614	91	615	92
rect	614	92	615	93
rect	614	93	615	94
rect	614	94	615	95
rect	614	95	615	96
rect	614	96	615	97
rect	614	97	615	98
rect	614	98	615	99
rect	614	99	615	100
rect	614	100	615	101
rect	614	101	615	102
rect	614	102	615	103
rect	614	103	615	104
rect	614	104	615	105
rect	614	105	615	106
rect	614	106	615	107
rect	614	107	615	108
rect	614	108	615	109
rect	614	109	615	110
rect	614	110	615	111
rect	614	111	615	112
rect	614	112	615	113
rect	614	113	615	114
rect	614	114	615	115
rect	614	115	615	116
rect	614	116	615	117
rect	614	117	615	118
rect	614	118	615	119
rect	614	119	615	120
rect	614	120	615	121
rect	614	121	615	122
rect	614	122	615	123
rect	614	123	615	124
rect	614	124	615	125
rect	614	125	615	126
rect	614	126	615	127
rect	614	127	615	128
rect	614	128	615	129
rect	614	129	615	130
rect	614	130	615	131
rect	614	131	615	132
rect	614	132	615	133
rect	614	133	615	134
rect	614	134	615	135
rect	614	135	615	136
rect	614	136	615	137
rect	614	137	615	138
rect	614	138	615	139
rect	614	139	615	140
rect	614	140	615	141
rect	614	141	615	142
rect	614	142	615	143
rect	614	143	615	144
rect	614	144	615	145
rect	614	145	615	146
rect	614	146	615	147
rect	614	147	615	148
rect	614	148	615	149
rect	614	149	615	150
rect	614	150	615	151
rect	614	151	615	152
rect	614	152	615	153
rect	614	153	615	154
rect	614	154	615	155
rect	614	155	615	156
rect	614	156	615	157
rect	614	157	615	158
rect	614	158	615	159
rect	614	159	615	160
rect	614	160	615	161
rect	614	161	615	162
rect	614	162	615	163
rect	614	163	615	164
rect	614	164	615	165
rect	614	165	615	166
rect	614	166	615	167
rect	614	167	615	168
rect	614	168	615	169
rect	614	169	615	170
rect	614	170	615	171
rect	614	171	615	172
rect	614	172	615	173
rect	614	173	615	174
rect	614	174	615	175
rect	614	175	615	176
rect	614	176	615	177
rect	614	177	615	178
rect	614	178	615	179
rect	614	179	615	180
rect	614	180	615	181
rect	614	181	615	182
rect	614	182	615	183
rect	614	183	615	184
rect	614	184	615	185
rect	614	185	615	186
rect	614	186	615	187
rect	614	187	615	188
rect	614	188	615	189
rect	614	189	615	190
rect	614	190	615	191
rect	614	191	615	192
rect	614	192	615	193
rect	614	193	615	194
rect	614	194	615	195
rect	614	195	615	196
rect	614	196	615	197
rect	614	197	615	198
rect	614	198	615	199
rect	614	199	615	200
rect	614	200	615	201
rect	614	201	615	202
rect	614	202	615	203
rect	614	203	615	204
rect	614	204	615	205
rect	614	205	615	206
rect	614	206	615	207
rect	614	207	615	208
rect	614	208	615	209
rect	614	209	615	210
rect	614	210	615	211
rect	614	211	615	212
rect	614	212	615	213
rect	614	213	615	214
rect	614	214	615	215
rect	614	215	615	216
rect	614	216	615	217
rect	614	217	615	218
rect	614	218	615	219
rect	614	219	615	220
rect	614	220	615	221
rect	614	221	615	222
rect	614	222	615	223
rect	614	223	615	224
rect	614	224	615	225
rect	614	225	615	226
rect	614	226	615	227
rect	614	227	615	228
rect	614	228	615	229
rect	614	229	615	230
rect	614	230	615	231
rect	614	231	615	232
rect	614	232	615	233
rect	614	233	615	234
rect	614	234	615	235
rect	614	235	615	236
rect	614	236	615	237
rect	614	237	615	238
rect	614	238	615	239
rect	614	239	615	240
rect	615	0	616	1
rect	615	1	616	2
rect	615	2	616	3
rect	615	3	616	4
rect	615	4	616	5
rect	615	5	616	6
rect	615	6	616	7
rect	615	7	616	8
rect	615	8	616	9
rect	615	9	616	10
rect	615	10	616	11
rect	615	11	616	12
rect	615	12	616	13
rect	615	13	616	14
rect	615	14	616	15
rect	615	15	616	16
rect	615	16	616	17
rect	615	17	616	18
rect	615	18	616	19
rect	615	19	616	20
rect	615	20	616	21
rect	615	21	616	22
rect	615	22	616	23
rect	615	23	616	24
rect	615	24	616	25
rect	615	25	616	26
rect	615	26	616	27
rect	615	27	616	28
rect	615	28	616	29
rect	615	29	616	30
rect	615	30	616	31
rect	615	31	616	32
rect	615	32	616	33
rect	615	33	616	34
rect	615	34	616	35
rect	615	35	616	36
rect	615	36	616	37
rect	615	37	616	38
rect	615	38	616	39
rect	615	39	616	40
rect	615	40	616	41
rect	615	41	616	42
rect	615	42	616	43
rect	615	43	616	44
rect	615	44	616	45
rect	615	45	616	46
rect	615	46	616	47
rect	615	47	616	48
rect	615	48	616	49
rect	615	49	616	50
rect	615	50	616	51
rect	615	51	616	52
rect	615	52	616	53
rect	615	53	616	54
rect	615	54	616	55
rect	615	55	616	56
rect	615	56	616	57
rect	615	57	616	58
rect	615	58	616	59
rect	615	59	616	60
rect	615	60	616	61
rect	615	61	616	62
rect	615	62	616	63
rect	615	63	616	64
rect	615	64	616	65
rect	615	65	616	66
rect	615	66	616	67
rect	615	67	616	68
rect	615	68	616	69
rect	615	69	616	70
rect	615	70	616	71
rect	615	71	616	72
rect	615	72	616	73
rect	615	73	616	74
rect	615	74	616	75
rect	615	75	616	76
rect	615	76	616	77
rect	615	77	616	78
rect	615	78	616	79
rect	615	79	616	80
rect	615	80	616	81
rect	615	81	616	82
rect	615	82	616	83
rect	615	83	616	84
rect	615	84	616	85
rect	615	85	616	86
rect	615	86	616	87
rect	615	87	616	88
rect	615	88	616	89
rect	615	89	616	90
rect	615	90	616	91
rect	615	91	616	92
rect	615	92	616	93
rect	615	93	616	94
rect	615	94	616	95
rect	615	95	616	96
rect	615	96	616	97
rect	615	97	616	98
rect	615	98	616	99
rect	615	99	616	100
rect	615	100	616	101
rect	615	101	616	102
rect	615	102	616	103
rect	615	103	616	104
rect	615	104	616	105
rect	615	105	616	106
rect	615	106	616	107
rect	615	107	616	108
rect	615	108	616	109
rect	615	109	616	110
rect	615	110	616	111
rect	615	111	616	112
rect	615	112	616	113
rect	615	113	616	114
rect	615	114	616	115
rect	615	115	616	116
rect	615	116	616	117
rect	615	117	616	118
rect	615	118	616	119
rect	615	119	616	120
rect	615	120	616	121
rect	615	121	616	122
rect	615	122	616	123
rect	615	123	616	124
rect	615	124	616	125
rect	615	125	616	126
rect	615	126	616	127
rect	615	127	616	128
rect	615	128	616	129
rect	615	129	616	130
rect	615	130	616	131
rect	615	131	616	132
rect	615	132	616	133
rect	615	133	616	134
rect	615	134	616	135
rect	615	135	616	136
rect	615	136	616	137
rect	615	137	616	138
rect	615	138	616	139
rect	615	139	616	140
rect	615	140	616	141
rect	615	141	616	142
rect	615	142	616	143
rect	615	143	616	144
rect	615	144	616	145
rect	615	145	616	146
rect	615	146	616	147
rect	615	147	616	148
rect	615	148	616	149
rect	615	149	616	150
rect	615	150	616	151
rect	615	151	616	152
rect	615	152	616	153
rect	615	153	616	154
rect	615	154	616	155
rect	615	155	616	156
rect	615	156	616	157
rect	615	157	616	158
rect	615	158	616	159
rect	615	159	616	160
rect	615	160	616	161
rect	615	161	616	162
rect	615	162	616	163
rect	615	163	616	164
rect	615	164	616	165
rect	615	165	616	166
rect	615	166	616	167
rect	615	167	616	168
rect	615	168	616	169
rect	615	169	616	170
rect	615	170	616	171
rect	615	171	616	172
rect	615	172	616	173
rect	615	173	616	174
rect	615	174	616	175
rect	615	175	616	176
rect	615	176	616	177
rect	615	177	616	178
rect	615	178	616	179
rect	615	179	616	180
rect	615	180	616	181
rect	615	181	616	182
rect	615	182	616	183
rect	615	183	616	184
rect	615	184	616	185
rect	615	185	616	186
rect	615	186	616	187
rect	615	187	616	188
rect	615	188	616	189
rect	615	189	616	190
rect	615	190	616	191
rect	615	191	616	192
rect	615	192	616	193
rect	615	193	616	194
rect	615	194	616	195
rect	615	195	616	196
rect	615	196	616	197
rect	615	197	616	198
rect	615	198	616	199
rect	615	199	616	200
rect	615	200	616	201
rect	615	201	616	202
rect	615	202	616	203
rect	615	203	616	204
rect	615	204	616	205
rect	615	205	616	206
rect	615	206	616	207
rect	615	207	616	208
rect	615	208	616	209
rect	615	209	616	210
rect	615	210	616	211
rect	615	211	616	212
rect	615	212	616	213
rect	615	213	616	214
rect	615	214	616	215
rect	615	215	616	216
rect	615	216	616	217
rect	615	217	616	218
rect	615	218	616	219
rect	615	219	616	220
rect	615	220	616	221
rect	615	221	616	222
rect	615	222	616	223
rect	615	223	616	224
rect	615	224	616	225
rect	615	225	616	226
rect	615	226	616	227
rect	615	227	616	228
rect	615	228	616	229
rect	615	229	616	230
rect	615	230	616	231
rect	615	231	616	232
rect	615	232	616	233
rect	615	233	616	234
rect	615	234	616	235
rect	615	235	616	236
rect	615	236	616	237
rect	615	237	616	238
rect	615	238	616	239
rect	615	239	616	240
rect	616	0	617	1
rect	616	1	617	2
rect	616	2	617	3
rect	616	3	617	4
rect	616	4	617	5
rect	616	5	617	6
rect	616	6	617	7
rect	616	7	617	8
rect	616	8	617	9
rect	616	9	617	10
rect	616	10	617	11
rect	616	11	617	12
rect	616	12	617	13
rect	616	13	617	14
rect	616	14	617	15
rect	616	15	617	16
rect	616	16	617	17
rect	616	17	617	18
rect	616	18	617	19
rect	616	19	617	20
rect	616	20	617	21
rect	616	21	617	22
rect	616	22	617	23
rect	616	23	617	24
rect	616	24	617	25
rect	616	25	617	26
rect	616	26	617	27
rect	616	27	617	28
rect	616	28	617	29
rect	616	29	617	30
rect	616	30	617	31
rect	616	31	617	32
rect	616	32	617	33
rect	616	33	617	34
rect	616	34	617	35
rect	616	35	617	36
rect	616	36	617	37
rect	616	37	617	38
rect	616	38	617	39
rect	616	39	617	40
rect	616	40	617	41
rect	616	41	617	42
rect	616	42	617	43
rect	616	43	617	44
rect	616	44	617	45
rect	616	45	617	46
rect	616	46	617	47
rect	616	47	617	48
rect	616	48	617	49
rect	616	49	617	50
rect	616	50	617	51
rect	616	51	617	52
rect	616	52	617	53
rect	616	53	617	54
rect	616	54	617	55
rect	616	55	617	56
rect	616	56	617	57
rect	616	57	617	58
rect	616	58	617	59
rect	616	59	617	60
rect	616	60	617	61
rect	616	61	617	62
rect	616	62	617	63
rect	616	63	617	64
rect	616	64	617	65
rect	616	65	617	66
rect	616	66	617	67
rect	616	67	617	68
rect	616	68	617	69
rect	616	69	617	70
rect	616	70	617	71
rect	616	71	617	72
rect	616	72	617	73
rect	616	73	617	74
rect	616	74	617	75
rect	616	75	617	76
rect	616	76	617	77
rect	616	77	617	78
rect	616	78	617	79
rect	616	79	617	80
rect	616	80	617	81
rect	616	81	617	82
rect	616	82	617	83
rect	616	83	617	84
rect	616	84	617	85
rect	616	85	617	86
rect	616	86	617	87
rect	616	87	617	88
rect	616	88	617	89
rect	616	89	617	90
rect	616	90	617	91
rect	616	91	617	92
rect	616	92	617	93
rect	616	93	617	94
rect	616	94	617	95
rect	616	95	617	96
rect	616	96	617	97
rect	616	97	617	98
rect	616	98	617	99
rect	616	99	617	100
rect	616	100	617	101
rect	616	101	617	102
rect	616	102	617	103
rect	616	103	617	104
rect	616	104	617	105
rect	616	105	617	106
rect	616	106	617	107
rect	616	107	617	108
rect	616	108	617	109
rect	616	109	617	110
rect	616	110	617	111
rect	616	111	617	112
rect	616	112	617	113
rect	616	113	617	114
rect	616	114	617	115
rect	616	115	617	116
rect	616	116	617	117
rect	616	117	617	118
rect	616	118	617	119
rect	616	119	617	120
rect	616	120	617	121
rect	616	121	617	122
rect	616	122	617	123
rect	616	123	617	124
rect	616	124	617	125
rect	616	125	617	126
rect	616	126	617	127
rect	616	127	617	128
rect	616	128	617	129
rect	616	129	617	130
rect	616	130	617	131
rect	616	131	617	132
rect	616	132	617	133
rect	616	133	617	134
rect	616	134	617	135
rect	616	135	617	136
rect	616	136	617	137
rect	616	137	617	138
rect	616	138	617	139
rect	616	139	617	140
rect	616	140	617	141
rect	616	141	617	142
rect	616	142	617	143
rect	616	143	617	144
rect	616	144	617	145
rect	616	145	617	146
rect	616	146	617	147
rect	616	147	617	148
rect	616	148	617	149
rect	616	149	617	150
rect	616	150	617	151
rect	616	151	617	152
rect	616	152	617	153
rect	616	153	617	154
rect	616	154	617	155
rect	616	155	617	156
rect	616	156	617	157
rect	616	157	617	158
rect	616	158	617	159
rect	616	159	617	160
rect	616	160	617	161
rect	616	161	617	162
rect	616	162	617	163
rect	616	163	617	164
rect	616	164	617	165
rect	616	165	617	166
rect	616	166	617	167
rect	616	167	617	168
rect	616	168	617	169
rect	616	169	617	170
rect	616	170	617	171
rect	616	171	617	172
rect	616	172	617	173
rect	616	173	617	174
rect	616	174	617	175
rect	616	175	617	176
rect	616	176	617	177
rect	616	177	617	178
rect	616	178	617	179
rect	616	179	617	180
rect	616	180	617	181
rect	616	181	617	182
rect	616	182	617	183
rect	616	183	617	184
rect	616	184	617	185
rect	616	185	617	186
rect	616	186	617	187
rect	616	187	617	188
rect	616	188	617	189
rect	616	189	617	190
rect	616	190	617	191
rect	616	191	617	192
rect	616	192	617	193
rect	616	193	617	194
rect	616	194	617	195
rect	616	195	617	196
rect	616	196	617	197
rect	616	197	617	198
rect	616	198	617	199
rect	616	199	617	200
rect	616	200	617	201
rect	616	201	617	202
rect	616	202	617	203
rect	616	203	617	204
rect	616	204	617	205
rect	616	205	617	206
rect	616	206	617	207
rect	616	207	617	208
rect	616	208	617	209
rect	616	209	617	210
rect	616	210	617	211
rect	616	211	617	212
rect	616	212	617	213
rect	616	213	617	214
rect	616	214	617	215
rect	616	215	617	216
rect	616	216	617	217
rect	616	217	617	218
rect	616	218	617	219
rect	616	219	617	220
rect	616	220	617	221
rect	616	221	617	222
rect	616	222	617	223
rect	616	223	617	224
rect	616	224	617	225
rect	616	225	617	226
rect	616	226	617	227
rect	616	227	617	228
rect	616	228	617	229
rect	616	229	617	230
rect	616	230	617	231
rect	616	231	617	232
rect	616	232	617	233
rect	616	233	617	234
rect	616	234	617	235
rect	616	235	617	236
rect	616	236	617	237
rect	616	237	617	238
rect	616	238	617	239
rect	616	239	617	240
rect	617	0	618	1
rect	617	1	618	2
rect	617	2	618	3
rect	617	3	618	4
rect	617	4	618	5
rect	617	5	618	6
rect	617	6	618	7
rect	617	7	618	8
rect	617	8	618	9
rect	617	9	618	10
rect	617	10	618	11
rect	617	11	618	12
rect	617	12	618	13
rect	617	13	618	14
rect	617	14	618	15
rect	617	15	618	16
rect	617	16	618	17
rect	617	17	618	18
rect	617	18	618	19
rect	617	19	618	20
rect	617	20	618	21
rect	617	21	618	22
rect	617	22	618	23
rect	617	23	618	24
rect	617	24	618	25
rect	617	25	618	26
rect	617	26	618	27
rect	617	27	618	28
rect	617	28	618	29
rect	617	29	618	30
rect	617	30	618	31
rect	617	31	618	32
rect	617	32	618	33
rect	617	33	618	34
rect	617	34	618	35
rect	617	35	618	36
rect	617	36	618	37
rect	617	37	618	38
rect	617	38	618	39
rect	617	39	618	40
rect	617	40	618	41
rect	617	41	618	42
rect	617	42	618	43
rect	617	43	618	44
rect	617	44	618	45
rect	617	45	618	46
rect	617	46	618	47
rect	617	47	618	48
rect	617	48	618	49
rect	617	49	618	50
rect	617	50	618	51
rect	617	51	618	52
rect	617	52	618	53
rect	617	53	618	54
rect	617	54	618	55
rect	617	55	618	56
rect	617	56	618	57
rect	617	57	618	58
rect	617	58	618	59
rect	617	59	618	60
rect	617	60	618	61
rect	617	61	618	62
rect	617	62	618	63
rect	617	63	618	64
rect	617	64	618	65
rect	617	65	618	66
rect	617	66	618	67
rect	617	67	618	68
rect	617	68	618	69
rect	617	69	618	70
rect	617	70	618	71
rect	617	71	618	72
rect	617	72	618	73
rect	617	73	618	74
rect	617	74	618	75
rect	617	75	618	76
rect	617	76	618	77
rect	617	77	618	78
rect	617	78	618	79
rect	617	79	618	80
rect	617	80	618	81
rect	617	81	618	82
rect	617	82	618	83
rect	617	83	618	84
rect	617	84	618	85
rect	617	85	618	86
rect	617	86	618	87
rect	617	87	618	88
rect	617	88	618	89
rect	617	89	618	90
rect	617	90	618	91
rect	617	91	618	92
rect	617	92	618	93
rect	617	93	618	94
rect	617	94	618	95
rect	617	95	618	96
rect	617	96	618	97
rect	617	97	618	98
rect	617	98	618	99
rect	617	99	618	100
rect	617	100	618	101
rect	617	101	618	102
rect	617	102	618	103
rect	617	103	618	104
rect	617	104	618	105
rect	617	105	618	106
rect	617	106	618	107
rect	617	107	618	108
rect	617	108	618	109
rect	617	109	618	110
rect	617	110	618	111
rect	617	111	618	112
rect	617	112	618	113
rect	617	113	618	114
rect	617	114	618	115
rect	617	115	618	116
rect	617	116	618	117
rect	617	117	618	118
rect	617	118	618	119
rect	617	119	618	120
rect	617	120	618	121
rect	617	121	618	122
rect	617	122	618	123
rect	617	123	618	124
rect	617	124	618	125
rect	617	125	618	126
rect	617	126	618	127
rect	617	127	618	128
rect	617	128	618	129
rect	617	129	618	130
rect	617	130	618	131
rect	617	131	618	132
rect	617	132	618	133
rect	617	133	618	134
rect	617	134	618	135
rect	617	135	618	136
rect	617	136	618	137
rect	617	137	618	138
rect	617	138	618	139
rect	617	139	618	140
rect	617	140	618	141
rect	617	141	618	142
rect	617	142	618	143
rect	617	143	618	144
rect	617	144	618	145
rect	617	145	618	146
rect	617	146	618	147
rect	617	147	618	148
rect	617	148	618	149
rect	617	149	618	150
rect	617	150	618	151
rect	617	151	618	152
rect	617	152	618	153
rect	617	153	618	154
rect	617	154	618	155
rect	617	155	618	156
rect	617	156	618	157
rect	617	157	618	158
rect	617	158	618	159
rect	617	159	618	160
rect	617	160	618	161
rect	617	161	618	162
rect	617	162	618	163
rect	617	163	618	164
rect	617	164	618	165
rect	617	165	618	166
rect	617	166	618	167
rect	617	167	618	168
rect	617	168	618	169
rect	617	169	618	170
rect	617	170	618	171
rect	617	171	618	172
rect	617	172	618	173
rect	617	173	618	174
rect	617	174	618	175
rect	617	175	618	176
rect	617	176	618	177
rect	617	177	618	178
rect	617	178	618	179
rect	617	179	618	180
rect	617	180	618	181
rect	617	181	618	182
rect	617	182	618	183
rect	617	183	618	184
rect	617	184	618	185
rect	617	185	618	186
rect	617	186	618	187
rect	617	187	618	188
rect	617	188	618	189
rect	617	189	618	190
rect	617	190	618	191
rect	617	191	618	192
rect	617	192	618	193
rect	617	193	618	194
rect	617	194	618	195
rect	617	195	618	196
rect	617	196	618	197
rect	617	197	618	198
rect	617	198	618	199
rect	617	199	618	200
rect	617	200	618	201
rect	617	201	618	202
rect	617	202	618	203
rect	617	203	618	204
rect	617	204	618	205
rect	617	205	618	206
rect	617	206	618	207
rect	617	207	618	208
rect	617	208	618	209
rect	617	209	618	210
rect	617	210	618	211
rect	617	211	618	212
rect	617	212	618	213
rect	617	213	618	214
rect	617	214	618	215
rect	617	215	618	216
rect	617	216	618	217
rect	617	217	618	218
rect	617	218	618	219
rect	617	219	618	220
rect	617	220	618	221
rect	617	221	618	222
rect	617	222	618	223
rect	617	223	618	224
rect	617	224	618	225
rect	617	225	618	226
rect	617	226	618	227
rect	617	227	618	228
rect	617	228	618	229
rect	617	229	618	230
rect	617	230	618	231
rect	617	231	618	232
rect	617	232	618	233
rect	617	233	618	234
rect	617	234	618	235
rect	617	235	618	236
rect	617	236	618	237
rect	617	237	618	238
rect	617	238	618	239
rect	617	239	618	240
rect	629	0	630	1
rect	629	1	630	2
rect	629	2	630	3
rect	629	3	630	4
rect	629	4	630	5
rect	629	5	630	6
rect	629	6	630	7
rect	629	7	630	8
rect	629	8	630	9
rect	629	9	630	10
rect	629	10	630	11
rect	629	11	630	12
rect	629	12	630	13
rect	629	13	630	14
rect	629	14	630	15
rect	629	15	630	16
rect	629	16	630	17
rect	629	17	630	18
rect	629	18	630	19
rect	629	19	630	20
rect	629	20	630	21
rect	629	21	630	22
rect	629	22	630	23
rect	629	23	630	24
rect	629	24	630	25
rect	629	25	630	26
rect	629	26	630	27
rect	629	27	630	28
rect	629	28	630	29
rect	629	29	630	30
rect	629	30	630	31
rect	629	31	630	32
rect	629	32	630	33
rect	629	33	630	34
rect	629	34	630	35
rect	629	35	630	36
rect	629	36	630	37
rect	629	37	630	38
rect	629	38	630	39
rect	629	39	630	40
rect	629	40	630	41
rect	629	41	630	42
rect	629	42	630	43
rect	629	43	630	44
rect	629	44	630	45
rect	629	45	630	46
rect	629	46	630	47
rect	629	47	630	48
rect	629	48	630	49
rect	629	49	630	50
rect	629	50	630	51
rect	629	51	630	52
rect	629	52	630	53
rect	629	53	630	54
rect	629	54	630	55
rect	629	55	630	56
rect	629	56	630	57
rect	629	57	630	58
rect	629	58	630	59
rect	629	59	630	60
rect	629	60	630	61
rect	629	61	630	62
rect	629	62	630	63
rect	629	63	630	64
rect	629	64	630	65
rect	629	65	630	66
rect	629	66	630	67
rect	629	67	630	68
rect	629	68	630	69
rect	629	69	630	70
rect	629	70	630	71
rect	629	71	630	72
rect	629	72	630	73
rect	629	73	630	74
rect	629	74	630	75
rect	629	75	630	76
rect	629	76	630	77
rect	629	77	630	78
rect	629	78	630	79
rect	629	79	630	80
rect	629	80	630	81
rect	629	81	630	82
rect	629	82	630	83
rect	629	83	630	84
rect	629	84	630	85
rect	629	85	630	86
rect	629	86	630	87
rect	629	87	630	88
rect	629	88	630	89
rect	629	89	630	90
rect	629	90	630	91
rect	629	91	630	92
rect	629	92	630	93
rect	629	93	630	94
rect	629	94	630	95
rect	629	95	630	96
rect	629	96	630	97
rect	629	97	630	98
rect	629	98	630	99
rect	629	99	630	100
rect	629	100	630	101
rect	629	101	630	102
rect	629	102	630	103
rect	629	103	630	104
rect	629	104	630	105
rect	629	105	630	106
rect	629	106	630	107
rect	629	107	630	108
rect	629	108	630	109
rect	629	109	630	110
rect	629	110	630	111
rect	629	111	630	112
rect	629	112	630	113
rect	629	113	630	114
rect	629	114	630	115
rect	629	115	630	116
rect	629	116	630	117
rect	629	117	630	118
rect	629	118	630	119
rect	629	119	630	120
rect	629	120	630	121
rect	629	121	630	122
rect	629	122	630	123
rect	629	123	630	124
rect	629	124	630	125
rect	629	125	630	126
rect	629	126	630	127
rect	629	127	630	128
rect	629	128	630	129
rect	629	129	630	130
rect	629	130	630	131
rect	629	131	630	132
rect	629	132	630	133
rect	629	133	630	134
rect	629	134	630	135
rect	629	135	630	136
rect	629	136	630	137
rect	629	137	630	138
rect	629	138	630	139
rect	629	139	630	140
rect	629	140	630	141
rect	629	141	630	142
rect	629	142	630	143
rect	629	143	630	144
rect	629	144	630	145
rect	629	145	630	146
rect	629	146	630	147
rect	629	147	630	148
rect	629	148	630	149
rect	629	149	630	150
rect	629	150	630	151
rect	629	151	630	152
rect	629	152	630	153
rect	629	153	630	154
rect	629	154	630	155
rect	629	155	630	156
rect	629	156	630	157
rect	629	157	630	158
rect	629	158	630	159
rect	629	159	630	160
rect	629	160	630	161
rect	629	161	630	162
rect	629	162	630	163
rect	629	163	630	164
rect	629	164	630	165
rect	629	165	630	166
rect	629	166	630	167
rect	629	167	630	168
rect	629	168	630	169
rect	629	169	630	170
rect	629	170	630	171
rect	629	171	630	172
rect	629	172	630	173
rect	629	173	630	174
rect	629	174	630	175
rect	629	175	630	176
rect	629	176	630	177
rect	629	177	630	178
rect	629	178	630	179
rect	629	179	630	180
rect	629	180	630	181
rect	629	181	630	182
rect	629	182	630	183
rect	629	183	630	184
rect	629	184	630	185
rect	629	185	630	186
rect	629	186	630	187
rect	629	187	630	188
rect	629	188	630	189
rect	629	189	630	190
rect	629	190	630	191
rect	629	191	630	192
rect	629	192	630	193
rect	629	193	630	194
rect	629	194	630	195
rect	629	195	630	196
rect	629	196	630	197
rect	629	197	630	198
rect	629	198	630	199
rect	629	199	630	200
rect	629	200	630	201
rect	629	201	630	202
rect	629	202	630	203
rect	629	203	630	204
rect	629	204	630	205
rect	629	205	630	206
rect	629	206	630	207
rect	629	207	630	208
rect	629	208	630	209
rect	629	209	630	210
rect	629	210	630	211
rect	629	211	630	212
rect	629	212	630	213
rect	629	213	630	214
rect	629	214	630	215
rect	629	215	630	216
rect	629	216	630	217
rect	629	217	630	218
rect	629	218	630	219
rect	630	0	631	1
rect	630	1	631	2
rect	630	2	631	3
rect	630	3	631	4
rect	630	4	631	5
rect	630	5	631	6
rect	630	6	631	7
rect	630	7	631	8
rect	630	8	631	9
rect	630	9	631	10
rect	630	10	631	11
rect	630	11	631	12
rect	630	12	631	13
rect	630	13	631	14
rect	630	14	631	15
rect	630	15	631	16
rect	630	16	631	17
rect	630	17	631	18
rect	630	18	631	19
rect	630	19	631	20
rect	630	20	631	21
rect	630	21	631	22
rect	630	22	631	23
rect	630	23	631	24
rect	630	24	631	25
rect	630	25	631	26
rect	630	26	631	27
rect	630	27	631	28
rect	630	28	631	29
rect	630	29	631	30
rect	630	30	631	31
rect	630	31	631	32
rect	630	32	631	33
rect	630	33	631	34
rect	630	34	631	35
rect	630	35	631	36
rect	630	36	631	37
rect	630	37	631	38
rect	630	38	631	39
rect	630	39	631	40
rect	630	40	631	41
rect	630	41	631	42
rect	630	42	631	43
rect	630	43	631	44
rect	630	44	631	45
rect	630	45	631	46
rect	630	46	631	47
rect	630	47	631	48
rect	630	48	631	49
rect	630	49	631	50
rect	630	50	631	51
rect	630	51	631	52
rect	630	52	631	53
rect	630	53	631	54
rect	630	54	631	55
rect	630	55	631	56
rect	630	56	631	57
rect	630	57	631	58
rect	630	58	631	59
rect	630	59	631	60
rect	630	60	631	61
rect	630	61	631	62
rect	630	62	631	63
rect	630	63	631	64
rect	630	64	631	65
rect	630	65	631	66
rect	630	66	631	67
rect	630	67	631	68
rect	630	68	631	69
rect	630	69	631	70
rect	630	70	631	71
rect	630	71	631	72
rect	630	72	631	73
rect	630	73	631	74
rect	630	74	631	75
rect	630	75	631	76
rect	630	76	631	77
rect	630	77	631	78
rect	630	78	631	79
rect	630	79	631	80
rect	630	80	631	81
rect	630	81	631	82
rect	630	82	631	83
rect	630	83	631	84
rect	630	84	631	85
rect	630	85	631	86
rect	630	86	631	87
rect	630	87	631	88
rect	630	88	631	89
rect	630	89	631	90
rect	630	90	631	91
rect	630	91	631	92
rect	630	92	631	93
rect	630	93	631	94
rect	630	94	631	95
rect	630	95	631	96
rect	630	96	631	97
rect	630	97	631	98
rect	630	98	631	99
rect	630	99	631	100
rect	630	100	631	101
rect	630	101	631	102
rect	630	102	631	103
rect	630	103	631	104
rect	630	104	631	105
rect	630	105	631	106
rect	630	106	631	107
rect	630	107	631	108
rect	630	108	631	109
rect	630	109	631	110
rect	630	110	631	111
rect	630	111	631	112
rect	630	112	631	113
rect	630	113	631	114
rect	630	114	631	115
rect	630	115	631	116
rect	630	116	631	117
rect	630	117	631	118
rect	630	118	631	119
rect	630	119	631	120
rect	630	120	631	121
rect	630	121	631	122
rect	630	122	631	123
rect	630	123	631	124
rect	630	124	631	125
rect	630	125	631	126
rect	630	126	631	127
rect	630	127	631	128
rect	630	128	631	129
rect	630	129	631	130
rect	630	130	631	131
rect	630	131	631	132
rect	630	132	631	133
rect	630	133	631	134
rect	630	134	631	135
rect	630	135	631	136
rect	630	136	631	137
rect	630	137	631	138
rect	630	138	631	139
rect	630	139	631	140
rect	630	140	631	141
rect	630	141	631	142
rect	630	142	631	143
rect	630	143	631	144
rect	630	144	631	145
rect	630	145	631	146
rect	630	146	631	147
rect	630	147	631	148
rect	630	148	631	149
rect	630	149	631	150
rect	630	150	631	151
rect	630	151	631	152
rect	630	152	631	153
rect	630	153	631	154
rect	630	154	631	155
rect	630	155	631	156
rect	630	156	631	157
rect	630	157	631	158
rect	630	158	631	159
rect	630	159	631	160
rect	630	160	631	161
rect	630	161	631	162
rect	630	162	631	163
rect	630	163	631	164
rect	630	164	631	165
rect	630	165	631	166
rect	630	166	631	167
rect	630	167	631	168
rect	630	168	631	169
rect	630	169	631	170
rect	630	170	631	171
rect	630	171	631	172
rect	630	172	631	173
rect	630	173	631	174
rect	630	174	631	175
rect	630	175	631	176
rect	630	176	631	177
rect	630	177	631	178
rect	630	178	631	179
rect	630	179	631	180
rect	630	180	631	181
rect	630	181	631	182
rect	630	182	631	183
rect	630	183	631	184
rect	630	184	631	185
rect	630	185	631	186
rect	630	186	631	187
rect	630	187	631	188
rect	630	188	631	189
rect	630	189	631	190
rect	630	190	631	191
rect	630	191	631	192
rect	630	192	631	193
rect	630	193	631	194
rect	630	194	631	195
rect	630	195	631	196
rect	630	196	631	197
rect	630	197	631	198
rect	630	198	631	199
rect	630	199	631	200
rect	630	200	631	201
rect	630	201	631	202
rect	630	202	631	203
rect	630	203	631	204
rect	630	204	631	205
rect	630	205	631	206
rect	630	206	631	207
rect	630	207	631	208
rect	630	208	631	209
rect	630	209	631	210
rect	630	210	631	211
rect	630	211	631	212
rect	630	212	631	213
rect	630	213	631	214
rect	630	214	631	215
rect	630	215	631	216
rect	630	216	631	217
rect	630	217	631	218
rect	630	218	631	219
rect	631	0	632	1
rect	631	1	632	2
rect	631	2	632	3
rect	631	3	632	4
rect	631	4	632	5
rect	631	5	632	6
rect	631	6	632	7
rect	631	7	632	8
rect	631	8	632	9
rect	631	9	632	10
rect	631	10	632	11
rect	631	11	632	12
rect	631	12	632	13
rect	631	13	632	14
rect	631	14	632	15
rect	631	15	632	16
rect	631	16	632	17
rect	631	17	632	18
rect	631	18	632	19
rect	631	19	632	20
rect	631	20	632	21
rect	631	21	632	22
rect	631	22	632	23
rect	631	23	632	24
rect	631	24	632	25
rect	631	25	632	26
rect	631	26	632	27
rect	631	27	632	28
rect	631	28	632	29
rect	631	29	632	30
rect	631	30	632	31
rect	631	31	632	32
rect	631	32	632	33
rect	631	33	632	34
rect	631	34	632	35
rect	631	35	632	36
rect	631	36	632	37
rect	631	37	632	38
rect	631	38	632	39
rect	631	39	632	40
rect	631	40	632	41
rect	631	41	632	42
rect	631	42	632	43
rect	631	43	632	44
rect	631	44	632	45
rect	631	45	632	46
rect	631	46	632	47
rect	631	47	632	48
rect	631	48	632	49
rect	631	49	632	50
rect	631	50	632	51
rect	631	51	632	52
rect	631	52	632	53
rect	631	53	632	54
rect	631	54	632	55
rect	631	55	632	56
rect	631	56	632	57
rect	631	57	632	58
rect	631	58	632	59
rect	631	59	632	60
rect	631	60	632	61
rect	631	61	632	62
rect	631	62	632	63
rect	631	63	632	64
rect	631	64	632	65
rect	631	65	632	66
rect	631	66	632	67
rect	631	67	632	68
rect	631	68	632	69
rect	631	69	632	70
rect	631	70	632	71
rect	631	71	632	72
rect	631	72	632	73
rect	631	73	632	74
rect	631	74	632	75
rect	631	75	632	76
rect	631	76	632	77
rect	631	77	632	78
rect	631	78	632	79
rect	631	79	632	80
rect	631	80	632	81
rect	631	81	632	82
rect	631	82	632	83
rect	631	83	632	84
rect	631	84	632	85
rect	631	85	632	86
rect	631	86	632	87
rect	631	87	632	88
rect	631	88	632	89
rect	631	89	632	90
rect	631	90	632	91
rect	631	91	632	92
rect	631	92	632	93
rect	631	93	632	94
rect	631	94	632	95
rect	631	95	632	96
rect	631	96	632	97
rect	631	97	632	98
rect	631	98	632	99
rect	631	99	632	100
rect	631	100	632	101
rect	631	101	632	102
rect	631	102	632	103
rect	631	103	632	104
rect	631	104	632	105
rect	631	105	632	106
rect	631	106	632	107
rect	631	107	632	108
rect	631	108	632	109
rect	631	109	632	110
rect	631	110	632	111
rect	631	111	632	112
rect	631	112	632	113
rect	631	113	632	114
rect	631	114	632	115
rect	631	115	632	116
rect	631	116	632	117
rect	631	117	632	118
rect	631	118	632	119
rect	631	119	632	120
rect	631	120	632	121
rect	631	121	632	122
rect	631	122	632	123
rect	631	123	632	124
rect	631	124	632	125
rect	631	125	632	126
rect	631	126	632	127
rect	631	127	632	128
rect	631	128	632	129
rect	631	129	632	130
rect	631	130	632	131
rect	631	131	632	132
rect	631	132	632	133
rect	631	133	632	134
rect	631	134	632	135
rect	631	135	632	136
rect	631	136	632	137
rect	631	137	632	138
rect	631	138	632	139
rect	631	139	632	140
rect	631	140	632	141
rect	631	141	632	142
rect	631	142	632	143
rect	631	143	632	144
rect	631	144	632	145
rect	631	145	632	146
rect	631	146	632	147
rect	631	147	632	148
rect	631	148	632	149
rect	631	149	632	150
rect	631	150	632	151
rect	631	151	632	152
rect	631	152	632	153
rect	631	153	632	154
rect	631	154	632	155
rect	631	155	632	156
rect	631	156	632	157
rect	631	157	632	158
rect	631	158	632	159
rect	631	159	632	160
rect	631	160	632	161
rect	631	161	632	162
rect	631	162	632	163
rect	631	163	632	164
rect	631	164	632	165
rect	631	165	632	166
rect	631	166	632	167
rect	631	167	632	168
rect	631	168	632	169
rect	631	169	632	170
rect	631	170	632	171
rect	631	171	632	172
rect	631	172	632	173
rect	631	173	632	174
rect	631	174	632	175
rect	631	175	632	176
rect	631	176	632	177
rect	631	177	632	178
rect	631	178	632	179
rect	631	179	632	180
rect	631	180	632	181
rect	631	181	632	182
rect	631	182	632	183
rect	631	183	632	184
rect	631	184	632	185
rect	631	185	632	186
rect	631	186	632	187
rect	631	187	632	188
rect	631	188	632	189
rect	631	189	632	190
rect	631	190	632	191
rect	631	191	632	192
rect	631	192	632	193
rect	631	193	632	194
rect	631	194	632	195
rect	631	195	632	196
rect	631	196	632	197
rect	631	197	632	198
rect	631	198	632	199
rect	631	199	632	200
rect	631	200	632	201
rect	631	201	632	202
rect	631	202	632	203
rect	631	203	632	204
rect	631	204	632	205
rect	631	205	632	206
rect	631	206	632	207
rect	631	207	632	208
rect	631	208	632	209
rect	631	209	632	210
rect	631	210	632	211
rect	631	211	632	212
rect	631	212	632	213
rect	631	213	632	214
rect	631	214	632	215
rect	631	215	632	216
rect	631	216	632	217
rect	631	217	632	218
rect	631	218	632	219
rect	632	0	633	1
rect	632	1	633	2
rect	632	2	633	3
rect	632	3	633	4
rect	632	4	633	5
rect	632	5	633	6
rect	632	6	633	7
rect	632	7	633	8
rect	632	8	633	9
rect	632	9	633	10
rect	632	10	633	11
rect	632	11	633	12
rect	632	12	633	13
rect	632	13	633	14
rect	632	14	633	15
rect	632	15	633	16
rect	632	16	633	17
rect	632	17	633	18
rect	632	18	633	19
rect	632	19	633	20
rect	632	20	633	21
rect	632	21	633	22
rect	632	22	633	23
rect	632	23	633	24
rect	632	24	633	25
rect	632	25	633	26
rect	632	26	633	27
rect	632	27	633	28
rect	632	28	633	29
rect	632	29	633	30
rect	632	30	633	31
rect	632	31	633	32
rect	632	32	633	33
rect	632	33	633	34
rect	632	34	633	35
rect	632	35	633	36
rect	632	36	633	37
rect	632	37	633	38
rect	632	38	633	39
rect	632	39	633	40
rect	632	40	633	41
rect	632	41	633	42
rect	632	42	633	43
rect	632	43	633	44
rect	632	44	633	45
rect	632	45	633	46
rect	632	46	633	47
rect	632	47	633	48
rect	632	48	633	49
rect	632	49	633	50
rect	632	50	633	51
rect	632	51	633	52
rect	632	52	633	53
rect	632	53	633	54
rect	632	54	633	55
rect	632	55	633	56
rect	632	56	633	57
rect	632	57	633	58
rect	632	58	633	59
rect	632	59	633	60
rect	632	60	633	61
rect	632	61	633	62
rect	632	62	633	63
rect	632	63	633	64
rect	632	64	633	65
rect	632	65	633	66
rect	632	66	633	67
rect	632	67	633	68
rect	632	68	633	69
rect	632	69	633	70
rect	632	70	633	71
rect	632	71	633	72
rect	632	72	633	73
rect	632	73	633	74
rect	632	74	633	75
rect	632	75	633	76
rect	632	76	633	77
rect	632	77	633	78
rect	632	78	633	79
rect	632	79	633	80
rect	632	80	633	81
rect	632	81	633	82
rect	632	82	633	83
rect	632	83	633	84
rect	632	84	633	85
rect	632	85	633	86
rect	632	86	633	87
rect	632	87	633	88
rect	632	88	633	89
rect	632	89	633	90
rect	632	90	633	91
rect	632	91	633	92
rect	632	92	633	93
rect	632	93	633	94
rect	632	94	633	95
rect	632	95	633	96
rect	632	96	633	97
rect	632	97	633	98
rect	632	98	633	99
rect	632	99	633	100
rect	632	100	633	101
rect	632	101	633	102
rect	632	102	633	103
rect	632	103	633	104
rect	632	104	633	105
rect	632	105	633	106
rect	632	106	633	107
rect	632	107	633	108
rect	632	108	633	109
rect	632	109	633	110
rect	632	110	633	111
rect	632	111	633	112
rect	632	112	633	113
rect	632	113	633	114
rect	632	114	633	115
rect	632	115	633	116
rect	632	116	633	117
rect	632	117	633	118
rect	632	118	633	119
rect	632	119	633	120
rect	632	120	633	121
rect	632	121	633	122
rect	632	122	633	123
rect	632	123	633	124
rect	632	124	633	125
rect	632	125	633	126
rect	632	126	633	127
rect	632	127	633	128
rect	632	128	633	129
rect	632	129	633	130
rect	632	130	633	131
rect	632	131	633	132
rect	632	132	633	133
rect	632	133	633	134
rect	632	134	633	135
rect	632	135	633	136
rect	632	136	633	137
rect	632	137	633	138
rect	632	138	633	139
rect	632	139	633	140
rect	632	140	633	141
rect	632	141	633	142
rect	632	142	633	143
rect	632	143	633	144
rect	632	144	633	145
rect	632	145	633	146
rect	632	146	633	147
rect	632	147	633	148
rect	632	148	633	149
rect	632	149	633	150
rect	632	150	633	151
rect	632	151	633	152
rect	632	152	633	153
rect	632	153	633	154
rect	632	154	633	155
rect	632	155	633	156
rect	632	156	633	157
rect	632	157	633	158
rect	632	158	633	159
rect	632	159	633	160
rect	632	160	633	161
rect	632	161	633	162
rect	632	162	633	163
rect	632	163	633	164
rect	632	164	633	165
rect	632	165	633	166
rect	632	166	633	167
rect	632	167	633	168
rect	632	168	633	169
rect	632	169	633	170
rect	632	170	633	171
rect	632	171	633	172
rect	632	172	633	173
rect	632	173	633	174
rect	632	174	633	175
rect	632	175	633	176
rect	632	176	633	177
rect	632	177	633	178
rect	632	178	633	179
rect	632	179	633	180
rect	632	180	633	181
rect	632	181	633	182
rect	632	182	633	183
rect	632	183	633	184
rect	632	184	633	185
rect	632	185	633	186
rect	632	186	633	187
rect	632	187	633	188
rect	632	188	633	189
rect	632	189	633	190
rect	632	190	633	191
rect	632	191	633	192
rect	632	192	633	193
rect	632	193	633	194
rect	632	194	633	195
rect	632	195	633	196
rect	632	196	633	197
rect	632	197	633	198
rect	632	198	633	199
rect	632	199	633	200
rect	632	200	633	201
rect	632	201	633	202
rect	632	202	633	203
rect	632	203	633	204
rect	632	204	633	205
rect	632	205	633	206
rect	632	206	633	207
rect	632	207	633	208
rect	632	208	633	209
rect	632	209	633	210
rect	632	210	633	211
rect	632	211	633	212
rect	632	212	633	213
rect	632	213	633	214
rect	632	214	633	215
rect	632	215	633	216
rect	632	216	633	217
rect	632	217	633	218
rect	632	218	633	219
rect	633	0	634	1
rect	633	1	634	2
rect	633	2	634	3
rect	633	3	634	4
rect	633	4	634	5
rect	633	5	634	6
rect	633	6	634	7
rect	633	7	634	8
rect	633	8	634	9
rect	633	9	634	10
rect	633	10	634	11
rect	633	11	634	12
rect	633	12	634	13
rect	633	13	634	14
rect	633	14	634	15
rect	633	15	634	16
rect	633	16	634	17
rect	633	17	634	18
rect	633	18	634	19
rect	633	19	634	20
rect	633	20	634	21
rect	633	21	634	22
rect	633	22	634	23
rect	633	23	634	24
rect	633	24	634	25
rect	633	25	634	26
rect	633	26	634	27
rect	633	27	634	28
rect	633	28	634	29
rect	633	29	634	30
rect	633	30	634	31
rect	633	31	634	32
rect	633	32	634	33
rect	633	33	634	34
rect	633	34	634	35
rect	633	35	634	36
rect	633	36	634	37
rect	633	37	634	38
rect	633	38	634	39
rect	633	39	634	40
rect	633	40	634	41
rect	633	41	634	42
rect	633	42	634	43
rect	633	43	634	44
rect	633	44	634	45
rect	633	45	634	46
rect	633	46	634	47
rect	633	47	634	48
rect	633	48	634	49
rect	633	49	634	50
rect	633	50	634	51
rect	633	51	634	52
rect	633	52	634	53
rect	633	53	634	54
rect	633	54	634	55
rect	633	55	634	56
rect	633	56	634	57
rect	633	57	634	58
rect	633	58	634	59
rect	633	59	634	60
rect	633	60	634	61
rect	633	61	634	62
rect	633	62	634	63
rect	633	63	634	64
rect	633	64	634	65
rect	633	65	634	66
rect	633	66	634	67
rect	633	67	634	68
rect	633	68	634	69
rect	633	69	634	70
rect	633	70	634	71
rect	633	71	634	72
rect	633	72	634	73
rect	633	73	634	74
rect	633	74	634	75
rect	633	75	634	76
rect	633	76	634	77
rect	633	77	634	78
rect	633	78	634	79
rect	633	79	634	80
rect	633	80	634	81
rect	633	81	634	82
rect	633	82	634	83
rect	633	83	634	84
rect	633	84	634	85
rect	633	85	634	86
rect	633	86	634	87
rect	633	87	634	88
rect	633	88	634	89
rect	633	89	634	90
rect	633	90	634	91
rect	633	91	634	92
rect	633	92	634	93
rect	633	93	634	94
rect	633	94	634	95
rect	633	95	634	96
rect	633	96	634	97
rect	633	97	634	98
rect	633	98	634	99
rect	633	99	634	100
rect	633	100	634	101
rect	633	101	634	102
rect	633	102	634	103
rect	633	103	634	104
rect	633	104	634	105
rect	633	105	634	106
rect	633	106	634	107
rect	633	107	634	108
rect	633	108	634	109
rect	633	109	634	110
rect	633	110	634	111
rect	633	111	634	112
rect	633	112	634	113
rect	633	113	634	114
rect	633	114	634	115
rect	633	115	634	116
rect	633	116	634	117
rect	633	117	634	118
rect	633	118	634	119
rect	633	119	634	120
rect	633	120	634	121
rect	633	121	634	122
rect	633	122	634	123
rect	633	123	634	124
rect	633	124	634	125
rect	633	125	634	126
rect	633	126	634	127
rect	633	127	634	128
rect	633	128	634	129
rect	633	129	634	130
rect	633	130	634	131
rect	633	131	634	132
rect	633	132	634	133
rect	633	133	634	134
rect	633	134	634	135
rect	633	135	634	136
rect	633	136	634	137
rect	633	137	634	138
rect	633	138	634	139
rect	633	139	634	140
rect	633	140	634	141
rect	633	141	634	142
rect	633	142	634	143
rect	633	143	634	144
rect	633	144	634	145
rect	633	145	634	146
rect	633	146	634	147
rect	633	147	634	148
rect	633	148	634	149
rect	633	149	634	150
rect	633	150	634	151
rect	633	151	634	152
rect	633	152	634	153
rect	633	153	634	154
rect	633	154	634	155
rect	633	155	634	156
rect	633	156	634	157
rect	633	157	634	158
rect	633	158	634	159
rect	633	159	634	160
rect	633	160	634	161
rect	633	161	634	162
rect	633	162	634	163
rect	633	163	634	164
rect	633	164	634	165
rect	633	165	634	166
rect	633	166	634	167
rect	633	167	634	168
rect	633	168	634	169
rect	633	169	634	170
rect	633	170	634	171
rect	633	171	634	172
rect	633	172	634	173
rect	633	173	634	174
rect	633	174	634	175
rect	633	175	634	176
rect	633	176	634	177
rect	633	177	634	178
rect	633	178	634	179
rect	633	179	634	180
rect	633	180	634	181
rect	633	181	634	182
rect	633	182	634	183
rect	633	183	634	184
rect	633	184	634	185
rect	633	185	634	186
rect	633	186	634	187
rect	633	187	634	188
rect	633	188	634	189
rect	633	189	634	190
rect	633	190	634	191
rect	633	191	634	192
rect	633	192	634	193
rect	633	193	634	194
rect	633	194	634	195
rect	633	195	634	196
rect	633	196	634	197
rect	633	197	634	198
rect	633	198	634	199
rect	633	199	634	200
rect	633	200	634	201
rect	633	201	634	202
rect	633	202	634	203
rect	633	203	634	204
rect	633	204	634	205
rect	633	205	634	206
rect	633	206	634	207
rect	633	207	634	208
rect	633	208	634	209
rect	633	209	634	210
rect	633	210	634	211
rect	633	211	634	212
rect	633	212	634	213
rect	633	213	634	214
rect	633	214	634	215
rect	633	215	634	216
rect	633	216	634	217
rect	633	217	634	218
rect	633	218	634	219
rect	634	0	635	1
rect	634	1	635	2
rect	634	2	635	3
rect	634	3	635	4
rect	634	4	635	5
rect	634	5	635	6
rect	634	6	635	7
rect	634	7	635	8
rect	634	8	635	9
rect	634	9	635	10
rect	634	10	635	11
rect	634	11	635	12
rect	634	12	635	13
rect	634	13	635	14
rect	634	14	635	15
rect	634	15	635	16
rect	634	16	635	17
rect	634	17	635	18
rect	634	18	635	19
rect	634	19	635	20
rect	634	20	635	21
rect	634	21	635	22
rect	634	22	635	23
rect	634	23	635	24
rect	634	24	635	25
rect	634	25	635	26
rect	634	26	635	27
rect	634	27	635	28
rect	634	28	635	29
rect	634	29	635	30
rect	634	30	635	31
rect	634	31	635	32
rect	634	32	635	33
rect	634	33	635	34
rect	634	34	635	35
rect	634	35	635	36
rect	634	36	635	37
rect	634	37	635	38
rect	634	38	635	39
rect	634	39	635	40
rect	634	40	635	41
rect	634	41	635	42
rect	634	42	635	43
rect	634	43	635	44
rect	634	44	635	45
rect	634	45	635	46
rect	634	46	635	47
rect	634	47	635	48
rect	634	48	635	49
rect	634	49	635	50
rect	634	50	635	51
rect	634	51	635	52
rect	634	52	635	53
rect	634	53	635	54
rect	634	54	635	55
rect	634	55	635	56
rect	634	56	635	57
rect	634	57	635	58
rect	634	58	635	59
rect	634	59	635	60
rect	634	60	635	61
rect	634	61	635	62
rect	634	62	635	63
rect	634	63	635	64
rect	634	64	635	65
rect	634	65	635	66
rect	634	66	635	67
rect	634	67	635	68
rect	634	68	635	69
rect	634	69	635	70
rect	634	70	635	71
rect	634	71	635	72
rect	634	72	635	73
rect	634	73	635	74
rect	634	74	635	75
rect	634	75	635	76
rect	634	76	635	77
rect	634	77	635	78
rect	634	78	635	79
rect	634	79	635	80
rect	634	80	635	81
rect	634	81	635	82
rect	634	82	635	83
rect	634	83	635	84
rect	634	84	635	85
rect	634	85	635	86
rect	634	86	635	87
rect	634	87	635	88
rect	634	88	635	89
rect	634	89	635	90
rect	634	90	635	91
rect	634	91	635	92
rect	634	92	635	93
rect	634	93	635	94
rect	634	94	635	95
rect	634	95	635	96
rect	634	96	635	97
rect	634	97	635	98
rect	634	98	635	99
rect	634	99	635	100
rect	634	100	635	101
rect	634	101	635	102
rect	634	102	635	103
rect	634	103	635	104
rect	634	104	635	105
rect	634	105	635	106
rect	634	106	635	107
rect	634	107	635	108
rect	634	108	635	109
rect	634	109	635	110
rect	634	110	635	111
rect	634	111	635	112
rect	634	112	635	113
rect	634	113	635	114
rect	634	114	635	115
rect	634	115	635	116
rect	634	116	635	117
rect	634	117	635	118
rect	634	118	635	119
rect	634	119	635	120
rect	634	120	635	121
rect	634	121	635	122
rect	634	122	635	123
rect	634	123	635	124
rect	634	124	635	125
rect	634	125	635	126
rect	634	126	635	127
rect	634	127	635	128
rect	634	128	635	129
rect	634	129	635	130
rect	634	130	635	131
rect	634	131	635	132
rect	634	132	635	133
rect	634	133	635	134
rect	634	134	635	135
rect	634	135	635	136
rect	634	136	635	137
rect	634	137	635	138
rect	634	138	635	139
rect	634	139	635	140
rect	634	140	635	141
rect	634	141	635	142
rect	634	142	635	143
rect	634	143	635	144
rect	634	144	635	145
rect	634	145	635	146
rect	634	146	635	147
rect	634	147	635	148
rect	634	148	635	149
rect	634	149	635	150
rect	634	150	635	151
rect	634	151	635	152
rect	634	152	635	153
rect	634	153	635	154
rect	634	154	635	155
rect	634	155	635	156
rect	634	156	635	157
rect	634	157	635	158
rect	634	158	635	159
rect	634	159	635	160
rect	634	160	635	161
rect	634	161	635	162
rect	634	162	635	163
rect	634	163	635	164
rect	634	164	635	165
rect	634	165	635	166
rect	634	166	635	167
rect	634	167	635	168
rect	634	168	635	169
rect	634	169	635	170
rect	634	170	635	171
rect	634	171	635	172
rect	634	172	635	173
rect	634	173	635	174
rect	634	174	635	175
rect	634	175	635	176
rect	634	176	635	177
rect	634	177	635	178
rect	634	178	635	179
rect	634	179	635	180
rect	634	180	635	181
rect	634	181	635	182
rect	634	182	635	183
rect	634	183	635	184
rect	634	184	635	185
rect	634	185	635	186
rect	634	186	635	187
rect	634	187	635	188
rect	634	188	635	189
rect	634	189	635	190
rect	634	190	635	191
rect	634	191	635	192
rect	634	192	635	193
rect	634	193	635	194
rect	634	194	635	195
rect	634	195	635	196
rect	634	196	635	197
rect	634	197	635	198
rect	634	198	635	199
rect	634	199	635	200
rect	634	200	635	201
rect	634	201	635	202
rect	634	202	635	203
rect	634	203	635	204
rect	634	204	635	205
rect	634	205	635	206
rect	634	206	635	207
rect	634	207	635	208
rect	634	208	635	209
rect	634	209	635	210
rect	634	210	635	211
rect	634	211	635	212
rect	634	212	635	213
rect	634	213	635	214
rect	634	214	635	215
rect	634	215	635	216
rect	634	216	635	217
rect	634	217	635	218
rect	634	218	635	219
rect	648	0	649	1
rect	648	1	649	2
rect	648	2	649	3
rect	648	3	649	4
rect	648	4	649	5
rect	648	5	649	6
rect	648	6	649	7
rect	648	7	649	8
rect	648	8	649	9
rect	648	9	649	10
rect	648	10	649	11
rect	648	11	649	12
rect	648	12	649	13
rect	648	13	649	14
rect	648	14	649	15
rect	648	15	649	16
rect	648	16	649	17
rect	648	17	649	18
rect	648	18	649	19
rect	648	19	649	20
rect	648	20	649	21
rect	648	21	649	22
rect	648	22	649	23
rect	648	23	649	24
rect	648	24	649	25
rect	648	25	649	26
rect	648	26	649	27
rect	648	27	649	28
rect	648	28	649	29
rect	648	29	649	30
rect	648	30	649	31
rect	648	31	649	32
rect	648	32	649	33
rect	648	33	649	34
rect	648	34	649	35
rect	648	35	649	36
rect	648	36	649	37
rect	648	37	649	38
rect	648	38	649	39
rect	648	39	649	40
rect	648	40	649	41
rect	648	41	649	42
rect	648	42	649	43
rect	648	43	649	44
rect	648	44	649	45
rect	648	45	649	46
rect	648	46	649	47
rect	648	47	649	48
rect	648	48	649	49
rect	648	49	649	50
rect	648	50	649	51
rect	648	51	649	52
rect	648	52	649	53
rect	648	53	649	54
rect	648	54	649	55
rect	648	55	649	56
rect	648	56	649	57
rect	648	57	649	58
rect	648	58	649	59
rect	648	59	649	60
rect	648	60	649	61
rect	648	61	649	62
rect	648	62	649	63
rect	648	63	649	64
rect	648	64	649	65
rect	648	65	649	66
rect	648	66	649	67
rect	648	67	649	68
rect	648	68	649	69
rect	648	69	649	70
rect	648	70	649	71
rect	648	71	649	72
rect	648	72	649	73
rect	648	73	649	74
rect	648	74	649	75
rect	648	75	649	76
rect	648	76	649	77
rect	648	77	649	78
rect	648	78	649	79
rect	648	79	649	80
rect	648	80	649	81
rect	648	81	649	82
rect	648	82	649	83
rect	648	83	649	84
rect	648	84	649	85
rect	648	85	649	86
rect	648	86	649	87
rect	648	87	649	88
rect	648	88	649	89
rect	648	89	649	90
rect	648	90	649	91
rect	648	91	649	92
rect	648	92	649	93
rect	648	93	649	94
rect	648	94	649	95
rect	648	95	649	96
rect	648	96	649	97
rect	648	97	649	98
rect	648	98	649	99
rect	648	99	649	100
rect	648	100	649	101
rect	648	101	649	102
rect	648	102	649	103
rect	648	103	649	104
rect	648	104	649	105
rect	648	105	649	106
rect	648	106	649	107
rect	648	107	649	108
rect	648	108	649	109
rect	648	109	649	110
rect	648	110	649	111
rect	648	111	649	112
rect	648	112	649	113
rect	648	113	649	114
rect	648	114	649	115
rect	648	115	649	116
rect	648	116	649	117
rect	648	117	649	118
rect	648	118	649	119
rect	648	119	649	120
rect	648	120	649	121
rect	648	121	649	122
rect	648	122	649	123
rect	648	123	649	124
rect	648	124	649	125
rect	648	125	649	126
rect	648	126	649	127
rect	648	127	649	128
rect	648	128	649	129
rect	648	129	649	130
rect	648	130	649	131
rect	648	131	649	132
rect	648	132	649	133
rect	648	133	649	134
rect	648	134	649	135
rect	648	135	649	136
rect	648	136	649	137
rect	648	137	649	138
rect	648	138	649	139
rect	648	139	649	140
rect	648	140	649	141
rect	648	141	649	142
rect	648	142	649	143
rect	648	143	649	144
rect	648	144	649	145
rect	648	145	649	146
rect	648	146	649	147
rect	648	147	649	148
rect	648	148	649	149
rect	648	149	649	150
rect	648	150	649	151
rect	648	151	649	152
rect	648	152	649	153
rect	648	153	649	154
rect	648	154	649	155
rect	648	155	649	156
rect	648	156	649	157
rect	648	157	649	158
rect	648	158	649	159
rect	648	159	649	160
rect	648	160	649	161
rect	648	161	649	162
rect	648	162	649	163
rect	648	163	649	164
rect	648	164	649	165
rect	648	165	649	166
rect	648	166	649	167
rect	648	167	649	168
rect	648	168	649	169
rect	648	169	649	170
rect	648	170	649	171
rect	648	171	649	172
rect	648	172	649	173
rect	648	173	649	174
rect	648	174	649	175
rect	648	175	649	176
rect	648	176	649	177
rect	648	177	649	178
rect	648	178	649	179
rect	648	179	649	180
rect	648	180	649	181
rect	648	181	649	182
rect	648	182	649	183
rect	648	183	649	184
rect	648	184	649	185
rect	648	185	649	186
rect	648	186	649	187
rect	648	187	649	188
rect	648	188	649	189
rect	648	189	649	190
rect	648	190	649	191
rect	648	191	649	192
rect	648	192	649	193
rect	648	193	649	194
rect	648	194	649	195
rect	649	0	650	1
rect	649	1	650	2
rect	649	2	650	3
rect	649	3	650	4
rect	649	4	650	5
rect	649	5	650	6
rect	649	6	650	7
rect	649	7	650	8
rect	649	8	650	9
rect	649	9	650	10
rect	649	10	650	11
rect	649	11	650	12
rect	649	12	650	13
rect	649	13	650	14
rect	649	14	650	15
rect	649	15	650	16
rect	649	16	650	17
rect	649	17	650	18
rect	649	18	650	19
rect	649	19	650	20
rect	649	20	650	21
rect	649	21	650	22
rect	649	22	650	23
rect	649	23	650	24
rect	649	24	650	25
rect	649	25	650	26
rect	649	26	650	27
rect	649	27	650	28
rect	649	28	650	29
rect	649	29	650	30
rect	649	30	650	31
rect	649	31	650	32
rect	649	32	650	33
rect	649	33	650	34
rect	649	34	650	35
rect	649	35	650	36
rect	649	36	650	37
rect	649	37	650	38
rect	649	38	650	39
rect	649	39	650	40
rect	649	40	650	41
rect	649	41	650	42
rect	649	42	650	43
rect	649	43	650	44
rect	649	44	650	45
rect	649	45	650	46
rect	649	46	650	47
rect	649	47	650	48
rect	649	48	650	49
rect	649	49	650	50
rect	649	50	650	51
rect	649	51	650	52
rect	649	52	650	53
rect	649	53	650	54
rect	649	54	650	55
rect	649	55	650	56
rect	649	56	650	57
rect	649	57	650	58
rect	649	58	650	59
rect	649	59	650	60
rect	649	60	650	61
rect	649	61	650	62
rect	649	62	650	63
rect	649	63	650	64
rect	649	64	650	65
rect	649	65	650	66
rect	649	66	650	67
rect	649	67	650	68
rect	649	68	650	69
rect	649	69	650	70
rect	649	70	650	71
rect	649	71	650	72
rect	649	72	650	73
rect	649	73	650	74
rect	649	74	650	75
rect	649	75	650	76
rect	649	76	650	77
rect	649	77	650	78
rect	649	78	650	79
rect	649	79	650	80
rect	649	80	650	81
rect	649	81	650	82
rect	649	82	650	83
rect	649	83	650	84
rect	649	84	650	85
rect	649	85	650	86
rect	649	86	650	87
rect	649	87	650	88
rect	649	88	650	89
rect	649	89	650	90
rect	649	90	650	91
rect	649	91	650	92
rect	649	92	650	93
rect	649	93	650	94
rect	649	94	650	95
rect	649	95	650	96
rect	649	96	650	97
rect	649	97	650	98
rect	649	98	650	99
rect	649	99	650	100
rect	649	100	650	101
rect	649	101	650	102
rect	649	102	650	103
rect	649	103	650	104
rect	649	104	650	105
rect	649	105	650	106
rect	649	106	650	107
rect	649	107	650	108
rect	649	108	650	109
rect	649	109	650	110
rect	649	110	650	111
rect	649	111	650	112
rect	649	112	650	113
rect	649	113	650	114
rect	649	114	650	115
rect	649	115	650	116
rect	649	116	650	117
rect	649	117	650	118
rect	649	118	650	119
rect	649	119	650	120
rect	649	120	650	121
rect	649	121	650	122
rect	649	122	650	123
rect	649	123	650	124
rect	649	124	650	125
rect	649	125	650	126
rect	649	126	650	127
rect	649	127	650	128
rect	649	128	650	129
rect	649	129	650	130
rect	649	130	650	131
rect	649	131	650	132
rect	649	132	650	133
rect	649	133	650	134
rect	649	134	650	135
rect	649	135	650	136
rect	649	136	650	137
rect	649	137	650	138
rect	649	138	650	139
rect	649	139	650	140
rect	649	140	650	141
rect	649	141	650	142
rect	649	142	650	143
rect	649	143	650	144
rect	649	144	650	145
rect	649	145	650	146
rect	649	146	650	147
rect	649	147	650	148
rect	649	148	650	149
rect	649	149	650	150
rect	649	150	650	151
rect	649	151	650	152
rect	649	152	650	153
rect	649	153	650	154
rect	649	154	650	155
rect	649	155	650	156
rect	649	156	650	157
rect	649	157	650	158
rect	649	158	650	159
rect	649	159	650	160
rect	649	160	650	161
rect	649	161	650	162
rect	649	162	650	163
rect	649	163	650	164
rect	649	164	650	165
rect	649	165	650	166
rect	649	166	650	167
rect	649	167	650	168
rect	649	168	650	169
rect	649	169	650	170
rect	649	170	650	171
rect	649	171	650	172
rect	649	172	650	173
rect	649	173	650	174
rect	649	174	650	175
rect	649	175	650	176
rect	649	176	650	177
rect	649	177	650	178
rect	649	178	650	179
rect	649	179	650	180
rect	649	180	650	181
rect	649	181	650	182
rect	649	182	650	183
rect	649	183	650	184
rect	649	184	650	185
rect	649	185	650	186
rect	649	186	650	187
rect	649	187	650	188
rect	649	188	650	189
rect	649	189	650	190
rect	649	190	650	191
rect	649	191	650	192
rect	649	192	650	193
rect	649	193	650	194
rect	649	194	650	195
rect	650	0	651	1
rect	650	1	651	2
rect	650	2	651	3
rect	650	3	651	4
rect	650	4	651	5
rect	650	5	651	6
rect	650	6	651	7
rect	650	7	651	8
rect	650	8	651	9
rect	650	9	651	10
rect	650	10	651	11
rect	650	11	651	12
rect	650	12	651	13
rect	650	13	651	14
rect	650	14	651	15
rect	650	15	651	16
rect	650	16	651	17
rect	650	17	651	18
rect	650	18	651	19
rect	650	19	651	20
rect	650	20	651	21
rect	650	21	651	22
rect	650	22	651	23
rect	650	23	651	24
rect	650	24	651	25
rect	650	25	651	26
rect	650	26	651	27
rect	650	27	651	28
rect	650	28	651	29
rect	650	29	651	30
rect	650	30	651	31
rect	650	31	651	32
rect	650	32	651	33
rect	650	33	651	34
rect	650	34	651	35
rect	650	35	651	36
rect	650	36	651	37
rect	650	37	651	38
rect	650	38	651	39
rect	650	39	651	40
rect	650	40	651	41
rect	650	41	651	42
rect	650	42	651	43
rect	650	43	651	44
rect	650	44	651	45
rect	650	45	651	46
rect	650	46	651	47
rect	650	47	651	48
rect	650	48	651	49
rect	650	49	651	50
rect	650	50	651	51
rect	650	51	651	52
rect	650	52	651	53
rect	650	53	651	54
rect	650	54	651	55
rect	650	55	651	56
rect	650	56	651	57
rect	650	57	651	58
rect	650	58	651	59
rect	650	59	651	60
rect	650	60	651	61
rect	650	61	651	62
rect	650	62	651	63
rect	650	63	651	64
rect	650	64	651	65
rect	650	65	651	66
rect	650	66	651	67
rect	650	67	651	68
rect	650	68	651	69
rect	650	69	651	70
rect	650	70	651	71
rect	650	71	651	72
rect	650	72	651	73
rect	650	73	651	74
rect	650	74	651	75
rect	650	75	651	76
rect	650	76	651	77
rect	650	77	651	78
rect	650	78	651	79
rect	650	79	651	80
rect	650	80	651	81
rect	650	81	651	82
rect	650	82	651	83
rect	650	83	651	84
rect	650	84	651	85
rect	650	85	651	86
rect	650	86	651	87
rect	650	87	651	88
rect	650	88	651	89
rect	650	89	651	90
rect	650	90	651	91
rect	650	91	651	92
rect	650	92	651	93
rect	650	93	651	94
rect	650	94	651	95
rect	650	95	651	96
rect	650	96	651	97
rect	650	97	651	98
rect	650	98	651	99
rect	650	99	651	100
rect	650	100	651	101
rect	650	101	651	102
rect	650	102	651	103
rect	650	103	651	104
rect	650	104	651	105
rect	650	105	651	106
rect	650	106	651	107
rect	650	107	651	108
rect	650	108	651	109
rect	650	109	651	110
rect	650	110	651	111
rect	650	111	651	112
rect	650	112	651	113
rect	650	113	651	114
rect	650	114	651	115
rect	650	115	651	116
rect	650	116	651	117
rect	650	117	651	118
rect	650	118	651	119
rect	650	119	651	120
rect	650	120	651	121
rect	650	121	651	122
rect	650	122	651	123
rect	650	123	651	124
rect	650	124	651	125
rect	650	125	651	126
rect	650	126	651	127
rect	650	127	651	128
rect	650	128	651	129
rect	650	129	651	130
rect	650	130	651	131
rect	650	131	651	132
rect	650	132	651	133
rect	650	133	651	134
rect	650	134	651	135
rect	650	135	651	136
rect	650	136	651	137
rect	650	137	651	138
rect	650	138	651	139
rect	650	139	651	140
rect	650	140	651	141
rect	650	141	651	142
rect	650	142	651	143
rect	650	143	651	144
rect	650	144	651	145
rect	650	145	651	146
rect	650	146	651	147
rect	650	147	651	148
rect	650	148	651	149
rect	650	149	651	150
rect	650	150	651	151
rect	650	151	651	152
rect	650	152	651	153
rect	650	153	651	154
rect	650	154	651	155
rect	650	155	651	156
rect	650	156	651	157
rect	650	157	651	158
rect	650	158	651	159
rect	650	159	651	160
rect	650	160	651	161
rect	650	161	651	162
rect	650	162	651	163
rect	650	163	651	164
rect	650	164	651	165
rect	650	165	651	166
rect	650	166	651	167
rect	650	167	651	168
rect	650	168	651	169
rect	650	169	651	170
rect	650	170	651	171
rect	650	171	651	172
rect	650	172	651	173
rect	650	173	651	174
rect	650	174	651	175
rect	650	175	651	176
rect	650	176	651	177
rect	650	177	651	178
rect	650	178	651	179
rect	650	179	651	180
rect	650	180	651	181
rect	650	181	651	182
rect	650	182	651	183
rect	650	183	651	184
rect	650	184	651	185
rect	650	185	651	186
rect	650	186	651	187
rect	650	187	651	188
rect	650	188	651	189
rect	650	189	651	190
rect	650	190	651	191
rect	650	191	651	192
rect	650	192	651	193
rect	650	193	651	194
rect	650	194	651	195
rect	651	0	652	1
rect	651	1	652	2
rect	651	2	652	3
rect	651	3	652	4
rect	651	4	652	5
rect	651	5	652	6
rect	651	6	652	7
rect	651	7	652	8
rect	651	8	652	9
rect	651	9	652	10
rect	651	10	652	11
rect	651	11	652	12
rect	651	12	652	13
rect	651	13	652	14
rect	651	14	652	15
rect	651	15	652	16
rect	651	16	652	17
rect	651	17	652	18
rect	651	18	652	19
rect	651	19	652	20
rect	651	20	652	21
rect	651	21	652	22
rect	651	22	652	23
rect	651	23	652	24
rect	651	24	652	25
rect	651	25	652	26
rect	651	26	652	27
rect	651	27	652	28
rect	651	28	652	29
rect	651	29	652	30
rect	651	30	652	31
rect	651	31	652	32
rect	651	32	652	33
rect	651	33	652	34
rect	651	34	652	35
rect	651	35	652	36
rect	651	36	652	37
rect	651	37	652	38
rect	651	38	652	39
rect	651	39	652	40
rect	651	40	652	41
rect	651	41	652	42
rect	651	42	652	43
rect	651	43	652	44
rect	651	44	652	45
rect	651	45	652	46
rect	651	46	652	47
rect	651	47	652	48
rect	651	48	652	49
rect	651	49	652	50
rect	651	50	652	51
rect	651	51	652	52
rect	651	52	652	53
rect	651	53	652	54
rect	651	54	652	55
rect	651	55	652	56
rect	651	56	652	57
rect	651	57	652	58
rect	651	58	652	59
rect	651	59	652	60
rect	651	60	652	61
rect	651	61	652	62
rect	651	62	652	63
rect	651	63	652	64
rect	651	64	652	65
rect	651	65	652	66
rect	651	66	652	67
rect	651	67	652	68
rect	651	68	652	69
rect	651	69	652	70
rect	651	70	652	71
rect	651	71	652	72
rect	651	72	652	73
rect	651	73	652	74
rect	651	74	652	75
rect	651	75	652	76
rect	651	76	652	77
rect	651	77	652	78
rect	651	78	652	79
rect	651	79	652	80
rect	651	80	652	81
rect	651	81	652	82
rect	651	82	652	83
rect	651	83	652	84
rect	651	84	652	85
rect	651	85	652	86
rect	651	86	652	87
rect	651	87	652	88
rect	651	88	652	89
rect	651	89	652	90
rect	651	90	652	91
rect	651	91	652	92
rect	651	92	652	93
rect	651	93	652	94
rect	651	94	652	95
rect	651	95	652	96
rect	651	96	652	97
rect	651	97	652	98
rect	651	98	652	99
rect	651	99	652	100
rect	651	100	652	101
rect	651	101	652	102
rect	651	102	652	103
rect	651	103	652	104
rect	651	104	652	105
rect	651	105	652	106
rect	651	106	652	107
rect	651	107	652	108
rect	651	108	652	109
rect	651	109	652	110
rect	651	110	652	111
rect	651	111	652	112
rect	651	112	652	113
rect	651	113	652	114
rect	651	114	652	115
rect	651	115	652	116
rect	651	116	652	117
rect	651	117	652	118
rect	651	118	652	119
rect	651	119	652	120
rect	651	120	652	121
rect	651	121	652	122
rect	651	122	652	123
rect	651	123	652	124
rect	651	124	652	125
rect	651	125	652	126
rect	651	126	652	127
rect	651	127	652	128
rect	651	128	652	129
rect	651	129	652	130
rect	651	130	652	131
rect	651	131	652	132
rect	651	132	652	133
rect	651	133	652	134
rect	651	134	652	135
rect	651	135	652	136
rect	651	136	652	137
rect	651	137	652	138
rect	651	138	652	139
rect	651	139	652	140
rect	651	140	652	141
rect	651	141	652	142
rect	651	142	652	143
rect	651	143	652	144
rect	651	144	652	145
rect	651	145	652	146
rect	651	146	652	147
rect	651	147	652	148
rect	651	148	652	149
rect	651	149	652	150
rect	651	150	652	151
rect	651	151	652	152
rect	651	152	652	153
rect	651	153	652	154
rect	651	154	652	155
rect	651	155	652	156
rect	651	156	652	157
rect	651	157	652	158
rect	651	158	652	159
rect	651	159	652	160
rect	651	160	652	161
rect	651	161	652	162
rect	651	162	652	163
rect	651	163	652	164
rect	651	164	652	165
rect	651	165	652	166
rect	651	166	652	167
rect	651	167	652	168
rect	651	168	652	169
rect	651	169	652	170
rect	651	170	652	171
rect	651	171	652	172
rect	651	172	652	173
rect	651	173	652	174
rect	651	174	652	175
rect	651	175	652	176
rect	651	176	652	177
rect	651	177	652	178
rect	651	178	652	179
rect	651	179	652	180
rect	651	180	652	181
rect	651	181	652	182
rect	651	182	652	183
rect	651	183	652	184
rect	651	184	652	185
rect	651	185	652	186
rect	651	186	652	187
rect	651	187	652	188
rect	651	188	652	189
rect	651	189	652	190
rect	651	190	652	191
rect	651	191	652	192
rect	651	192	652	193
rect	651	193	652	194
rect	651	194	652	195
rect	652	0	653	1
rect	652	1	653	2
rect	652	2	653	3
rect	652	3	653	4
rect	652	4	653	5
rect	652	5	653	6
rect	652	6	653	7
rect	652	7	653	8
rect	652	8	653	9
rect	652	9	653	10
rect	652	10	653	11
rect	652	11	653	12
rect	652	12	653	13
rect	652	13	653	14
rect	652	14	653	15
rect	652	15	653	16
rect	652	16	653	17
rect	652	17	653	18
rect	652	18	653	19
rect	652	19	653	20
rect	652	20	653	21
rect	652	21	653	22
rect	652	22	653	23
rect	652	23	653	24
rect	652	24	653	25
rect	652	25	653	26
rect	652	26	653	27
rect	652	27	653	28
rect	652	28	653	29
rect	652	29	653	30
rect	652	30	653	31
rect	652	31	653	32
rect	652	32	653	33
rect	652	33	653	34
rect	652	34	653	35
rect	652	35	653	36
rect	652	36	653	37
rect	652	37	653	38
rect	652	38	653	39
rect	652	39	653	40
rect	652	40	653	41
rect	652	41	653	42
rect	652	42	653	43
rect	652	43	653	44
rect	652	44	653	45
rect	652	45	653	46
rect	652	46	653	47
rect	652	47	653	48
rect	652	48	653	49
rect	652	49	653	50
rect	652	50	653	51
rect	652	51	653	52
rect	652	52	653	53
rect	652	53	653	54
rect	652	54	653	55
rect	652	55	653	56
rect	652	56	653	57
rect	652	57	653	58
rect	652	58	653	59
rect	652	59	653	60
rect	652	60	653	61
rect	652	61	653	62
rect	652	62	653	63
rect	652	63	653	64
rect	652	64	653	65
rect	652	65	653	66
rect	652	66	653	67
rect	652	67	653	68
rect	652	68	653	69
rect	652	69	653	70
rect	652	70	653	71
rect	652	71	653	72
rect	652	72	653	73
rect	652	73	653	74
rect	652	74	653	75
rect	652	75	653	76
rect	652	76	653	77
rect	652	77	653	78
rect	652	78	653	79
rect	652	79	653	80
rect	652	80	653	81
rect	652	81	653	82
rect	652	82	653	83
rect	652	83	653	84
rect	652	84	653	85
rect	652	85	653	86
rect	652	86	653	87
rect	652	87	653	88
rect	652	88	653	89
rect	652	89	653	90
rect	652	90	653	91
rect	652	91	653	92
rect	652	92	653	93
rect	652	93	653	94
rect	652	94	653	95
rect	652	95	653	96
rect	652	96	653	97
rect	652	97	653	98
rect	652	98	653	99
rect	652	99	653	100
rect	652	100	653	101
rect	652	101	653	102
rect	652	102	653	103
rect	652	103	653	104
rect	652	104	653	105
rect	652	105	653	106
rect	652	106	653	107
rect	652	107	653	108
rect	652	108	653	109
rect	652	109	653	110
rect	652	110	653	111
rect	652	111	653	112
rect	652	112	653	113
rect	652	113	653	114
rect	652	114	653	115
rect	652	115	653	116
rect	652	116	653	117
rect	652	117	653	118
rect	652	118	653	119
rect	652	119	653	120
rect	652	120	653	121
rect	652	121	653	122
rect	652	122	653	123
rect	652	123	653	124
rect	652	124	653	125
rect	652	125	653	126
rect	652	126	653	127
rect	652	127	653	128
rect	652	128	653	129
rect	652	129	653	130
rect	652	130	653	131
rect	652	131	653	132
rect	652	132	653	133
rect	652	133	653	134
rect	652	134	653	135
rect	652	135	653	136
rect	652	136	653	137
rect	652	137	653	138
rect	652	138	653	139
rect	652	139	653	140
rect	652	140	653	141
rect	652	141	653	142
rect	652	142	653	143
rect	652	143	653	144
rect	652	144	653	145
rect	652	145	653	146
rect	652	146	653	147
rect	652	147	653	148
rect	652	148	653	149
rect	652	149	653	150
rect	652	150	653	151
rect	652	151	653	152
rect	652	152	653	153
rect	652	153	653	154
rect	652	154	653	155
rect	652	155	653	156
rect	652	156	653	157
rect	652	157	653	158
rect	652	158	653	159
rect	652	159	653	160
rect	652	160	653	161
rect	652	161	653	162
rect	652	162	653	163
rect	652	163	653	164
rect	652	164	653	165
rect	652	165	653	166
rect	652	166	653	167
rect	652	167	653	168
rect	652	168	653	169
rect	652	169	653	170
rect	652	170	653	171
rect	652	171	653	172
rect	652	172	653	173
rect	652	173	653	174
rect	652	174	653	175
rect	652	175	653	176
rect	652	176	653	177
rect	652	177	653	178
rect	652	178	653	179
rect	652	179	653	180
rect	652	180	653	181
rect	652	181	653	182
rect	652	182	653	183
rect	652	183	653	184
rect	652	184	653	185
rect	652	185	653	186
rect	652	186	653	187
rect	652	187	653	188
rect	652	188	653	189
rect	652	189	653	190
rect	652	190	653	191
rect	652	191	653	192
rect	652	192	653	193
rect	652	193	653	194
rect	652	194	653	195
rect	653	0	654	1
rect	653	1	654	2
rect	653	2	654	3
rect	653	3	654	4
rect	653	4	654	5
rect	653	5	654	6
rect	653	6	654	7
rect	653	7	654	8
rect	653	8	654	9
rect	653	9	654	10
rect	653	10	654	11
rect	653	11	654	12
rect	653	12	654	13
rect	653	13	654	14
rect	653	14	654	15
rect	653	15	654	16
rect	653	16	654	17
rect	653	17	654	18
rect	653	18	654	19
rect	653	19	654	20
rect	653	20	654	21
rect	653	21	654	22
rect	653	22	654	23
rect	653	23	654	24
rect	653	24	654	25
rect	653	25	654	26
rect	653	26	654	27
rect	653	27	654	28
rect	653	28	654	29
rect	653	29	654	30
rect	653	30	654	31
rect	653	31	654	32
rect	653	32	654	33
rect	653	33	654	34
rect	653	34	654	35
rect	653	35	654	36
rect	653	36	654	37
rect	653	37	654	38
rect	653	38	654	39
rect	653	39	654	40
rect	653	40	654	41
rect	653	41	654	42
rect	653	42	654	43
rect	653	43	654	44
rect	653	44	654	45
rect	653	45	654	46
rect	653	46	654	47
rect	653	47	654	48
rect	653	48	654	49
rect	653	49	654	50
rect	653	50	654	51
rect	653	51	654	52
rect	653	52	654	53
rect	653	53	654	54
rect	653	54	654	55
rect	653	55	654	56
rect	653	56	654	57
rect	653	57	654	58
rect	653	58	654	59
rect	653	59	654	60
rect	653	60	654	61
rect	653	61	654	62
rect	653	62	654	63
rect	653	63	654	64
rect	653	64	654	65
rect	653	65	654	66
rect	653	66	654	67
rect	653	67	654	68
rect	653	68	654	69
rect	653	69	654	70
rect	653	70	654	71
rect	653	71	654	72
rect	653	72	654	73
rect	653	73	654	74
rect	653	74	654	75
rect	653	75	654	76
rect	653	76	654	77
rect	653	77	654	78
rect	653	78	654	79
rect	653	79	654	80
rect	653	80	654	81
rect	653	81	654	82
rect	653	82	654	83
rect	653	83	654	84
rect	653	84	654	85
rect	653	85	654	86
rect	653	86	654	87
rect	653	87	654	88
rect	653	88	654	89
rect	653	89	654	90
rect	653	90	654	91
rect	653	91	654	92
rect	653	92	654	93
rect	653	93	654	94
rect	653	94	654	95
rect	653	95	654	96
rect	653	96	654	97
rect	653	97	654	98
rect	653	98	654	99
rect	653	99	654	100
rect	653	100	654	101
rect	653	101	654	102
rect	653	102	654	103
rect	653	103	654	104
rect	653	104	654	105
rect	653	105	654	106
rect	653	106	654	107
rect	653	107	654	108
rect	653	108	654	109
rect	653	109	654	110
rect	653	110	654	111
rect	653	111	654	112
rect	653	112	654	113
rect	653	113	654	114
rect	653	114	654	115
rect	653	115	654	116
rect	653	116	654	117
rect	653	117	654	118
rect	653	118	654	119
rect	653	119	654	120
rect	653	120	654	121
rect	653	121	654	122
rect	653	122	654	123
rect	653	123	654	124
rect	653	124	654	125
rect	653	125	654	126
rect	653	126	654	127
rect	653	127	654	128
rect	653	128	654	129
rect	653	129	654	130
rect	653	130	654	131
rect	653	131	654	132
rect	653	132	654	133
rect	653	133	654	134
rect	653	134	654	135
rect	653	135	654	136
rect	653	136	654	137
rect	653	137	654	138
rect	653	138	654	139
rect	653	139	654	140
rect	653	140	654	141
rect	653	141	654	142
rect	653	142	654	143
rect	653	143	654	144
rect	653	144	654	145
rect	653	145	654	146
rect	653	146	654	147
rect	653	147	654	148
rect	653	148	654	149
rect	653	149	654	150
rect	653	150	654	151
rect	653	151	654	152
rect	653	152	654	153
rect	653	153	654	154
rect	653	154	654	155
rect	653	155	654	156
rect	653	156	654	157
rect	653	157	654	158
rect	653	158	654	159
rect	653	159	654	160
rect	653	160	654	161
rect	653	161	654	162
rect	653	162	654	163
rect	653	163	654	164
rect	653	164	654	165
rect	653	165	654	166
rect	653	166	654	167
rect	653	167	654	168
rect	653	168	654	169
rect	653	169	654	170
rect	653	170	654	171
rect	653	171	654	172
rect	653	172	654	173
rect	653	173	654	174
rect	653	174	654	175
rect	653	175	654	176
rect	653	176	654	177
rect	653	177	654	178
rect	653	178	654	179
rect	653	179	654	180
rect	653	180	654	181
rect	653	181	654	182
rect	653	182	654	183
rect	653	183	654	184
rect	653	184	654	185
rect	653	185	654	186
rect	653	186	654	187
rect	653	187	654	188
rect	653	188	654	189
rect	653	189	654	190
rect	653	190	654	191
rect	653	191	654	192
rect	653	192	654	193
rect	653	193	654	194
rect	653	194	654	195
rect	661	0	662	1
rect	661	1	662	2
rect	661	2	662	3
rect	661	3	662	4
rect	661	4	662	5
rect	661	5	662	6
rect	661	6	662	7
rect	661	7	662	8
rect	661	8	662	9
rect	661	9	662	10
rect	661	10	662	11
rect	661	11	662	12
rect	661	12	662	13
rect	661	13	662	14
rect	661	14	662	15
rect	661	15	662	16
rect	661	16	662	17
rect	661	17	662	18
rect	661	18	662	19
rect	661	19	662	20
rect	661	20	662	21
rect	661	21	662	22
rect	661	22	662	23
rect	661	23	662	24
rect	661	24	662	25
rect	661	25	662	26
rect	661	26	662	27
rect	661	27	662	28
rect	661	28	662	29
rect	661	29	662	30
rect	661	30	662	31
rect	661	31	662	32
rect	661	32	662	33
rect	661	33	662	34
rect	661	34	662	35
rect	661	35	662	36
rect	661	36	662	37
rect	661	37	662	38
rect	661	38	662	39
rect	661	39	662	40
rect	661	40	662	41
rect	661	41	662	42
rect	661	42	662	43
rect	661	43	662	44
rect	661	44	662	45
rect	661	45	662	46
rect	661	46	662	47
rect	661	47	662	48
rect	661	48	662	49
rect	661	49	662	50
rect	661	50	662	51
rect	661	51	662	52
rect	661	52	662	53
rect	661	53	662	54
rect	661	54	662	55
rect	661	55	662	56
rect	661	56	662	57
rect	661	57	662	58
rect	661	58	662	59
rect	661	59	662	60
rect	661	60	662	61
rect	661	61	662	62
rect	661	62	662	63
rect	661	63	662	64
rect	661	64	662	65
rect	661	65	662	66
rect	661	66	662	67
rect	661	67	662	68
rect	661	68	662	69
rect	661	69	662	70
rect	661	70	662	71
rect	661	71	662	72
rect	661	72	662	73
rect	661	73	662	74
rect	661	74	662	75
rect	661	75	662	76
rect	661	76	662	77
rect	661	77	662	78
rect	661	78	662	79
rect	661	79	662	80
rect	661	80	662	81
rect	661	81	662	82
rect	661	82	662	83
rect	661	83	662	84
rect	661	84	662	85
rect	661	85	662	86
rect	661	86	662	87
rect	661	87	662	88
rect	661	88	662	89
rect	661	89	662	90
rect	661	90	662	91
rect	661	91	662	92
rect	661	92	662	93
rect	661	93	662	94
rect	661	94	662	95
rect	661	95	662	96
rect	661	96	662	97
rect	661	97	662	98
rect	661	98	662	99
rect	661	99	662	100
rect	661	100	662	101
rect	661	101	662	102
rect	661	102	662	103
rect	661	103	662	104
rect	661	104	662	105
rect	661	105	662	106
rect	661	106	662	107
rect	661	107	662	108
rect	661	108	662	109
rect	661	109	662	110
rect	661	110	662	111
rect	661	111	662	112
rect	661	112	662	113
rect	661	113	662	114
rect	661	114	662	115
rect	661	115	662	116
rect	661	116	662	117
rect	661	117	662	118
rect	661	118	662	119
rect	661	119	662	120
rect	661	120	662	121
rect	661	121	662	122
rect	661	122	662	123
rect	661	123	662	124
rect	661	124	662	125
rect	661	125	662	126
rect	661	126	662	127
rect	661	127	662	128
rect	661	128	662	129
rect	661	129	662	130
rect	661	130	662	131
rect	661	131	662	132
rect	661	132	662	133
rect	661	133	662	134
rect	661	134	662	135
rect	661	135	662	136
rect	661	136	662	137
rect	661	137	662	138
rect	661	138	662	139
rect	661	139	662	140
rect	661	140	662	141
rect	661	141	662	142
rect	661	142	662	143
rect	661	143	662	144
rect	661	144	662	145
rect	661	145	662	146
rect	661	146	662	147
rect	661	147	662	148
rect	661	148	662	149
rect	661	149	662	150
rect	661	150	662	151
rect	661	151	662	152
rect	661	152	662	153
rect	661	153	662	154
rect	661	154	662	155
rect	661	155	662	156
rect	661	156	662	157
rect	661	157	662	158
rect	661	158	662	159
rect	661	159	662	160
rect	661	160	662	161
rect	661	161	662	162
rect	661	162	662	163
rect	661	163	662	164
rect	661	164	662	165
rect	661	165	662	166
rect	661	166	662	167
rect	661	167	662	168
rect	662	0	663	1
rect	662	1	663	2
rect	662	2	663	3
rect	662	3	663	4
rect	662	4	663	5
rect	662	5	663	6
rect	662	6	663	7
rect	662	7	663	8
rect	662	8	663	9
rect	662	9	663	10
rect	662	10	663	11
rect	662	11	663	12
rect	662	12	663	13
rect	662	13	663	14
rect	662	14	663	15
rect	662	15	663	16
rect	662	16	663	17
rect	662	17	663	18
rect	662	18	663	19
rect	662	19	663	20
rect	662	20	663	21
rect	662	21	663	22
rect	662	22	663	23
rect	662	23	663	24
rect	662	24	663	25
rect	662	25	663	26
rect	662	26	663	27
rect	662	27	663	28
rect	662	28	663	29
rect	662	29	663	30
rect	662	30	663	31
rect	662	31	663	32
rect	662	32	663	33
rect	662	33	663	34
rect	662	34	663	35
rect	662	35	663	36
rect	662	36	663	37
rect	662	37	663	38
rect	662	38	663	39
rect	662	39	663	40
rect	662	40	663	41
rect	662	41	663	42
rect	662	42	663	43
rect	662	43	663	44
rect	662	44	663	45
rect	662	45	663	46
rect	662	46	663	47
rect	662	47	663	48
rect	662	48	663	49
rect	662	49	663	50
rect	662	50	663	51
rect	662	51	663	52
rect	662	52	663	53
rect	662	53	663	54
rect	662	54	663	55
rect	662	55	663	56
rect	662	56	663	57
rect	662	57	663	58
rect	662	58	663	59
rect	662	59	663	60
rect	662	60	663	61
rect	662	61	663	62
rect	662	62	663	63
rect	662	63	663	64
rect	662	64	663	65
rect	662	65	663	66
rect	662	66	663	67
rect	662	67	663	68
rect	662	68	663	69
rect	662	69	663	70
rect	662	70	663	71
rect	662	71	663	72
rect	662	72	663	73
rect	662	73	663	74
rect	662	74	663	75
rect	662	75	663	76
rect	662	76	663	77
rect	662	77	663	78
rect	662	78	663	79
rect	662	79	663	80
rect	662	80	663	81
rect	662	81	663	82
rect	662	82	663	83
rect	662	83	663	84
rect	662	84	663	85
rect	662	85	663	86
rect	662	86	663	87
rect	662	87	663	88
rect	662	88	663	89
rect	662	89	663	90
rect	662	90	663	91
rect	662	91	663	92
rect	662	92	663	93
rect	662	93	663	94
rect	662	94	663	95
rect	662	95	663	96
rect	662	96	663	97
rect	662	97	663	98
rect	662	98	663	99
rect	662	99	663	100
rect	662	100	663	101
rect	662	101	663	102
rect	662	102	663	103
rect	662	103	663	104
rect	662	104	663	105
rect	662	105	663	106
rect	662	106	663	107
rect	662	107	663	108
rect	662	108	663	109
rect	662	109	663	110
rect	662	110	663	111
rect	662	111	663	112
rect	662	112	663	113
rect	662	113	663	114
rect	662	114	663	115
rect	662	115	663	116
rect	662	116	663	117
rect	662	117	663	118
rect	662	118	663	119
rect	662	119	663	120
rect	662	120	663	121
rect	662	121	663	122
rect	662	122	663	123
rect	662	123	663	124
rect	662	124	663	125
rect	662	125	663	126
rect	662	126	663	127
rect	662	127	663	128
rect	662	128	663	129
rect	662	129	663	130
rect	662	130	663	131
rect	662	131	663	132
rect	662	132	663	133
rect	662	133	663	134
rect	662	134	663	135
rect	662	135	663	136
rect	662	136	663	137
rect	662	137	663	138
rect	662	138	663	139
rect	662	139	663	140
rect	662	140	663	141
rect	662	141	663	142
rect	662	142	663	143
rect	662	143	663	144
rect	662	144	663	145
rect	662	145	663	146
rect	662	146	663	147
rect	662	147	663	148
rect	662	148	663	149
rect	662	149	663	150
rect	662	150	663	151
rect	662	151	663	152
rect	662	152	663	153
rect	662	153	663	154
rect	662	154	663	155
rect	662	155	663	156
rect	662	156	663	157
rect	662	157	663	158
rect	662	158	663	159
rect	662	159	663	160
rect	662	160	663	161
rect	662	161	663	162
rect	662	162	663	163
rect	662	163	663	164
rect	662	164	663	165
rect	662	165	663	166
rect	662	166	663	167
rect	662	167	663	168
rect	663	0	664	1
rect	663	1	664	2
rect	663	2	664	3
rect	663	3	664	4
rect	663	4	664	5
rect	663	5	664	6
rect	663	6	664	7
rect	663	7	664	8
rect	663	8	664	9
rect	663	9	664	10
rect	663	10	664	11
rect	663	11	664	12
rect	663	12	664	13
rect	663	13	664	14
rect	663	14	664	15
rect	663	15	664	16
rect	663	16	664	17
rect	663	17	664	18
rect	663	18	664	19
rect	663	19	664	20
rect	663	20	664	21
rect	663	21	664	22
rect	663	22	664	23
rect	663	23	664	24
rect	663	24	664	25
rect	663	25	664	26
rect	663	26	664	27
rect	663	27	664	28
rect	663	28	664	29
rect	663	29	664	30
rect	663	30	664	31
rect	663	31	664	32
rect	663	32	664	33
rect	663	33	664	34
rect	663	34	664	35
rect	663	35	664	36
rect	663	36	664	37
rect	663	37	664	38
rect	663	38	664	39
rect	663	39	664	40
rect	663	40	664	41
rect	663	41	664	42
rect	663	42	664	43
rect	663	43	664	44
rect	663	44	664	45
rect	663	45	664	46
rect	663	46	664	47
rect	663	47	664	48
rect	663	48	664	49
rect	663	49	664	50
rect	663	50	664	51
rect	663	51	664	52
rect	663	52	664	53
rect	663	53	664	54
rect	663	54	664	55
rect	663	55	664	56
rect	663	56	664	57
rect	663	57	664	58
rect	663	58	664	59
rect	663	59	664	60
rect	663	60	664	61
rect	663	61	664	62
rect	663	62	664	63
rect	663	63	664	64
rect	663	64	664	65
rect	663	65	664	66
rect	663	66	664	67
rect	663	67	664	68
rect	663	68	664	69
rect	663	69	664	70
rect	663	70	664	71
rect	663	71	664	72
rect	663	72	664	73
rect	663	73	664	74
rect	663	74	664	75
rect	663	75	664	76
rect	663	76	664	77
rect	663	77	664	78
rect	663	78	664	79
rect	663	79	664	80
rect	663	80	664	81
rect	663	81	664	82
rect	663	82	664	83
rect	663	83	664	84
rect	663	84	664	85
rect	663	85	664	86
rect	663	86	664	87
rect	663	87	664	88
rect	663	88	664	89
rect	663	89	664	90
rect	663	90	664	91
rect	663	91	664	92
rect	663	92	664	93
rect	663	93	664	94
rect	663	94	664	95
rect	663	95	664	96
rect	663	96	664	97
rect	663	97	664	98
rect	663	98	664	99
rect	663	99	664	100
rect	663	100	664	101
rect	663	101	664	102
rect	663	102	664	103
rect	663	103	664	104
rect	663	104	664	105
rect	663	105	664	106
rect	663	106	664	107
rect	663	107	664	108
rect	663	108	664	109
rect	663	109	664	110
rect	663	110	664	111
rect	663	111	664	112
rect	663	112	664	113
rect	663	113	664	114
rect	663	114	664	115
rect	663	115	664	116
rect	663	116	664	117
rect	663	117	664	118
rect	663	118	664	119
rect	663	119	664	120
rect	663	120	664	121
rect	663	121	664	122
rect	663	122	664	123
rect	663	123	664	124
rect	663	124	664	125
rect	663	125	664	126
rect	663	126	664	127
rect	663	127	664	128
rect	663	128	664	129
rect	663	129	664	130
rect	663	130	664	131
rect	663	131	664	132
rect	663	132	664	133
rect	663	133	664	134
rect	663	134	664	135
rect	663	135	664	136
rect	663	136	664	137
rect	663	137	664	138
rect	663	138	664	139
rect	663	139	664	140
rect	663	140	664	141
rect	663	141	664	142
rect	663	142	664	143
rect	663	143	664	144
rect	663	144	664	145
rect	663	145	664	146
rect	663	146	664	147
rect	663	147	664	148
rect	663	148	664	149
rect	663	149	664	150
rect	663	150	664	151
rect	663	151	664	152
rect	663	152	664	153
rect	663	153	664	154
rect	663	154	664	155
rect	663	155	664	156
rect	663	156	664	157
rect	663	157	664	158
rect	663	158	664	159
rect	663	159	664	160
rect	663	160	664	161
rect	663	161	664	162
rect	663	162	664	163
rect	663	163	664	164
rect	663	164	664	165
rect	663	165	664	166
rect	663	166	664	167
rect	663	167	664	168
rect	664	0	665	1
rect	664	1	665	2
rect	664	2	665	3
rect	664	3	665	4
rect	664	4	665	5
rect	664	5	665	6
rect	664	6	665	7
rect	664	7	665	8
rect	664	8	665	9
rect	664	9	665	10
rect	664	10	665	11
rect	664	11	665	12
rect	664	12	665	13
rect	664	13	665	14
rect	664	14	665	15
rect	664	15	665	16
rect	664	16	665	17
rect	664	17	665	18
rect	664	18	665	19
rect	664	19	665	20
rect	664	20	665	21
rect	664	21	665	22
rect	664	22	665	23
rect	664	23	665	24
rect	664	24	665	25
rect	664	25	665	26
rect	664	26	665	27
rect	664	27	665	28
rect	664	28	665	29
rect	664	29	665	30
rect	664	30	665	31
rect	664	31	665	32
rect	664	32	665	33
rect	664	33	665	34
rect	664	34	665	35
rect	664	35	665	36
rect	664	36	665	37
rect	664	37	665	38
rect	664	38	665	39
rect	664	39	665	40
rect	664	40	665	41
rect	664	41	665	42
rect	664	42	665	43
rect	664	43	665	44
rect	664	44	665	45
rect	664	45	665	46
rect	664	46	665	47
rect	664	47	665	48
rect	664	48	665	49
rect	664	49	665	50
rect	664	50	665	51
rect	664	51	665	52
rect	664	52	665	53
rect	664	53	665	54
rect	664	54	665	55
rect	664	55	665	56
rect	664	56	665	57
rect	664	57	665	58
rect	664	58	665	59
rect	664	59	665	60
rect	664	60	665	61
rect	664	61	665	62
rect	664	62	665	63
rect	664	63	665	64
rect	664	64	665	65
rect	664	65	665	66
rect	664	66	665	67
rect	664	67	665	68
rect	664	68	665	69
rect	664	69	665	70
rect	664	70	665	71
rect	664	71	665	72
rect	664	72	665	73
rect	664	73	665	74
rect	664	74	665	75
rect	664	75	665	76
rect	664	76	665	77
rect	664	77	665	78
rect	664	78	665	79
rect	664	79	665	80
rect	664	80	665	81
rect	664	81	665	82
rect	664	82	665	83
rect	664	83	665	84
rect	664	84	665	85
rect	664	85	665	86
rect	664	86	665	87
rect	664	87	665	88
rect	664	88	665	89
rect	664	89	665	90
rect	664	90	665	91
rect	664	91	665	92
rect	664	92	665	93
rect	664	93	665	94
rect	664	94	665	95
rect	664	95	665	96
rect	664	96	665	97
rect	664	97	665	98
rect	664	98	665	99
rect	664	99	665	100
rect	664	100	665	101
rect	664	101	665	102
rect	664	102	665	103
rect	664	103	665	104
rect	664	104	665	105
rect	664	105	665	106
rect	664	106	665	107
rect	664	107	665	108
rect	664	108	665	109
rect	664	109	665	110
rect	664	110	665	111
rect	664	111	665	112
rect	664	112	665	113
rect	664	113	665	114
rect	664	114	665	115
rect	664	115	665	116
rect	664	116	665	117
rect	664	117	665	118
rect	664	118	665	119
rect	664	119	665	120
rect	664	120	665	121
rect	664	121	665	122
rect	664	122	665	123
rect	664	123	665	124
rect	664	124	665	125
rect	664	125	665	126
rect	664	126	665	127
rect	664	127	665	128
rect	664	128	665	129
rect	664	129	665	130
rect	664	130	665	131
rect	664	131	665	132
rect	664	132	665	133
rect	664	133	665	134
rect	664	134	665	135
rect	664	135	665	136
rect	664	136	665	137
rect	664	137	665	138
rect	664	138	665	139
rect	664	139	665	140
rect	664	140	665	141
rect	664	141	665	142
rect	664	142	665	143
rect	664	143	665	144
rect	664	144	665	145
rect	664	145	665	146
rect	664	146	665	147
rect	664	147	665	148
rect	664	148	665	149
rect	664	149	665	150
rect	664	150	665	151
rect	664	151	665	152
rect	664	152	665	153
rect	664	153	665	154
rect	664	154	665	155
rect	664	155	665	156
rect	664	156	665	157
rect	664	157	665	158
rect	664	158	665	159
rect	664	159	665	160
rect	664	160	665	161
rect	664	161	665	162
rect	664	162	665	163
rect	664	163	665	164
rect	664	164	665	165
rect	664	165	665	166
rect	664	166	665	167
rect	664	167	665	168
rect	665	0	666	1
rect	665	1	666	2
rect	665	2	666	3
rect	665	3	666	4
rect	665	4	666	5
rect	665	5	666	6
rect	665	6	666	7
rect	665	7	666	8
rect	665	8	666	9
rect	665	9	666	10
rect	665	10	666	11
rect	665	11	666	12
rect	665	12	666	13
rect	665	13	666	14
rect	665	14	666	15
rect	665	15	666	16
rect	665	16	666	17
rect	665	17	666	18
rect	665	18	666	19
rect	665	19	666	20
rect	665	20	666	21
rect	665	21	666	22
rect	665	22	666	23
rect	665	23	666	24
rect	665	24	666	25
rect	665	25	666	26
rect	665	26	666	27
rect	665	27	666	28
rect	665	28	666	29
rect	665	29	666	30
rect	665	30	666	31
rect	665	31	666	32
rect	665	32	666	33
rect	665	33	666	34
rect	665	34	666	35
rect	665	35	666	36
rect	665	36	666	37
rect	665	37	666	38
rect	665	38	666	39
rect	665	39	666	40
rect	665	40	666	41
rect	665	41	666	42
rect	665	42	666	43
rect	665	43	666	44
rect	665	44	666	45
rect	665	45	666	46
rect	665	46	666	47
rect	665	47	666	48
rect	665	48	666	49
rect	665	49	666	50
rect	665	50	666	51
rect	665	51	666	52
rect	665	52	666	53
rect	665	53	666	54
rect	665	54	666	55
rect	665	55	666	56
rect	665	56	666	57
rect	665	57	666	58
rect	665	58	666	59
rect	665	59	666	60
rect	665	60	666	61
rect	665	61	666	62
rect	665	62	666	63
rect	665	63	666	64
rect	665	64	666	65
rect	665	65	666	66
rect	665	66	666	67
rect	665	67	666	68
rect	665	68	666	69
rect	665	69	666	70
rect	665	70	666	71
rect	665	71	666	72
rect	665	72	666	73
rect	665	73	666	74
rect	665	74	666	75
rect	665	75	666	76
rect	665	76	666	77
rect	665	77	666	78
rect	665	78	666	79
rect	665	79	666	80
rect	665	80	666	81
rect	665	81	666	82
rect	665	82	666	83
rect	665	83	666	84
rect	665	84	666	85
rect	665	85	666	86
rect	665	86	666	87
rect	665	87	666	88
rect	665	88	666	89
rect	665	89	666	90
rect	665	90	666	91
rect	665	91	666	92
rect	665	92	666	93
rect	665	93	666	94
rect	665	94	666	95
rect	665	95	666	96
rect	665	96	666	97
rect	665	97	666	98
rect	665	98	666	99
rect	665	99	666	100
rect	665	100	666	101
rect	665	101	666	102
rect	665	102	666	103
rect	665	103	666	104
rect	665	104	666	105
rect	665	105	666	106
rect	665	106	666	107
rect	665	107	666	108
rect	665	108	666	109
rect	665	109	666	110
rect	665	110	666	111
rect	665	111	666	112
rect	665	112	666	113
rect	665	113	666	114
rect	665	114	666	115
rect	665	115	666	116
rect	665	116	666	117
rect	665	117	666	118
rect	665	118	666	119
rect	665	119	666	120
rect	665	120	666	121
rect	665	121	666	122
rect	665	122	666	123
rect	665	123	666	124
rect	665	124	666	125
rect	665	125	666	126
rect	665	126	666	127
rect	665	127	666	128
rect	665	128	666	129
rect	665	129	666	130
rect	665	130	666	131
rect	665	131	666	132
rect	665	132	666	133
rect	665	133	666	134
rect	665	134	666	135
rect	665	135	666	136
rect	665	136	666	137
rect	665	137	666	138
rect	665	138	666	139
rect	665	139	666	140
rect	665	140	666	141
rect	665	141	666	142
rect	665	142	666	143
rect	665	143	666	144
rect	665	144	666	145
rect	665	145	666	146
rect	665	146	666	147
rect	665	147	666	148
rect	665	148	666	149
rect	665	149	666	150
rect	665	150	666	151
rect	665	151	666	152
rect	665	152	666	153
rect	665	153	666	154
rect	665	154	666	155
rect	665	155	666	156
rect	665	156	666	157
rect	665	157	666	158
rect	665	158	666	159
rect	665	159	666	160
rect	665	160	666	161
rect	665	161	666	162
rect	665	162	666	163
rect	665	163	666	164
rect	665	164	666	165
rect	665	165	666	166
rect	665	166	666	167
rect	665	167	666	168
rect	666	0	667	1
rect	666	1	667	2
rect	666	2	667	3
rect	666	3	667	4
rect	666	4	667	5
rect	666	5	667	6
rect	666	6	667	7
rect	666	7	667	8
rect	666	8	667	9
rect	666	9	667	10
rect	666	10	667	11
rect	666	11	667	12
rect	666	12	667	13
rect	666	13	667	14
rect	666	14	667	15
rect	666	15	667	16
rect	666	16	667	17
rect	666	17	667	18
rect	666	18	667	19
rect	666	19	667	20
rect	666	20	667	21
rect	666	21	667	22
rect	666	22	667	23
rect	666	23	667	24
rect	666	24	667	25
rect	666	25	667	26
rect	666	26	667	27
rect	666	27	667	28
rect	666	28	667	29
rect	666	29	667	30
rect	666	30	667	31
rect	666	31	667	32
rect	666	32	667	33
rect	666	33	667	34
rect	666	34	667	35
rect	666	35	667	36
rect	666	36	667	37
rect	666	37	667	38
rect	666	38	667	39
rect	666	39	667	40
rect	666	40	667	41
rect	666	41	667	42
rect	666	42	667	43
rect	666	43	667	44
rect	666	44	667	45
rect	666	45	667	46
rect	666	46	667	47
rect	666	47	667	48
rect	666	48	667	49
rect	666	49	667	50
rect	666	50	667	51
rect	666	51	667	52
rect	666	52	667	53
rect	666	53	667	54
rect	666	54	667	55
rect	666	55	667	56
rect	666	56	667	57
rect	666	57	667	58
rect	666	58	667	59
rect	666	59	667	60
rect	666	60	667	61
rect	666	61	667	62
rect	666	62	667	63
rect	666	63	667	64
rect	666	64	667	65
rect	666	65	667	66
rect	666	66	667	67
rect	666	67	667	68
rect	666	68	667	69
rect	666	69	667	70
rect	666	70	667	71
rect	666	71	667	72
rect	666	72	667	73
rect	666	73	667	74
rect	666	74	667	75
rect	666	75	667	76
rect	666	76	667	77
rect	666	77	667	78
rect	666	78	667	79
rect	666	79	667	80
rect	666	80	667	81
rect	666	81	667	82
rect	666	82	667	83
rect	666	83	667	84
rect	666	84	667	85
rect	666	85	667	86
rect	666	86	667	87
rect	666	87	667	88
rect	666	88	667	89
rect	666	89	667	90
rect	666	90	667	91
rect	666	91	667	92
rect	666	92	667	93
rect	666	93	667	94
rect	666	94	667	95
rect	666	95	667	96
rect	666	96	667	97
rect	666	97	667	98
rect	666	98	667	99
rect	666	99	667	100
rect	666	100	667	101
rect	666	101	667	102
rect	666	102	667	103
rect	666	103	667	104
rect	666	104	667	105
rect	666	105	667	106
rect	666	106	667	107
rect	666	107	667	108
rect	666	108	667	109
rect	666	109	667	110
rect	666	110	667	111
rect	666	111	667	112
rect	666	112	667	113
rect	666	113	667	114
rect	666	114	667	115
rect	666	115	667	116
rect	666	116	667	117
rect	666	117	667	118
rect	666	118	667	119
rect	666	119	667	120
rect	666	120	667	121
rect	666	121	667	122
rect	666	122	667	123
rect	666	123	667	124
rect	666	124	667	125
rect	666	125	667	126
rect	666	126	667	127
rect	666	127	667	128
rect	666	128	667	129
rect	666	129	667	130
rect	666	130	667	131
rect	666	131	667	132
rect	666	132	667	133
rect	666	133	667	134
rect	666	134	667	135
rect	666	135	667	136
rect	666	136	667	137
rect	666	137	667	138
rect	666	138	667	139
rect	666	139	667	140
rect	666	140	667	141
rect	666	141	667	142
rect	666	142	667	143
rect	666	143	667	144
rect	666	144	667	145
rect	666	145	667	146
rect	666	146	667	147
rect	666	147	667	148
rect	666	148	667	149
rect	666	149	667	150
rect	666	150	667	151
rect	666	151	667	152
rect	666	152	667	153
rect	666	153	667	154
rect	666	154	667	155
rect	666	155	667	156
rect	666	156	667	157
rect	666	157	667	158
rect	666	158	667	159
rect	666	159	667	160
rect	666	160	667	161
rect	666	161	667	162
rect	666	162	667	163
rect	666	163	667	164
rect	666	164	667	165
rect	666	165	667	166
rect	666	166	667	167
rect	666	167	667	168
<< metal1 >>
rect	621	188	622	189
rect	621	189	622	190
rect	621	190	622	191
rect	621	191	622	192
rect	621	192	622	193
<< metal2 >>
rect	1	121	2	122
rect	1	172	2	173
rect	2	121	3	122
rect	2	172	3	173
rect	3	52	4	53
rect	3	58	4	59
rect	3	109	4	110
rect	3	115	4	116
rect	3	118	4	119
rect	3	121	4	122
rect	3	124	4	125
rect	3	136	4	137
rect	3	145	4	146
rect	3	172	4	173
rect	4	52	5	53
rect	4	58	5	59
rect	4	109	5	110
rect	4	115	5	116
rect	4	118	5	119
rect	4	121	5	122
rect	4	124	5	125
rect	4	136	5	137
rect	4	145	5	146
rect	4	172	5	173
rect	5	7	6	8
rect	5	52	6	53
rect	5	58	6	59
rect	5	79	6	80
rect	5	85	6	86
rect	5	91	6	92
rect	5	106	6	107
rect	5	109	6	110
rect	5	115	6	116
rect	5	118	6	119
rect	5	121	6	122
rect	5	124	6	125
rect	5	136	6	137
rect	5	142	6	143
rect	5	145	6	146
rect	5	172	6	173
rect	12	1	13	2
rect	12	4	13	5
rect	12	7	13	8
rect	12	13	13	14
rect	12	25	13	26
rect	12	28	13	29
rect	12	52	13	53
rect	12	67	13	68
rect	12	73	13	74
rect	12	79	13	80
rect	12	91	13	92
rect	12	94	13	95
rect	12	100	13	101
rect	12	106	13	107
rect	12	109	13	110
rect	12	118	13	119
rect	12	121	13	122
rect	12	124	13	125
rect	12	130	13	131
rect	12	145	13	146
rect	12	172	13	173
rect	13	1	14	2
rect	13	4	14	5
rect	13	7	14	8
rect	13	13	14	14
rect	13	25	14	26
rect	13	28	14	29
rect	13	52	14	53
rect	13	67	14	68
rect	13	73	14	74
rect	13	79	14	80
rect	13	91	14	92
rect	13	94	14	95
rect	13	100	14	101
rect	13	106	14	107
rect	13	109	14	110
rect	13	118	14	119
rect	13	121	14	122
rect	13	124	14	125
rect	13	145	14	146
rect	13	172	14	173
rect	14	1	15	2
rect	14	4	15	5
rect	14	7	15	8
rect	14	13	15	14
rect	14	25	15	26
rect	14	28	15	29
rect	14	52	15	53
rect	14	67	15	68
rect	14	73	15	74
rect	14	79	15	80
rect	14	91	15	92
rect	14	94	15	95
rect	14	100	15	101
rect	14	106	15	107
rect	14	109	15	110
rect	14	118	15	119
rect	14	121	15	122
rect	14	124	15	125
rect	14	145	15	146
rect	14	172	15	173
rect	14	202	15	203
rect	15	1	16	2
rect	15	4	16	5
rect	15	7	16	8
rect	15	13	16	14
rect	15	25	16	26
rect	15	28	16	29
rect	15	52	16	53
rect	15	67	16	68
rect	15	73	16	74
rect	15	79	16	80
rect	15	91	16	92
rect	15	94	16	95
rect	15	100	16	101
rect	15	106	16	107
rect	15	109	16	110
rect	15	118	16	119
rect	15	124	16	125
rect	15	145	16	146
rect	15	172	16	173
rect	15	202	16	203
rect	16	1	17	2
rect	16	4	17	5
rect	16	7	17	8
rect	16	13	17	14
rect	16	25	17	26
rect	16	28	17	29
rect	16	52	17	53
rect	16	67	17	68
rect	16	73	17	74
rect	16	79	17	80
rect	16	91	17	92
rect	16	94	17	95
rect	16	100	17	101
rect	16	106	17	107
rect	16	109	17	110
rect	16	118	17	119
rect	16	124	17	125
rect	16	145	17	146
rect	16	172	17	173
rect	16	202	17	203
rect	16	211	17	212
rect	17	1	18	2
rect	17	4	18	5
rect	17	7	18	8
rect	17	13	18	14
rect	17	25	18	26
rect	17	28	18	29
rect	17	52	18	53
rect	17	67	18	68
rect	17	73	18	74
rect	17	91	18	92
rect	17	94	18	95
rect	17	109	18	110
rect	17	124	18	125
rect	17	145	18	146
rect	17	202	18	203
rect	17	211	18	212
rect	18	1	19	2
rect	18	4	19	5
rect	18	7	19	8
rect	18	13	19	14
rect	18	25	19	26
rect	18	28	19	29
rect	18	52	19	53
rect	18	67	19	68
rect	18	73	19	74
rect	18	85	19	86
rect	18	91	19	92
rect	18	94	19	95
rect	18	109	19	110
rect	18	124	19	125
rect	18	130	19	131
rect	18	145	19	146
rect	18	178	19	179
rect	18	202	19	203
rect	18	211	19	212
rect	19	1	20	2
rect	19	4	20	5
rect	19	7	20	8
rect	19	13	20	14
rect	19	25	20	26
rect	19	28	20	29
rect	19	52	20	53
rect	19	67	20	68
rect	19	73	20	74
rect	19	85	20	86
rect	19	91	20	92
rect	19	94	20	95
rect	19	109	20	110
rect	19	124	20	125
rect	19	130	20	131
rect	19	145	20	146
rect	19	178	20	179
rect	19	202	20	203
rect	19	211	20	212
rect	20	1	21	2
rect	20	4	21	5
rect	20	7	21	8
rect	20	13	21	14
rect	20	25	21	26
rect	20	28	21	29
rect	20	52	21	53
rect	20	67	21	68
rect	20	73	21	74
rect	20	76	21	77
rect	20	85	21	86
rect	20	91	21	92
rect	20	94	21	95
rect	20	109	21	110
rect	20	124	21	125
rect	20	130	21	131
rect	20	145	21	146
rect	20	175	21	176
rect	20	178	21	179
rect	20	202	21	203
rect	20	211	21	212
rect	21	1	22	2
rect	21	4	22	5
rect	21	7	22	8
rect	21	13	22	14
rect	21	28	22	29
rect	21	52	22	53
rect	21	67	22	68
rect	21	73	22	74
rect	21	76	22	77
rect	21	85	22	86
rect	21	91	22	92
rect	21	94	22	95
rect	21	109	22	110
rect	21	124	22	125
rect	21	130	22	131
rect	21	145	22	146
rect	21	175	22	176
rect	21	178	22	179
rect	21	202	22	203
rect	21	211	22	212
rect	22	1	23	2
rect	22	4	23	5
rect	22	7	23	8
rect	22	13	23	14
rect	22	28	23	29
rect	22	52	23	53
rect	22	67	23	68
rect	22	73	23	74
rect	22	76	23	77
rect	22	85	23	86
rect	22	91	23	92
rect	22	94	23	95
rect	22	109	23	110
rect	22	124	23	125
rect	22	130	23	131
rect	22	145	23	146
rect	22	175	23	176
rect	22	178	23	179
rect	22	202	23	203
rect	22	211	23	212
rect	22	214	23	215
rect	23	1	24	2
rect	23	4	24	5
rect	23	7	24	8
rect	23	28	24	29
rect	23	52	24	53
rect	23	67	24	68
rect	23	73	24	74
rect	23	76	24	77
rect	23	85	24	86
rect	23	91	24	92
rect	23	94	24	95
rect	23	109	24	110
rect	23	124	24	125
rect	23	130	24	131
rect	23	145	24	146
rect	23	175	24	176
rect	23	178	24	179
rect	23	202	24	203
rect	23	211	24	212
rect	23	214	24	215
rect	24	1	25	2
rect	24	4	25	5
rect	24	7	25	8
rect	24	28	25	29
rect	24	52	25	53
rect	24	67	25	68
rect	24	73	25	74
rect	24	76	25	77
rect	24	85	25	86
rect	24	91	25	92
rect	24	94	25	95
rect	24	109	25	110
rect	24	124	25	125
rect	24	130	25	131
rect	24	145	25	146
rect	24	172	25	173
rect	24	175	25	176
rect	24	178	25	179
rect	24	202	25	203
rect	24	211	25	212
rect	24	214	25	215
rect	25	1	26	2
rect	25	7	26	8
rect	25	28	26	29
rect	25	67	26	68
rect	25	76	26	77
rect	25	85	26	86
rect	25	91	26	92
rect	25	130	26	131
rect	25	145	26	146
rect	25	172	26	173
rect	25	175	26	176
rect	25	178	26	179
rect	25	202	26	203
rect	25	211	26	212
rect	25	214	26	215
rect	26	1	27	2
rect	26	7	27	8
rect	26	28	27	29
rect	26	67	27	68
rect	26	76	27	77
rect	26	82	27	83
rect	26	85	27	86
rect	26	91	27	92
rect	26	106	27	107
rect	26	121	27	122
rect	26	130	27	131
rect	26	136	27	137
rect	26	145	27	146
rect	26	172	27	173
rect	26	175	27	176
rect	26	178	27	179
rect	26	202	27	203
rect	26	211	27	212
rect	26	214	27	215
rect	27	76	28	77
rect	27	82	28	83
rect	27	85	28	86
rect	27	106	28	107
rect	27	121	28	122
rect	27	130	28	131
rect	27	136	28	137
rect	27	172	28	173
rect	27	175	28	176
rect	27	178	28	179
rect	27	202	28	203
rect	27	211	28	212
rect	27	214	28	215
rect	28	10	29	11
rect	28	13	29	14
rect	28	16	29	17
rect	28	22	29	23
rect	28	25	29	26
rect	28	52	29	53
rect	28	55	29	56
rect	28	76	29	77
rect	28	79	29	80
rect	28	82	29	83
rect	28	85	29	86
rect	28	106	29	107
rect	28	109	29	110
rect	28	118	29	119
rect	28	121	29	122
rect	28	127	29	128
rect	28	130	29	131
rect	28	133	29	134
rect	28	136	29	137
rect	28	139	29	140
rect	28	163	29	164
rect	28	172	29	173
rect	28	175	29	176
rect	28	178	29	179
rect	28	187	29	188
rect	28	190	29	191
rect	28	202	29	203
rect	28	211	29	212
rect	28	214	29	215
rect	35	7	36	8
rect	35	13	36	14
rect	35	22	36	23
rect	35	25	36	26
rect	35	46	36	47
rect	35	52	36	53
rect	35	61	36	62
rect	35	79	36	80
rect	35	82	36	83
rect	35	85	36	86
rect	35	106	36	107
rect	35	109	36	110
rect	35	118	36	119
rect	35	121	36	122
rect	35	130	36	131
rect	35	133	36	134
rect	35	136	36	137
rect	35	145	36	146
rect	35	157	36	158
rect	35	163	36	164
rect	35	166	36	167
rect	35	172	36	173
rect	35	175	36	176
rect	35	178	36	179
rect	35	187	36	188
rect	35	202	36	203
rect	35	211	36	212
rect	35	214	36	215
rect	36	7	37	8
rect	36	13	37	14
rect	36	22	37	23
rect	36	25	37	26
rect	36	46	37	47
rect	36	52	37	53
rect	36	61	37	62
rect	36	79	37	80
rect	36	82	37	83
rect	36	85	37	86
rect	36	106	37	107
rect	36	109	37	110
rect	36	118	37	119
rect	36	121	37	122
rect	36	133	37	134
rect	36	136	37	137
rect	36	145	37	146
rect	36	157	37	158
rect	36	163	37	164
rect	36	166	37	167
rect	36	172	37	173
rect	36	175	37	176
rect	36	178	37	179
rect	36	187	37	188
rect	36	202	37	203
rect	36	211	37	212
rect	36	214	37	215
rect	37	7	38	8
rect	37	13	38	14
rect	37	22	38	23
rect	37	25	38	26
rect	37	46	38	47
rect	37	52	38	53
rect	37	61	38	62
rect	37	79	38	80
rect	37	82	38	83
rect	37	85	38	86
rect	37	106	38	107
rect	37	109	38	110
rect	37	118	38	119
rect	37	121	38	122
rect	37	133	38	134
rect	37	136	38	137
rect	37	142	38	143
rect	37	145	38	146
rect	37	157	38	158
rect	37	163	38	164
rect	37	166	38	167
rect	37	172	38	173
rect	37	175	38	176
rect	37	178	38	179
rect	37	187	38	188
rect	37	202	38	203
rect	37	211	38	212
rect	37	214	38	215
rect	38	7	39	8
rect	38	13	39	14
rect	38	22	39	23
rect	38	25	39	26
rect	38	46	39	47
rect	38	52	39	53
rect	38	61	39	62
rect	38	79	39	80
rect	38	82	39	83
rect	38	85	39	86
rect	38	106	39	107
rect	38	109	39	110
rect	38	118	39	119
rect	38	121	39	122
rect	38	133	39	134
rect	38	142	39	143
rect	38	145	39	146
rect	38	157	39	158
rect	38	163	39	164
rect	38	166	39	167
rect	38	172	39	173
rect	38	175	39	176
rect	38	178	39	179
rect	38	187	39	188
rect	38	202	39	203
rect	38	211	39	212
rect	38	214	39	215
rect	39	7	40	8
rect	39	13	40	14
rect	39	22	40	23
rect	39	25	40	26
rect	39	46	40	47
rect	39	52	40	53
rect	39	61	40	62
rect	39	79	40	80
rect	39	82	40	83
rect	39	85	40	86
rect	39	106	40	107
rect	39	109	40	110
rect	39	118	40	119
rect	39	121	40	122
rect	39	130	40	131
rect	39	133	40	134
rect	39	142	40	143
rect	39	145	40	146
rect	39	157	40	158
rect	39	163	40	164
rect	39	166	40	167
rect	39	172	40	173
rect	39	175	40	176
rect	39	178	40	179
rect	39	187	40	188
rect	39	202	40	203
rect	39	211	40	212
rect	39	214	40	215
rect	40	7	41	8
rect	40	13	41	14
rect	40	22	41	23
rect	40	25	41	26
rect	40	46	41	47
rect	40	52	41	53
rect	40	61	41	62
rect	40	79	41	80
rect	40	82	41	83
rect	40	85	41	86
rect	40	106	41	107
rect	40	109	41	110
rect	40	121	41	122
rect	40	130	41	131
rect	40	133	41	134
rect	40	142	41	143
rect	40	145	41	146
rect	40	163	41	164
rect	40	166	41	167
rect	40	172	41	173
rect	40	175	41	176
rect	40	178	41	179
rect	40	187	41	188
rect	40	202	41	203
rect	40	211	41	212
rect	40	214	41	215
rect	41	7	42	8
rect	41	13	42	14
rect	41	22	42	23
rect	41	25	42	26
rect	41	46	42	47
rect	41	52	42	53
rect	41	61	42	62
rect	41	79	42	80
rect	41	82	42	83
rect	41	85	42	86
rect	41	106	42	107
rect	41	109	42	110
rect	41	121	42	122
rect	41	130	42	131
rect	41	133	42	134
rect	41	142	42	143
rect	41	145	42	146
rect	41	154	42	155
rect	41	163	42	164
rect	41	166	42	167
rect	41	172	42	173
rect	41	175	42	176
rect	41	178	42	179
rect	41	187	42	188
rect	41	199	42	200
rect	41	202	42	203
rect	41	211	42	212
rect	41	214	42	215
rect	42	7	43	8
rect	42	13	43	14
rect	42	22	43	23
rect	42	25	43	26
rect	42	46	43	47
rect	42	52	43	53
rect	42	61	43	62
rect	42	79	43	80
rect	42	85	43	86
rect	42	106	43	107
rect	42	109	43	110
rect	42	121	43	122
rect	42	130	43	131
rect	42	133	43	134
rect	42	142	43	143
rect	42	145	43	146
rect	42	154	43	155
rect	42	163	43	164
rect	42	166	43	167
rect	42	172	43	173
rect	42	175	43	176
rect	42	178	43	179
rect	42	187	43	188
rect	42	199	43	200
rect	42	202	43	203
rect	42	211	43	212
rect	42	214	43	215
rect	43	7	44	8
rect	43	13	44	14
rect	43	22	44	23
rect	43	25	44	26
rect	43	46	44	47
rect	43	52	44	53
rect	43	61	44	62
rect	43	79	44	80
rect	43	85	44	86
rect	43	103	44	104
rect	43	106	44	107
rect	43	109	44	110
rect	43	112	44	113
rect	43	121	44	122
rect	43	130	44	131
rect	43	133	44	134
rect	43	142	44	143
rect	43	145	44	146
rect	43	154	44	155
rect	43	163	44	164
rect	43	166	44	167
rect	43	169	44	170
rect	43	172	44	173
rect	43	175	44	176
rect	43	178	44	179
rect	43	187	44	188
rect	43	199	44	200
rect	43	202	44	203
rect	43	211	44	212
rect	43	214	44	215
rect	44	7	45	8
rect	44	13	45	14
rect	44	22	45	23
rect	44	25	45	26
rect	44	46	45	47
rect	44	85	45	86
rect	44	103	45	104
rect	44	106	45	107
rect	44	112	45	113
rect	44	121	45	122
rect	44	130	45	131
rect	44	142	45	143
rect	44	154	45	155
rect	44	163	45	164
rect	44	166	45	167
rect	44	169	45	170
rect	44	172	45	173
rect	44	175	45	176
rect	44	178	45	179
rect	44	199	45	200
rect	44	202	45	203
rect	44	211	45	212
rect	44	214	45	215
rect	45	7	46	8
rect	45	13	46	14
rect	45	22	46	23
rect	45	25	46	26
rect	45	46	46	47
rect	45	55	46	56
rect	45	67	46	68
rect	45	85	46	86
rect	45	100	46	101
rect	45	103	46	104
rect	45	106	46	107
rect	45	112	46	113
rect	45	121	46	122
rect	45	124	46	125
rect	45	127	46	128
rect	45	130	46	131
rect	45	142	46	143
rect	45	154	46	155
rect	45	157	46	158
rect	45	163	46	164
rect	45	166	46	167
rect	45	169	46	170
rect	45	172	46	173
rect	45	175	46	176
rect	45	178	46	179
rect	45	199	46	200
rect	45	202	46	203
rect	45	208	46	209
rect	45	211	46	212
rect	45	214	46	215
rect	46	7	47	8
rect	46	25	47	26
rect	46	46	47	47
rect	46	55	47	56
rect	46	67	47	68
rect	46	85	47	86
rect	46	100	47	101
rect	46	103	47	104
rect	46	106	47	107
rect	46	112	47	113
rect	46	121	47	122
rect	46	124	47	125
rect	46	127	47	128
rect	46	130	47	131
rect	46	142	47	143
rect	46	154	47	155
rect	46	157	47	158
rect	46	163	47	164
rect	46	166	47	167
rect	46	169	47	170
rect	46	172	47	173
rect	46	175	47	176
rect	46	178	47	179
rect	46	199	47	200
rect	46	202	47	203
rect	46	208	47	209
rect	46	211	47	212
rect	46	214	47	215
rect	47	7	48	8
rect	47	16	48	17
rect	47	25	48	26
rect	47	31	48	32
rect	47	34	48	35
rect	47	46	48	47
rect	47	55	48	56
rect	47	67	48	68
rect	47	85	48	86
rect	47	100	48	101
rect	47	103	48	104
rect	47	106	48	107
rect	47	112	48	113
rect	47	121	48	122
rect	47	124	48	125
rect	47	127	48	128
rect	47	130	48	131
rect	47	142	48	143
rect	47	154	48	155
rect	47	157	48	158
rect	47	163	48	164
rect	47	166	48	167
rect	47	169	48	170
rect	47	172	48	173
rect	47	175	48	176
rect	47	178	48	179
rect	47	193	48	194
rect	47	199	48	200
rect	47	202	48	203
rect	47	208	48	209
rect	47	211	48	212
rect	47	214	48	215
rect	48	7	49	8
rect	48	16	49	17
rect	48	25	49	26
rect	48	31	49	32
rect	48	34	49	35
rect	48	46	49	47
rect	48	55	49	56
rect	48	67	49	68
rect	48	85	49	86
rect	48	100	49	101
rect	48	103	49	104
rect	48	106	49	107
rect	48	112	49	113
rect	48	121	49	122
rect	48	124	49	125
rect	48	127	49	128
rect	48	130	49	131
rect	48	142	49	143
rect	48	154	49	155
rect	48	157	49	158
rect	48	163	49	164
rect	48	166	49	167
rect	48	169	49	170
rect	48	172	49	173
rect	48	178	49	179
rect	48	193	49	194
rect	48	199	49	200
rect	48	202	49	203
rect	48	208	49	209
rect	48	214	49	215
rect	49	7	50	8
rect	49	10	50	11
rect	49	16	50	17
rect	49	25	50	26
rect	49	31	50	32
rect	49	34	50	35
rect	49	46	50	47
rect	49	55	50	56
rect	49	67	50	68
rect	49	85	50	86
rect	49	100	50	101
rect	49	103	50	104
rect	49	106	50	107
rect	49	112	50	113
rect	49	121	50	122
rect	49	124	50	125
rect	49	127	50	128
rect	49	130	50	131
rect	49	142	50	143
rect	49	145	50	146
rect	49	154	50	155
rect	49	157	50	158
rect	49	163	50	164
rect	49	166	50	167
rect	49	169	50	170
rect	49	172	50	173
rect	49	178	50	179
rect	49	190	50	191
rect	49	193	50	194
rect	49	199	50	200
rect	49	202	50	203
rect	49	208	50	209
rect	49	214	50	215
rect	49	238	50	239
rect	50	10	51	11
rect	50	16	51	17
rect	50	31	51	32
rect	50	34	51	35
rect	50	55	51	56
rect	50	67	51	68
rect	50	100	51	101
rect	50	103	51	104
rect	50	112	51	113
rect	50	121	51	122
rect	50	124	51	125
rect	50	127	51	128
rect	50	130	51	131
rect	50	142	51	143
rect	50	145	51	146
rect	50	154	51	155
rect	50	157	51	158
rect	50	169	51	170
rect	50	178	51	179
rect	50	190	51	191
rect	50	193	51	194
rect	50	199	51	200
rect	50	208	51	209
rect	50	238	51	239
rect	51	10	52	11
rect	51	13	52	14
rect	51	16	52	17
rect	51	19	52	20
rect	51	28	52	29
rect	51	31	52	32
rect	51	34	52	35
rect	51	40	52	41
rect	51	55	52	56
rect	51	64	52	65
rect	51	67	52	68
rect	51	76	52	77
rect	51	91	52	92
rect	51	97	52	98
rect	51	100	52	101
rect	51	103	52	104
rect	51	112	52	113
rect	51	121	52	122
rect	51	124	52	125
rect	51	127	52	128
rect	51	130	52	131
rect	51	139	52	140
rect	51	142	52	143
rect	51	145	52	146
rect	51	154	52	155
rect	51	157	52	158
rect	51	169	52	170
rect	51	178	52	179
rect	51	187	52	188
rect	51	190	52	191
rect	51	193	52	194
rect	51	199	52	200
rect	51	208	52	209
rect	51	211	52	212
rect	51	238	52	239
rect	51	241	52	242
rect	58	7	59	8
rect	58	13	59	14
rect	58	16	59	17
rect	58	19	59	20
rect	58	28	59	29
rect	58	31	59	32
rect	58	34	59	35
rect	58	40	59	41
rect	58	55	59	56
rect	58	61	59	62
rect	58	64	59	65
rect	58	67	59	68
rect	58	76	59	77
rect	58	79	59	80
rect	58	97	59	98
rect	58	100	59	101
rect	58	103	59	104
rect	58	112	59	113
rect	58	121	59	122
rect	58	124	59	125
rect	58	127	59	128
rect	58	130	59	131
rect	58	139	59	140
rect	58	142	59	143
rect	58	145	59	146
rect	58	154	59	155
rect	58	157	59	158
rect	58	163	59	164
rect	58	172	59	173
rect	58	175	59	176
rect	58	178	59	179
rect	58	187	59	188
rect	58	190	59	191
rect	58	199	59	200
rect	58	205	59	206
rect	58	208	59	209
rect	58	211	59	212
rect	58	220	59	221
rect	58	238	59	239
rect	58	241	59	242
rect	59	7	60	8
rect	59	13	60	14
rect	59	16	60	17
rect	59	19	60	20
rect	59	28	60	29
rect	59	31	60	32
rect	59	34	60	35
rect	59	40	60	41
rect	59	55	60	56
rect	59	61	60	62
rect	59	64	60	65
rect	59	67	60	68
rect	59	76	60	77
rect	59	79	60	80
rect	59	97	60	98
rect	59	100	60	101
rect	59	103	60	104
rect	59	112	60	113
rect	59	121	60	122
rect	59	124	60	125
rect	59	127	60	128
rect	59	130	60	131
rect	59	139	60	140
rect	59	142	60	143
rect	59	145	60	146
rect	59	154	60	155
rect	59	157	60	158
rect	59	163	60	164
rect	59	172	60	173
rect	59	175	60	176
rect	59	178	60	179
rect	59	187	60	188
rect	59	190	60	191
rect	59	205	60	206
rect	59	208	60	209
rect	59	211	60	212
rect	59	220	60	221
rect	59	238	60	239
rect	59	241	60	242
rect	60	7	61	8
rect	60	13	61	14
rect	60	16	61	17
rect	60	19	61	20
rect	60	28	61	29
rect	60	31	61	32
rect	60	34	61	35
rect	60	40	61	41
rect	60	55	61	56
rect	60	61	61	62
rect	60	64	61	65
rect	60	67	61	68
rect	60	76	61	77
rect	60	79	61	80
rect	60	97	61	98
rect	60	100	61	101
rect	60	103	61	104
rect	60	112	61	113
rect	60	121	61	122
rect	60	124	61	125
rect	60	127	61	128
rect	60	130	61	131
rect	60	139	61	140
rect	60	142	61	143
rect	60	145	61	146
rect	60	154	61	155
rect	60	157	61	158
rect	60	163	61	164
rect	60	172	61	173
rect	60	175	61	176
rect	60	178	61	179
rect	60	187	61	188
rect	60	190	61	191
rect	60	205	61	206
rect	60	208	61	209
rect	60	211	61	212
rect	60	220	61	221
rect	60	232	61	233
rect	60	238	61	239
rect	60	241	61	242
rect	61	7	62	8
rect	61	13	62	14
rect	61	16	62	17
rect	61	19	62	20
rect	61	28	62	29
rect	61	31	62	32
rect	61	34	62	35
rect	61	40	62	41
rect	61	55	62	56
rect	61	61	62	62
rect	61	64	62	65
rect	61	67	62	68
rect	61	76	62	77
rect	61	79	62	80
rect	61	97	62	98
rect	61	100	62	101
rect	61	103	62	104
rect	61	112	62	113
rect	61	124	62	125
rect	61	127	62	128
rect	61	130	62	131
rect	61	139	62	140
rect	61	142	62	143
rect	61	145	62	146
rect	61	154	62	155
rect	61	157	62	158
rect	61	163	62	164
rect	61	172	62	173
rect	61	175	62	176
rect	61	178	62	179
rect	61	187	62	188
rect	61	205	62	206
rect	61	208	62	209
rect	61	211	62	212
rect	61	220	62	221
rect	61	232	62	233
rect	61	238	62	239
rect	61	241	62	242
rect	62	7	63	8
rect	62	13	63	14
rect	62	16	63	17
rect	62	19	63	20
rect	62	28	63	29
rect	62	31	63	32
rect	62	34	63	35
rect	62	40	63	41
rect	62	55	63	56
rect	62	61	63	62
rect	62	64	63	65
rect	62	67	63	68
rect	62	76	63	77
rect	62	79	63	80
rect	62	97	63	98
rect	62	100	63	101
rect	62	103	63	104
rect	62	106	63	107
rect	62	112	63	113
rect	62	124	63	125
rect	62	127	63	128
rect	62	130	63	131
rect	62	139	63	140
rect	62	142	63	143
rect	62	145	63	146
rect	62	154	63	155
rect	62	157	63	158
rect	62	163	63	164
rect	62	172	63	173
rect	62	175	63	176
rect	62	178	63	179
rect	62	187	63	188
rect	62	199	63	200
rect	62	205	63	206
rect	62	208	63	209
rect	62	211	63	212
rect	62	220	63	221
rect	62	232	63	233
rect	62	238	63	239
rect	62	241	63	242
rect	63	7	64	8
rect	63	13	64	14
rect	63	16	64	17
rect	63	19	64	20
rect	63	28	64	29
rect	63	31	64	32
rect	63	34	64	35
rect	63	40	64	41
rect	63	55	64	56
rect	63	61	64	62
rect	63	64	64	65
rect	63	67	64	68
rect	63	76	64	77
rect	63	79	64	80
rect	63	97	64	98
rect	63	100	64	101
rect	63	106	64	107
rect	63	112	64	113
rect	63	124	64	125
rect	63	127	64	128
rect	63	130	64	131
rect	63	139	64	140
rect	63	142	64	143
rect	63	145	64	146
rect	63	154	64	155
rect	63	157	64	158
rect	63	163	64	164
rect	63	172	64	173
rect	63	175	64	176
rect	63	178	64	179
rect	63	187	64	188
rect	63	199	64	200
rect	63	208	64	209
rect	63	211	64	212
rect	63	220	64	221
rect	63	232	64	233
rect	63	238	64	239
rect	63	241	64	242
rect	64	7	65	8
rect	64	13	65	14
rect	64	16	65	17
rect	64	19	65	20
rect	64	28	65	29
rect	64	31	65	32
rect	64	34	65	35
rect	64	40	65	41
rect	64	55	65	56
rect	64	61	65	62
rect	64	64	65	65
rect	64	67	65	68
rect	64	76	65	77
rect	64	79	65	80
rect	64	97	65	98
rect	64	100	65	101
rect	64	106	65	107
rect	64	112	65	113
rect	64	124	65	125
rect	64	127	65	128
rect	64	130	65	131
rect	64	139	65	140
rect	64	142	65	143
rect	64	145	65	146
rect	64	154	65	155
rect	64	157	65	158
rect	64	163	65	164
rect	64	172	65	173
rect	64	175	65	176
rect	64	178	65	179
rect	64	187	65	188
rect	64	199	65	200
rect	64	208	65	209
rect	64	211	65	212
rect	64	220	65	221
rect	64	232	65	233
rect	64	238	65	239
rect	64	241	65	242
rect	65	7	66	8
rect	65	13	66	14
rect	65	16	66	17
rect	65	19	66	20
rect	65	31	66	32
rect	65	34	66	35
rect	65	40	66	41
rect	65	55	66	56
rect	65	61	66	62
rect	65	64	66	65
rect	65	67	66	68
rect	65	76	66	77
rect	65	79	66	80
rect	65	97	66	98
rect	65	100	66	101
rect	65	106	66	107
rect	65	124	66	125
rect	65	127	66	128
rect	65	130	66	131
rect	65	139	66	140
rect	65	142	66	143
rect	65	145	66	146
rect	65	157	66	158
rect	65	163	66	164
rect	65	172	66	173
rect	65	178	66	179
rect	65	187	66	188
rect	65	199	66	200
rect	65	208	66	209
rect	65	220	66	221
rect	65	232	66	233
rect	65	238	66	239
rect	65	241	66	242
rect	66	5	67	6
rect	66	7	67	8
rect	66	13	67	14
rect	66	16	67	17
rect	66	19	67	20
rect	66	31	67	32
rect	66	34	67	35
rect	66	40	67	41
rect	66	55	67	56
rect	66	61	67	62
rect	66	64	67	65
rect	66	67	67	68
rect	66	76	67	77
rect	66	79	67	80
rect	66	97	67	98
rect	66	100	67	101
rect	66	103	67	104
rect	66	106	67	107
rect	66	124	67	125
rect	66	127	67	128
rect	66	130	67	131
rect	66	139	67	140
rect	66	142	67	143
rect	66	145	67	146
rect	66	157	67	158
rect	66	163	67	164
rect	66	166	67	167
rect	66	172	67	173
rect	66	178	67	179
rect	66	187	67	188
rect	66	196	67	197
rect	66	199	67	200
rect	66	208	67	209
rect	66	217	67	218
rect	66	220	67	221
rect	66	232	67	233
rect	66	238	67	239
rect	66	241	67	242
rect	67	5	68	6
rect	67	7	68	8
rect	67	13	68	14
rect	67	19	68	20
rect	67	31	68	32
rect	67	34	68	35
rect	67	55	68	56
rect	67	61	68	62
rect	67	64	68	65
rect	67	67	68	68
rect	67	76	68	77
rect	67	79	68	80
rect	67	97	68	98
rect	67	103	68	104
rect	67	106	68	107
rect	67	124	68	125
rect	67	130	68	131
rect	67	142	68	143
rect	67	145	68	146
rect	67	157	68	158
rect	67	163	68	164
rect	67	166	68	167
rect	67	172	68	173
rect	67	196	68	197
rect	67	199	68	200
rect	67	208	68	209
rect	67	217	68	218
rect	67	220	68	221
rect	67	232	68	233
rect	67	238	68	239
rect	67	241	68	242
rect	68	5	69	6
rect	68	7	69	8
rect	68	13	69	14
rect	68	19	69	20
rect	68	28	69	29
rect	68	31	69	32
rect	68	34	69	35
rect	68	49	69	50
rect	68	55	69	56
rect	68	61	69	62
rect	68	64	69	65
rect	68	67	69	68
rect	68	76	69	77
rect	68	79	69	80
rect	68	97	69	98
rect	68	103	69	104
rect	68	106	69	107
rect	68	118	69	119
rect	68	121	69	122
rect	68	124	69	125
rect	68	130	69	131
rect	68	142	69	143
rect	68	145	69	146
rect	68	154	69	155
rect	68	157	69	158
rect	68	163	69	164
rect	68	166	69	167
rect	68	172	69	173
rect	68	175	69	176
rect	68	196	69	197
rect	68	199	69	200
rect	68	208	69	209
rect	68	211	69	212
rect	68	217	69	218
rect	68	220	69	221
rect	68	232	69	233
rect	68	238	69	239
rect	68	241	69	242
rect	69	5	70	6
rect	69	7	70	8
rect	69	19	70	20
rect	69	28	70	29
rect	69	34	70	35
rect	69	49	70	50
rect	69	55	70	56
rect	69	61	70	62
rect	69	64	70	65
rect	69	76	70	77
rect	69	79	70	80
rect	69	97	70	98
rect	69	103	70	104
rect	69	106	70	107
rect	69	118	70	119
rect	69	121	70	122
rect	69	124	70	125
rect	69	145	70	146
rect	69	154	70	155
rect	69	157	70	158
rect	69	163	70	164
rect	69	166	70	167
rect	69	172	70	173
rect	69	175	70	176
rect	69	196	70	197
rect	69	199	70	200
rect	69	208	70	209
rect	69	211	70	212
rect	69	217	70	218
rect	69	220	70	221
rect	69	232	70	233
rect	69	238	70	239
rect	70	5	71	6
rect	70	7	71	8
rect	70	19	71	20
rect	70	25	71	26
rect	70	28	71	29
rect	70	34	71	35
rect	70	40	71	41
rect	70	49	71	50
rect	70	55	71	56
rect	70	61	71	62
rect	70	64	71	65
rect	70	73	71	74
rect	70	76	71	77
rect	70	79	71	80
rect	70	97	71	98
rect	70	100	71	101
rect	70	103	71	104
rect	70	106	71	107
rect	70	112	71	113
rect	70	118	71	119
rect	70	121	71	122
rect	70	124	71	125
rect	70	127	71	128
rect	70	139	71	140
rect	70	145	71	146
rect	70	154	71	155
rect	70	157	71	158
rect	70	163	71	164
rect	70	166	71	167
rect	70	172	71	173
rect	70	175	71	176
rect	70	178	71	179
rect	70	181	71	182
rect	70	184	71	185
rect	70	190	71	191
rect	70	196	71	197
rect	70	199	71	200
rect	70	208	71	209
rect	70	211	71	212
rect	70	217	71	218
rect	70	220	71	221
rect	70	232	71	233
rect	70	238	71	239
rect	70	289	71	290
rect	71	5	72	6
rect	71	25	72	26
rect	71	28	72	29
rect	71	34	72	35
rect	71	40	72	41
rect	71	49	72	50
rect	71	55	72	56
rect	71	61	72	62
rect	71	73	72	74
rect	71	76	72	77
rect	71	79	72	80
rect	71	100	72	101
rect	71	103	72	104
rect	71	106	72	107
rect	71	112	72	113
rect	71	118	72	119
rect	71	121	72	122
rect	71	124	72	125
rect	71	127	72	128
rect	71	139	72	140
rect	71	154	72	155
rect	71	157	72	158
rect	71	163	72	164
rect	71	166	72	167
rect	71	175	72	176
rect	71	178	72	179
rect	71	181	72	182
rect	71	184	72	185
rect	71	190	72	191
rect	71	196	72	197
rect	71	199	72	200
rect	71	211	72	212
rect	71	217	72	218
rect	71	220	72	221
rect	71	232	72	233
rect	71	289	72	290
rect	72	5	73	6
rect	72	16	73	17
rect	72	25	73	26
rect	72	28	73	29
rect	72	31	73	32
rect	72	34	73	35
rect	72	40	73	41
rect	72	49	73	50
rect	72	55	73	56
rect	72	61	73	62
rect	72	73	73	74
rect	72	76	73	77
rect	72	79	73	80
rect	72	82	73	83
rect	72	85	73	86
rect	72	91	73	92
rect	72	100	73	101
rect	72	103	73	104
rect	72	106	73	107
rect	72	112	73	113
rect	72	115	73	116
rect	72	118	73	119
rect	72	121	73	122
rect	72	124	73	125
rect	72	127	73	128
rect	72	130	73	131
rect	72	136	73	137
rect	72	139	73	140
rect	72	142	73	143
rect	72	154	73	155
rect	72	157	73	158
rect	72	163	73	164
rect	72	166	73	167
rect	72	175	73	176
rect	72	178	73	179
rect	72	181	73	182
rect	72	184	73	185
rect	72	190	73	191
rect	72	193	73	194
rect	72	196	73	197
rect	72	199	73	200
rect	72	211	73	212
rect	72	214	73	215
rect	72	217	73	218
rect	72	220	73	221
rect	72	223	73	224
rect	72	229	73	230
rect	72	232	73	233
rect	72	286	73	287
rect	72	289	73	290
rect	73	16	74	17
rect	73	25	74	26
rect	73	28	74	29
rect	73	31	74	32
rect	73	40	74	41
rect	73	49	74	50
rect	73	73	74	74
rect	73	82	74	83
rect	73	85	74	86
rect	73	91	74	92
rect	73	100	74	101
rect	73	103	74	104
rect	73	106	74	107
rect	73	112	74	113
rect	73	115	74	116
rect	73	118	74	119
rect	73	121	74	122
rect	73	124	74	125
rect	73	127	74	128
rect	73	130	74	131
rect	73	136	74	137
rect	73	139	74	140
rect	73	142	74	143
rect	73	154	74	155
rect	73	157	74	158
rect	73	166	74	167
rect	73	175	74	176
rect	73	178	74	179
rect	73	181	74	182
rect	73	184	74	185
rect	73	190	74	191
rect	73	193	74	194
rect	73	196	74	197
rect	73	199	74	200
rect	73	211	74	212
rect	73	214	74	215
rect	73	217	74	218
rect	73	220	74	221
rect	73	223	74	224
rect	73	229	74	230
rect	73	232	74	233
rect	73	286	74	287
rect	73	289	74	290
rect	74	7	75	8
rect	74	10	75	11
rect	74	16	75	17
rect	74	19	75	20
rect	74	22	75	23
rect	74	25	75	26
rect	74	28	75	29
rect	74	31	75	32
rect	74	40	75	41
rect	74	49	75	50
rect	74	58	75	59
rect	74	67	75	68
rect	74	70	75	71
rect	74	73	75	74
rect	74	82	75	83
rect	74	85	75	86
rect	74	91	75	92
rect	74	100	75	101
rect	74	103	75	104
rect	74	106	75	107
rect	74	112	75	113
rect	74	115	75	116
rect	74	118	75	119
rect	74	121	75	122
rect	74	124	75	125
rect	74	127	75	128
rect	74	130	75	131
rect	74	136	75	137
rect	74	139	75	140
rect	74	142	75	143
rect	74	145	75	146
rect	74	154	75	155
rect	74	157	75	158
rect	74	166	75	167
rect	74	175	75	176
rect	74	178	75	179
rect	74	181	75	182
rect	74	184	75	185
rect	74	187	75	188
rect	74	190	75	191
rect	74	193	75	194
rect	74	196	75	197
rect	74	199	75	200
rect	74	208	75	209
rect	74	211	75	212
rect	74	214	75	215
rect	74	217	75	218
rect	74	220	75	221
rect	74	223	75	224
rect	74	226	75	227
rect	74	229	75	230
rect	74	232	75	233
rect	74	238	75	239
rect	74	241	75	242
rect	74	286	75	287
rect	74	289	75	290
rect	81	7	82	8
rect	81	16	82	17
rect	81	19	82	20
rect	81	22	82	23
rect	81	25	82	26
rect	81	28	82	29
rect	81	31	82	32
rect	81	34	82	35
rect	81	40	82	41
rect	81	49	82	50
rect	81	58	82	59
rect	81	67	82	68
rect	81	70	82	71
rect	81	73	82	74
rect	81	79	82	80
rect	81	82	82	83
rect	81	91	82	92
rect	81	100	82	101
rect	81	103	82	104
rect	81	106	82	107
rect	81	115	82	116
rect	81	118	82	119
rect	81	121	82	122
rect	81	124	82	125
rect	81	127	82	128
rect	81	136	82	137
rect	81	139	82	140
rect	81	142	82	143
rect	81	145	82	146
rect	81	154	82	155
rect	81	157	82	158
rect	81	166	82	167
rect	81	175	82	176
rect	81	178	82	179
rect	81	187	82	188
rect	81	190	82	191
rect	81	193	82	194
rect	81	196	82	197
rect	81	199	82	200
rect	81	202	82	203
rect	81	205	82	206
rect	81	208	82	209
rect	81	211	82	212
rect	81	214	82	215
rect	81	217	82	218
rect	81	220	82	221
rect	81	229	82	230
rect	81	232	82	233
rect	81	241	82	242
rect	81	253	82	254
rect	81	268	82	269
rect	81	286	82	287
rect	81	289	82	290
rect	82	7	83	8
rect	82	16	83	17
rect	82	19	83	20
rect	82	22	83	23
rect	82	25	83	26
rect	82	28	83	29
rect	82	31	83	32
rect	82	34	83	35
rect	82	40	83	41
rect	82	49	83	50
rect	82	58	83	59
rect	82	67	83	68
rect	82	70	83	71
rect	82	73	83	74
rect	82	79	83	80
rect	82	82	83	83
rect	82	91	83	92
rect	82	100	83	101
rect	82	103	83	104
rect	82	106	83	107
rect	82	115	83	116
rect	82	121	83	122
rect	82	124	83	125
rect	82	127	83	128
rect	82	136	83	137
rect	82	139	83	140
rect	82	142	83	143
rect	82	145	83	146
rect	82	154	83	155
rect	82	157	83	158
rect	82	166	83	167
rect	82	175	83	176
rect	82	178	83	179
rect	82	187	83	188
rect	82	190	83	191
rect	82	193	83	194
rect	82	196	83	197
rect	82	199	83	200
rect	82	202	83	203
rect	82	205	83	206
rect	82	211	83	212
rect	82	214	83	215
rect	82	217	83	218
rect	82	220	83	221
rect	82	229	83	230
rect	82	232	83	233
rect	82	241	83	242
rect	82	253	83	254
rect	82	268	83	269
rect	82	286	83	287
rect	82	289	83	290
rect	83	7	84	8
rect	83	16	84	17
rect	83	19	84	20
rect	83	22	84	23
rect	83	25	84	26
rect	83	28	84	29
rect	83	31	84	32
rect	83	34	84	35
rect	83	40	84	41
rect	83	49	84	50
rect	83	58	84	59
rect	83	67	84	68
rect	83	70	84	71
rect	83	73	84	74
rect	83	79	84	80
rect	83	82	84	83
rect	83	91	84	92
rect	83	100	84	101
rect	83	103	84	104
rect	83	106	84	107
rect	83	115	84	116
rect	83	121	84	122
rect	83	124	84	125
rect	83	127	84	128
rect	83	130	84	131
rect	83	136	84	137
rect	83	139	84	140
rect	83	142	84	143
rect	83	145	84	146
rect	83	154	84	155
rect	83	157	84	158
rect	83	166	84	167
rect	83	175	84	176
rect	83	178	84	179
rect	83	187	84	188
rect	83	190	84	191
rect	83	193	84	194
rect	83	196	84	197
rect	83	199	84	200
rect	83	202	84	203
rect	83	205	84	206
rect	83	211	84	212
rect	83	214	84	215
rect	83	217	84	218
rect	83	220	84	221
rect	83	226	84	227
rect	83	229	84	230
rect	83	232	84	233
rect	83	241	84	242
rect	83	253	84	254
rect	83	268	84	269
rect	83	286	84	287
rect	83	289	84	290
rect	84	7	85	8
rect	84	16	85	17
rect	84	19	85	20
rect	84	22	85	23
rect	84	25	85	26
rect	84	28	85	29
rect	84	31	85	32
rect	84	34	85	35
rect	84	40	85	41
rect	84	49	85	50
rect	84	58	85	59
rect	84	67	85	68
rect	84	70	85	71
rect	84	73	85	74
rect	84	79	85	80
rect	84	82	85	83
rect	84	91	85	92
rect	84	100	85	101
rect	84	103	85	104
rect	84	106	85	107
rect	84	115	85	116
rect	84	121	85	122
rect	84	124	85	125
rect	84	130	85	131
rect	84	136	85	137
rect	84	139	85	140
rect	84	142	85	143
rect	84	145	85	146
rect	84	154	85	155
rect	84	157	85	158
rect	84	166	85	167
rect	84	175	85	176
rect	84	178	85	179
rect	84	187	85	188
rect	84	190	85	191
rect	84	193	85	194
rect	84	196	85	197
rect	84	199	85	200
rect	84	202	85	203
rect	84	205	85	206
rect	84	211	85	212
rect	84	217	85	218
rect	84	220	85	221
rect	84	226	85	227
rect	84	229	85	230
rect	84	232	85	233
rect	84	241	85	242
rect	84	253	85	254
rect	84	268	85	269
rect	84	286	85	287
rect	84	289	85	290
rect	85	7	86	8
rect	85	16	86	17
rect	85	19	86	20
rect	85	22	86	23
rect	85	25	86	26
rect	85	28	86	29
rect	85	31	86	32
rect	85	34	86	35
rect	85	40	86	41
rect	85	49	86	50
rect	85	58	86	59
rect	85	67	86	68
rect	85	70	86	71
rect	85	73	86	74
rect	85	79	86	80
rect	85	82	86	83
rect	85	91	86	92
rect	85	100	86	101
rect	85	103	86	104
rect	85	106	86	107
rect	85	115	86	116
rect	85	118	86	119
rect	85	121	86	122
rect	85	124	86	125
rect	85	130	86	131
rect	85	136	86	137
rect	85	139	86	140
rect	85	142	86	143
rect	85	145	86	146
rect	85	154	86	155
rect	85	157	86	158
rect	85	166	86	167
rect	85	175	86	176
rect	85	178	86	179
rect	85	187	86	188
rect	85	190	86	191
rect	85	193	86	194
rect	85	196	86	197
rect	85	199	86	200
rect	85	202	86	203
rect	85	205	86	206
rect	85	208	86	209
rect	85	211	86	212
rect	85	217	86	218
rect	85	220	86	221
rect	85	226	86	227
rect	85	229	86	230
rect	85	232	86	233
rect	85	241	86	242
rect	85	253	86	254
rect	85	268	86	269
rect	85	286	86	287
rect	85	289	86	290
rect	86	7	87	8
rect	86	16	87	17
rect	86	19	87	20
rect	86	22	87	23
rect	86	25	87	26
rect	86	28	87	29
rect	86	31	87	32
rect	86	34	87	35
rect	86	40	87	41
rect	86	49	87	50
rect	86	58	87	59
rect	86	67	87	68
rect	86	70	87	71
rect	86	73	87	74
rect	86	79	87	80
rect	86	82	87	83
rect	86	91	87	92
rect	86	100	87	101
rect	86	103	87	104
rect	86	106	87	107
rect	86	118	87	119
rect	86	121	87	122
rect	86	124	87	125
rect	86	130	87	131
rect	86	136	87	137
rect	86	139	87	140
rect	86	142	87	143
rect	86	145	87	146
rect	86	154	87	155
rect	86	157	87	158
rect	86	166	87	167
rect	86	175	87	176
rect	86	178	87	179
rect	86	187	87	188
rect	86	190	87	191
rect	86	193	87	194
rect	86	199	87	200
rect	86	202	87	203
rect	86	205	87	206
rect	86	208	87	209
rect	86	211	87	212
rect	86	220	87	221
rect	86	226	87	227
rect	86	229	87	230
rect	86	232	87	233
rect	86	241	87	242
rect	86	253	87	254
rect	86	268	87	269
rect	86	286	87	287
rect	86	289	87	290
rect	87	7	88	8
rect	87	16	88	17
rect	87	19	88	20
rect	87	22	88	23
rect	87	25	88	26
rect	87	28	88	29
rect	87	31	88	32
rect	87	34	88	35
rect	87	40	88	41
rect	87	49	88	50
rect	87	58	88	59
rect	87	67	88	68
rect	87	70	88	71
rect	87	73	88	74
rect	87	79	88	80
rect	87	82	88	83
rect	87	91	88	92
rect	87	100	88	101
rect	87	103	88	104
rect	87	106	88	107
rect	87	118	88	119
rect	87	121	88	122
rect	87	124	88	125
rect	87	127	88	128
rect	87	130	88	131
rect	87	136	88	137
rect	87	139	88	140
rect	87	142	88	143
rect	87	145	88	146
rect	87	154	88	155
rect	87	157	88	158
rect	87	166	88	167
rect	87	175	88	176
rect	87	178	88	179
rect	87	187	88	188
rect	87	190	88	191
rect	87	193	88	194
rect	87	199	88	200
rect	87	202	88	203
rect	87	205	88	206
rect	87	208	88	209
rect	87	211	88	212
rect	87	214	88	215
rect	87	220	88	221
rect	87	226	88	227
rect	87	229	88	230
rect	87	232	88	233
rect	87	235	88	236
rect	87	241	88	242
rect	87	253	88	254
rect	87	268	88	269
rect	87	286	88	287
rect	87	289	88	290
rect	88	7	89	8
rect	88	16	89	17
rect	88	19	89	20
rect	88	22	89	23
rect	88	25	89	26
rect	88	28	89	29
rect	88	31	89	32
rect	88	34	89	35
rect	88	49	89	50
rect	88	58	89	59
rect	88	67	89	68
rect	88	70	89	71
rect	88	79	89	80
rect	88	82	89	83
rect	88	91	89	92
rect	88	100	89	101
rect	88	103	89	104
rect	88	118	89	119
rect	88	121	89	122
rect	88	124	89	125
rect	88	127	89	128
rect	88	130	89	131
rect	88	136	89	137
rect	88	139	89	140
rect	88	142	89	143
rect	88	145	89	146
rect	88	154	89	155
rect	88	157	89	158
rect	88	166	89	167
rect	88	175	89	176
rect	88	178	89	179
rect	88	187	89	188
rect	88	190	89	191
rect	88	193	89	194
rect	88	199	89	200
rect	88	202	89	203
rect	88	208	89	209
rect	88	214	89	215
rect	88	220	89	221
rect	88	226	89	227
rect	88	229	89	230
rect	88	232	89	233
rect	88	235	89	236
rect	88	241	89	242
rect	88	253	89	254
rect	88	268	89	269
rect	88	286	89	287
rect	88	289	89	290
rect	89	7	90	8
rect	89	16	90	17
rect	89	19	90	20
rect	89	22	90	23
rect	89	25	90	26
rect	89	28	90	29
rect	89	31	90	32
rect	89	34	90	35
rect	89	46	90	47
rect	89	49	90	50
rect	89	58	90	59
rect	89	67	90	68
rect	89	70	90	71
rect	89	76	90	77
rect	89	79	90	80
rect	89	82	90	83
rect	89	91	90	92
rect	89	100	90	101
rect	89	103	90	104
rect	89	115	90	116
rect	89	118	90	119
rect	89	121	90	122
rect	89	124	90	125
rect	89	127	90	128
rect	89	130	90	131
rect	89	136	90	137
rect	89	139	90	140
rect	89	142	90	143
rect	89	145	90	146
rect	89	154	90	155
rect	89	157	90	158
rect	89	166	90	167
rect	89	175	90	176
rect	89	178	90	179
rect	89	187	90	188
rect	89	190	90	191
rect	89	193	90	194
rect	89	196	90	197
rect	89	199	90	200
rect	89	202	90	203
rect	89	208	90	209
rect	89	214	90	215
rect	89	220	90	221
rect	89	226	90	227
rect	89	229	90	230
rect	89	232	90	233
rect	89	235	90	236
rect	89	241	90	242
rect	89	250	90	251
rect	89	253	90	254
rect	89	268	90	269
rect	89	286	90	287
rect	89	289	90	290
rect	90	7	91	8
rect	90	16	91	17
rect	90	19	91	20
rect	90	22	91	23
rect	90	28	91	29
rect	90	31	91	32
rect	90	34	91	35
rect	90	46	91	47
rect	90	58	91	59
rect	90	70	91	71
rect	90	76	91	77
rect	90	79	91	80
rect	90	82	91	83
rect	90	100	91	101
rect	90	103	91	104
rect	90	115	91	116
rect	90	118	91	119
rect	90	121	91	122
rect	90	124	91	125
rect	90	127	91	128
rect	90	130	91	131
rect	90	136	91	137
rect	90	139	91	140
rect	90	142	91	143
rect	90	154	91	155
rect	90	157	91	158
rect	90	166	91	167
rect	90	175	91	176
rect	90	178	91	179
rect	90	187	91	188
rect	90	190	91	191
rect	90	193	91	194
rect	90	196	91	197
rect	90	199	91	200
rect	90	208	91	209
rect	90	214	91	215
rect	90	226	91	227
rect	90	229	91	230
rect	90	232	91	233
rect	90	235	91	236
rect	90	241	91	242
rect	90	250	91	251
rect	90	253	91	254
rect	90	286	91	287
rect	90	289	91	290
rect	91	7	92	8
rect	91	16	92	17
rect	91	19	92	20
rect	91	22	92	23
rect	91	28	92	29
rect	91	31	92	32
rect	91	34	92	35
rect	91	43	92	44
rect	91	46	92	47
rect	91	58	92	59
rect	91	61	92	62
rect	91	70	92	71
rect	91	76	92	77
rect	91	79	92	80
rect	91	82	92	83
rect	91	85	92	86
rect	91	100	92	101
rect	91	103	92	104
rect	91	109	92	110
rect	91	115	92	116
rect	91	118	92	119
rect	91	121	92	122
rect	91	124	92	125
rect	91	127	92	128
rect	91	130	92	131
rect	91	136	92	137
rect	91	139	92	140
rect	91	142	92	143
rect	91	148	92	149
rect	91	154	92	155
rect	91	157	92	158
rect	91	166	92	167
rect	91	175	92	176
rect	91	178	92	179
rect	91	187	92	188
rect	91	190	92	191
rect	91	193	92	194
rect	91	196	92	197
rect	91	199	92	200
rect	91	205	92	206
rect	91	208	92	209
rect	91	211	92	212
rect	91	214	92	215
rect	91	226	92	227
rect	91	229	92	230
rect	91	232	92	233
rect	91	235	92	236
rect	91	241	92	242
rect	91	250	92	251
rect	91	253	92	254
rect	91	277	92	278
rect	91	286	92	287
rect	91	289	92	290
rect	92	7	93	8
rect	92	16	93	17
rect	92	22	93	23
rect	92	31	93	32
rect	92	34	93	35
rect	92	43	93	44
rect	92	46	93	47
rect	92	58	93	59
rect	92	61	93	62
rect	92	70	93	71
rect	92	76	93	77
rect	92	79	93	80
rect	92	82	93	83
rect	92	85	93	86
rect	92	100	93	101
rect	92	103	93	104
rect	92	109	93	110
rect	92	115	93	116
rect	92	118	93	119
rect	92	121	93	122
rect	92	124	93	125
rect	92	127	93	128
rect	92	130	93	131
rect	92	136	93	137
rect	92	139	93	140
rect	92	142	93	143
rect	92	148	93	149
rect	92	154	93	155
rect	92	157	93	158
rect	92	166	93	167
rect	92	175	93	176
rect	92	178	93	179
rect	92	187	93	188
rect	92	190	93	191
rect	92	193	93	194
rect	92	196	93	197
rect	92	205	93	206
rect	92	208	93	209
rect	92	211	93	212
rect	92	214	93	215
rect	92	226	93	227
rect	92	229	93	230
rect	92	235	93	236
rect	92	241	93	242
rect	92	250	93	251
rect	92	277	93	278
rect	92	286	93	287
rect	92	289	93	290
rect	93	7	94	8
rect	93	16	94	17
rect	93	22	94	23
rect	93	25	94	26
rect	93	31	94	32
rect	93	34	94	35
rect	93	43	94	44
rect	93	46	94	47
rect	93	49	94	50
rect	93	58	94	59
rect	93	61	94	62
rect	93	67	94	68
rect	93	70	94	71
rect	93	76	94	77
rect	93	79	94	80
rect	93	82	94	83
rect	93	85	94	86
rect	93	100	94	101
rect	93	103	94	104
rect	93	109	94	110
rect	93	115	94	116
rect	93	118	94	119
rect	93	121	94	122
rect	93	124	94	125
rect	93	127	94	128
rect	93	130	94	131
rect	93	136	94	137
rect	93	139	94	140
rect	93	142	94	143
rect	93	148	94	149
rect	93	154	94	155
rect	93	157	94	158
rect	93	166	94	167
rect	93	175	94	176
rect	93	178	94	179
rect	93	181	94	182
rect	93	187	94	188
rect	93	190	94	191
rect	93	193	94	194
rect	93	196	94	197
rect	93	205	94	206
rect	93	208	94	209
rect	93	211	94	212
rect	93	214	94	215
rect	93	217	94	218
rect	93	226	94	227
rect	93	229	94	230
rect	93	235	94	236
rect	93	238	94	239
rect	93	241	94	242
rect	93	250	94	251
rect	93	268	94	269
rect	93	277	94	278
rect	93	286	94	287
rect	93	289	94	290
rect	94	7	95	8
rect	94	16	95	17
rect	94	25	95	26
rect	94	43	95	44
rect	94	46	95	47
rect	94	49	95	50
rect	94	61	95	62
rect	94	67	95	68
rect	94	70	95	71
rect	94	76	95	77
rect	94	79	95	80
rect	94	85	95	86
rect	94	100	95	101
rect	94	109	95	110
rect	94	115	95	116
rect	94	118	95	119
rect	94	121	95	122
rect	94	124	95	125
rect	94	127	95	128
rect	94	130	95	131
rect	94	136	95	137
rect	94	139	95	140
rect	94	148	95	149
rect	94	154	95	155
rect	94	166	95	167
rect	94	175	95	176
rect	94	178	95	179
rect	94	181	95	182
rect	94	190	95	191
rect	94	193	95	194
rect	94	196	95	197
rect	94	205	95	206
rect	94	208	95	209
rect	94	211	95	212
rect	94	214	95	215
rect	94	217	95	218
rect	94	226	95	227
rect	94	235	95	236
rect	94	238	95	239
rect	94	241	95	242
rect	94	250	95	251
rect	94	268	95	269
rect	94	277	95	278
rect	94	286	95	287
rect	94	289	95	290
rect	95	7	96	8
rect	95	10	96	11
rect	95	16	96	17
rect	95	25	96	26
rect	95	28	96	29
rect	95	40	96	41
rect	95	43	96	44
rect	95	46	96	47
rect	95	49	96	50
rect	95	61	96	62
rect	95	67	96	68
rect	95	70	96	71
rect	95	73	96	74
rect	95	76	96	77
rect	95	79	96	80
rect	95	85	96	86
rect	95	94	96	95
rect	95	100	96	101
rect	95	106	96	107
rect	95	109	96	110
rect	95	115	96	116
rect	95	118	96	119
rect	95	121	96	122
rect	95	124	96	125
rect	95	127	96	128
rect	95	130	96	131
rect	95	136	96	137
rect	95	139	96	140
rect	95	145	96	146
rect	95	148	96	149
rect	95	154	96	155
rect	95	163	96	164
rect	95	166	96	167
rect	95	175	96	176
rect	95	178	96	179
rect	95	181	96	182
rect	95	190	96	191
rect	95	193	96	194
rect	95	196	96	197
rect	95	205	96	206
rect	95	208	96	209
rect	95	211	96	212
rect	95	214	96	215
rect	95	217	96	218
rect	95	220	96	221
rect	95	226	96	227
rect	95	235	96	236
rect	95	238	96	239
rect	95	241	96	242
rect	95	250	96	251
rect	95	253	96	254
rect	95	268	96	269
rect	95	277	96	278
rect	95	286	96	287
rect	95	289	96	290
rect	95	292	96	293
rect	95	298	96	299
rect	96	10	97	11
rect	96	25	97	26
rect	96	28	97	29
rect	96	40	97	41
rect	96	43	97	44
rect	96	46	97	47
rect	96	49	97	50
rect	96	61	97	62
rect	96	67	97	68
rect	96	73	97	74
rect	96	76	97	77
rect	96	85	97	86
rect	96	94	97	95
rect	96	100	97	101
rect	96	106	97	107
rect	96	109	97	110
rect	96	115	97	116
rect	96	118	97	119
rect	96	121	97	122
rect	96	124	97	125
rect	96	127	97	128
rect	96	130	97	131
rect	96	136	97	137
rect	96	145	97	146
rect	96	148	97	149
rect	96	163	97	164
rect	96	166	97	167
rect	96	175	97	176
rect	96	181	97	182
rect	96	190	97	191
rect	96	196	97	197
rect	96	205	97	206
rect	96	208	97	209
rect	96	211	97	212
rect	96	214	97	215
rect	96	217	97	218
rect	96	220	97	221
rect	96	226	97	227
rect	96	235	97	236
rect	96	238	97	239
rect	96	241	97	242
rect	96	250	97	251
rect	96	253	97	254
rect	96	268	97	269
rect	96	277	97	278
rect	96	286	97	287
rect	96	292	97	293
rect	96	298	97	299
rect	97	10	98	11
rect	97	13	98	14
rect	97	22	98	23
rect	97	25	98	26
rect	97	28	98	29
rect	97	31	98	32
rect	97	34	98	35
rect	97	40	98	41
rect	97	43	98	44
rect	97	46	98	47
rect	97	49	98	50
rect	97	55	98	56
rect	97	58	98	59
rect	97	61	98	62
rect	97	64	98	65
rect	97	67	98	68
rect	97	73	98	74
rect	97	76	98	77
rect	97	85	98	86
rect	97	94	98	95
rect	97	100	98	101
rect	97	103	98	104
rect	97	106	98	107
rect	97	109	98	110
rect	97	115	98	116
rect	97	118	98	119
rect	97	121	98	122
rect	97	124	98	125
rect	97	127	98	128
rect	97	130	98	131
rect	97	136	98	137
rect	97	142	98	143
rect	97	145	98	146
rect	97	148	98	149
rect	97	160	98	161
rect	97	163	98	164
rect	97	166	98	167
rect	97	175	98	176
rect	97	181	98	182
rect	97	187	98	188
rect	97	190	98	191
rect	97	196	98	197
rect	97	205	98	206
rect	97	208	98	209
rect	97	211	98	212
rect	97	214	98	215
rect	97	217	98	218
rect	97	220	98	221
rect	97	226	98	227
rect	97	232	98	233
rect	97	235	98	236
rect	97	238	98	239
rect	97	241	98	242
rect	97	250	98	251
rect	97	253	98	254
rect	97	268	98	269
rect	97	277	98	278
rect	97	286	98	287
rect	97	292	98	293
rect	97	298	98	299
rect	97	310	98	311
rect	98	10	99	11
rect	98	13	99	14
rect	98	22	99	23
rect	98	25	99	26
rect	98	28	99	29
rect	98	31	99	32
rect	98	34	99	35
rect	98	40	99	41
rect	98	43	99	44
rect	98	46	99	47
rect	98	49	99	50
rect	98	55	99	56
rect	98	58	99	59
rect	98	61	99	62
rect	98	64	99	65
rect	98	67	99	68
rect	98	73	99	74
rect	98	76	99	77
rect	98	85	99	86
rect	98	94	99	95
rect	98	103	99	104
rect	98	106	99	107
rect	98	109	99	110
rect	98	115	99	116
rect	98	118	99	119
rect	98	127	99	128
rect	98	130	99	131
rect	98	142	99	143
rect	98	145	99	146
rect	98	148	99	149
rect	98	160	99	161
rect	98	163	99	164
rect	98	181	99	182
rect	98	187	99	188
rect	98	196	99	197
rect	98	205	99	206
rect	98	208	99	209
rect	98	211	99	212
rect	98	214	99	215
rect	98	217	99	218
rect	98	220	99	221
rect	98	226	99	227
rect	98	232	99	233
rect	98	235	99	236
rect	98	238	99	239
rect	98	241	99	242
rect	98	250	99	251
rect	98	253	99	254
rect	98	268	99	269
rect	98	277	99	278
rect	98	292	99	293
rect	98	298	99	299
rect	98	310	99	311
rect	99	7	100	8
rect	99	10	100	11
rect	99	13	100	14
rect	99	22	100	23
rect	99	25	100	26
rect	99	28	100	29
rect	99	31	100	32
rect	99	34	100	35
rect	99	40	100	41
rect	99	43	100	44
rect	99	46	100	47
rect	99	49	100	50
rect	99	55	100	56
rect	99	58	100	59
rect	99	61	100	62
rect	99	64	100	65
rect	99	67	100	68
rect	99	73	100	74
rect	99	76	100	77
rect	99	85	100	86
rect	99	94	100	95
rect	99	103	100	104
rect	99	106	100	107
rect	99	109	100	110
rect	99	112	100	113
rect	99	115	100	116
rect	99	118	100	119
rect	99	127	100	128
rect	99	130	100	131
rect	99	133	100	134
rect	99	142	100	143
rect	99	145	100	146
rect	99	148	100	149
rect	99	157	100	158
rect	99	160	100	161
rect	99	163	100	164
rect	99	172	100	173
rect	99	181	100	182
rect	99	184	100	185
rect	99	187	100	188
rect	99	196	100	197
rect	99	205	100	206
rect	99	208	100	209
rect	99	211	100	212
rect	99	214	100	215
rect	99	217	100	218
rect	99	220	100	221
rect	99	226	100	227
rect	99	229	100	230
rect	99	232	100	233
rect	99	235	100	236
rect	99	238	100	239
rect	99	241	100	242
rect	99	250	100	251
rect	99	253	100	254
rect	99	268	100	269
rect	99	277	100	278
rect	99	292	100	293
rect	99	298	100	299
rect	99	307	100	308
rect	99	310	100	311
rect	106	13	107	14
rect	106	22	107	23
rect	106	25	107	26
rect	106	28	107	29
rect	106	31	107	32
rect	106	37	107	38
rect	106	40	107	41
rect	106	43	107	44
rect	106	46	107	47
rect	106	49	107	50
rect	106	58	107	59
rect	106	61	107	62
rect	106	64	107	65
rect	106	70	107	71
rect	106	73	107	74
rect	106	76	107	77
rect	106	85	107	86
rect	106	94	107	95
rect	106	103	107	104
rect	106	106	107	107
rect	106	109	107	110
rect	106	112	107	113
rect	106	115	107	116
rect	106	118	107	119
rect	106	124	107	125
rect	106	127	107	128
rect	106	130	107	131
rect	106	133	107	134
rect	106	136	107	137
rect	106	142	107	143
rect	106	145	107	146
rect	106	148	107	149
rect	106	154	107	155
rect	106	157	107	158
rect	106	160	107	161
rect	106	163	107	164
rect	106	166	107	167
rect	106	169	107	170
rect	106	172	107	173
rect	106	175	107	176
rect	106	181	107	182
rect	106	184	107	185
rect	106	187	107	188
rect	106	196	107	197
rect	106	205	107	206
rect	106	208	107	209
rect	106	211	107	212
rect	106	214	107	215
rect	106	217	107	218
rect	106	226	107	227
rect	106	229	107	230
rect	106	232	107	233
rect	106	235	107	236
rect	106	238	107	239
rect	106	241	107	242
rect	106	250	107	251
rect	106	253	107	254
rect	106	265	107	266
rect	106	268	107	269
rect	106	271	107	272
rect	106	277	107	278
rect	106	289	107	290
rect	106	292	107	293
rect	106	307	107	308
rect	106	310	107	311
rect	107	13	108	14
rect	107	22	108	23
rect	107	25	108	26
rect	107	28	108	29
rect	107	31	108	32
rect	107	37	108	38
rect	107	40	108	41
rect	107	43	108	44
rect	107	46	108	47
rect	107	49	108	50
rect	107	58	108	59
rect	107	61	108	62
rect	107	64	108	65
rect	107	70	108	71
rect	107	73	108	74
rect	107	76	108	77
rect	107	85	108	86
rect	107	94	108	95
rect	107	103	108	104
rect	107	106	108	107
rect	107	109	108	110
rect	107	112	108	113
rect	107	115	108	116
rect	107	118	108	119
rect	107	124	108	125
rect	107	127	108	128
rect	107	130	108	131
rect	107	133	108	134
rect	107	136	108	137
rect	107	142	108	143
rect	107	145	108	146
rect	107	154	108	155
rect	107	157	108	158
rect	107	160	108	161
rect	107	163	108	164
rect	107	166	108	167
rect	107	169	108	170
rect	107	172	108	173
rect	107	175	108	176
rect	107	181	108	182
rect	107	184	108	185
rect	107	187	108	188
rect	107	196	108	197
rect	107	205	108	206
rect	107	208	108	209
rect	107	211	108	212
rect	107	214	108	215
rect	107	217	108	218
rect	107	226	108	227
rect	107	229	108	230
rect	107	232	108	233
rect	107	235	108	236
rect	107	238	108	239
rect	107	241	108	242
rect	107	250	108	251
rect	107	253	108	254
rect	107	265	108	266
rect	107	268	108	269
rect	107	271	108	272
rect	107	277	108	278
rect	107	289	108	290
rect	107	292	108	293
rect	107	307	108	308
rect	107	310	108	311
rect	108	13	109	14
rect	108	22	109	23
rect	108	25	109	26
rect	108	28	109	29
rect	108	31	109	32
rect	108	37	109	38
rect	108	40	109	41
rect	108	43	109	44
rect	108	46	109	47
rect	108	49	109	50
rect	108	58	109	59
rect	108	61	109	62
rect	108	64	109	65
rect	108	70	109	71
rect	108	73	109	74
rect	108	76	109	77
rect	108	85	109	86
rect	108	94	109	95
rect	108	101	109	102
rect	108	103	109	104
rect	108	106	109	107
rect	108	109	109	110
rect	108	112	109	113
rect	108	115	109	116
rect	108	118	109	119
rect	108	124	109	125
rect	108	127	109	128
rect	108	130	109	131
rect	108	133	109	134
rect	108	136	109	137
rect	108	142	109	143
rect	108	145	109	146
rect	108	154	109	155
rect	108	157	109	158
rect	108	160	109	161
rect	108	163	109	164
rect	108	166	109	167
rect	108	169	109	170
rect	108	172	109	173
rect	108	175	109	176
rect	108	181	109	182
rect	108	184	109	185
rect	108	187	109	188
rect	108	196	109	197
rect	108	205	109	206
rect	108	208	109	209
rect	108	211	109	212
rect	108	214	109	215
rect	108	217	109	218
rect	108	226	109	227
rect	108	229	109	230
rect	108	232	109	233
rect	108	235	109	236
rect	108	238	109	239
rect	108	241	109	242
rect	108	250	109	251
rect	108	253	109	254
rect	108	265	109	266
rect	108	268	109	269
rect	108	271	109	272
rect	108	277	109	278
rect	108	289	109	290
rect	108	292	109	293
rect	108	307	109	308
rect	108	310	109	311
rect	109	13	110	14
rect	109	22	110	23
rect	109	25	110	26
rect	109	28	110	29
rect	109	31	110	32
rect	109	37	110	38
rect	109	40	110	41
rect	109	43	110	44
rect	109	46	110	47
rect	109	49	110	50
rect	109	58	110	59
rect	109	61	110	62
rect	109	64	110	65
rect	109	70	110	71
rect	109	73	110	74
rect	109	76	110	77
rect	109	85	110	86
rect	109	94	110	95
rect	109	101	110	102
rect	109	103	110	104
rect	109	106	110	107
rect	109	109	110	110
rect	109	112	110	113
rect	109	115	110	116
rect	109	118	110	119
rect	109	124	110	125
rect	109	127	110	128
rect	109	130	110	131
rect	109	133	110	134
rect	109	136	110	137
rect	109	142	110	143
rect	109	145	110	146
rect	109	157	110	158
rect	109	160	110	161
rect	109	163	110	164
rect	109	166	110	167
rect	109	169	110	170
rect	109	172	110	173
rect	109	175	110	176
rect	109	181	110	182
rect	109	184	110	185
rect	109	187	110	188
rect	109	196	110	197
rect	109	205	110	206
rect	109	208	110	209
rect	109	211	110	212
rect	109	214	110	215
rect	109	217	110	218
rect	109	226	110	227
rect	109	229	110	230
rect	109	232	110	233
rect	109	235	110	236
rect	109	238	110	239
rect	109	241	110	242
rect	109	250	110	251
rect	109	253	110	254
rect	109	265	110	266
rect	109	268	110	269
rect	109	271	110	272
rect	109	277	110	278
rect	109	289	110	290
rect	109	292	110	293
rect	109	307	110	308
rect	109	310	110	311
rect	110	13	111	14
rect	110	22	111	23
rect	110	25	111	26
rect	110	28	111	29
rect	110	31	111	32
rect	110	37	111	38
rect	110	40	111	41
rect	110	43	111	44
rect	110	46	111	47
rect	110	49	111	50
rect	110	58	111	59
rect	110	61	111	62
rect	110	64	111	65
rect	110	70	111	71
rect	110	73	111	74
rect	110	76	111	77
rect	110	85	111	86
rect	110	94	111	95
rect	110	101	111	102
rect	110	103	111	104
rect	110	106	111	107
rect	110	109	111	110
rect	110	112	111	113
rect	110	115	111	116
rect	110	118	111	119
rect	110	124	111	125
rect	110	127	111	128
rect	110	130	111	131
rect	110	133	111	134
rect	110	136	111	137
rect	110	142	111	143
rect	110	145	111	146
rect	110	148	111	149
rect	110	157	111	158
rect	110	160	111	161
rect	110	163	111	164
rect	110	166	111	167
rect	110	169	111	170
rect	110	172	111	173
rect	110	175	111	176
rect	110	181	111	182
rect	110	184	111	185
rect	110	187	111	188
rect	110	196	111	197
rect	110	205	111	206
rect	110	208	111	209
rect	110	211	111	212
rect	110	214	111	215
rect	110	217	111	218
rect	110	226	111	227
rect	110	229	111	230
rect	110	232	111	233
rect	110	235	111	236
rect	110	238	111	239
rect	110	241	111	242
rect	110	250	111	251
rect	110	253	111	254
rect	110	265	111	266
rect	110	268	111	269
rect	110	271	111	272
rect	110	277	111	278
rect	110	289	111	290
rect	110	292	111	293
rect	110	307	111	308
rect	110	310	111	311
rect	111	13	112	14
rect	111	22	112	23
rect	111	25	112	26
rect	111	28	112	29
rect	111	31	112	32
rect	111	37	112	38
rect	111	40	112	41
rect	111	43	112	44
rect	111	46	112	47
rect	111	49	112	50
rect	111	58	112	59
rect	111	61	112	62
rect	111	64	112	65
rect	111	70	112	71
rect	111	73	112	74
rect	111	76	112	77
rect	111	85	112	86
rect	111	94	112	95
rect	111	103	112	104
rect	111	106	112	107
rect	111	109	112	110
rect	111	112	112	113
rect	111	115	112	116
rect	111	118	112	119
rect	111	124	112	125
rect	111	127	112	128
rect	111	130	112	131
rect	111	133	112	134
rect	111	136	112	137
rect	111	142	112	143
rect	111	145	112	146
rect	111	148	112	149
rect	111	157	112	158
rect	111	160	112	161
rect	111	163	112	164
rect	111	166	112	167
rect	111	169	112	170
rect	111	172	112	173
rect	111	175	112	176
rect	111	181	112	182
rect	111	184	112	185
rect	111	187	112	188
rect	111	196	112	197
rect	111	205	112	206
rect	111	208	112	209
rect	111	211	112	212
rect	111	214	112	215
rect	111	217	112	218
rect	111	226	112	227
rect	111	229	112	230
rect	111	232	112	233
rect	111	235	112	236
rect	111	238	112	239
rect	111	241	112	242
rect	111	250	112	251
rect	111	253	112	254
rect	111	265	112	266
rect	111	268	112	269
rect	111	271	112	272
rect	111	277	112	278
rect	111	289	112	290
rect	111	292	112	293
rect	111	307	112	308
rect	111	310	112	311
rect	112	13	113	14
rect	112	22	113	23
rect	112	25	113	26
rect	112	28	113	29
rect	112	31	113	32
rect	112	37	113	38
rect	112	40	113	41
rect	112	43	113	44
rect	112	46	113	47
rect	112	49	113	50
rect	112	58	113	59
rect	112	61	113	62
rect	112	64	113	65
rect	112	70	113	71
rect	112	73	113	74
rect	112	76	113	77
rect	112	85	113	86
rect	112	94	113	95
rect	112	103	113	104
rect	112	106	113	107
rect	112	109	113	110
rect	112	112	113	113
rect	112	115	113	116
rect	112	118	113	119
rect	112	124	113	125
rect	112	127	113	128
rect	112	130	113	131
rect	112	133	113	134
rect	112	136	113	137
rect	112	142	113	143
rect	112	145	113	146
rect	112	148	113	149
rect	112	154	113	155
rect	112	157	113	158
rect	112	160	113	161
rect	112	163	113	164
rect	112	166	113	167
rect	112	169	113	170
rect	112	172	113	173
rect	112	175	113	176
rect	112	181	113	182
rect	112	184	113	185
rect	112	187	113	188
rect	112	196	113	197
rect	112	205	113	206
rect	112	208	113	209
rect	112	211	113	212
rect	112	214	113	215
rect	112	217	113	218
rect	112	226	113	227
rect	112	229	113	230
rect	112	232	113	233
rect	112	235	113	236
rect	112	238	113	239
rect	112	241	113	242
rect	112	250	113	251
rect	112	253	113	254
rect	112	265	113	266
rect	112	268	113	269
rect	112	271	113	272
rect	112	277	113	278
rect	112	289	113	290
rect	112	292	113	293
rect	112	307	113	308
rect	112	310	113	311
rect	113	13	114	14
rect	113	22	114	23
rect	113	25	114	26
rect	113	28	114	29
rect	113	31	114	32
rect	113	37	114	38
rect	113	40	114	41
rect	113	43	114	44
rect	113	46	114	47
rect	113	49	114	50
rect	113	58	114	59
rect	113	61	114	62
rect	113	64	114	65
rect	113	70	114	71
rect	113	73	114	74
rect	113	76	114	77
rect	113	85	114	86
rect	113	94	114	95
rect	113	106	114	107
rect	113	109	114	110
rect	113	112	114	113
rect	113	115	114	116
rect	113	118	114	119
rect	113	124	114	125
rect	113	127	114	128
rect	113	130	114	131
rect	113	133	114	134
rect	113	136	114	137
rect	113	142	114	143
rect	113	145	114	146
rect	113	148	114	149
rect	113	154	114	155
rect	113	157	114	158
rect	113	160	114	161
rect	113	163	114	164
rect	113	166	114	167
rect	113	169	114	170
rect	113	172	114	173
rect	113	175	114	176
rect	113	181	114	182
rect	113	184	114	185
rect	113	187	114	188
rect	113	196	114	197
rect	113	205	114	206
rect	113	208	114	209
rect	113	211	114	212
rect	113	214	114	215
rect	113	217	114	218
rect	113	226	114	227
rect	113	229	114	230
rect	113	232	114	233
rect	113	235	114	236
rect	113	238	114	239
rect	113	241	114	242
rect	113	253	114	254
rect	113	265	114	266
rect	113	268	114	269
rect	113	271	114	272
rect	113	277	114	278
rect	113	289	114	290
rect	113	292	114	293
rect	113	307	114	308
rect	113	310	114	311
rect	114	13	115	14
rect	114	22	115	23
rect	114	25	115	26
rect	114	28	115	29
rect	114	31	115	32
rect	114	37	115	38
rect	114	40	115	41
rect	114	43	115	44
rect	114	46	115	47
rect	114	49	115	50
rect	114	58	115	59
rect	114	61	115	62
rect	114	64	115	65
rect	114	70	115	71
rect	114	73	115	74
rect	114	76	115	77
rect	114	85	115	86
rect	114	94	115	95
rect	114	106	115	107
rect	114	109	115	110
rect	114	112	115	113
rect	114	115	115	116
rect	114	118	115	119
rect	114	121	115	122
rect	114	124	115	125
rect	114	127	115	128
rect	114	130	115	131
rect	114	133	115	134
rect	114	136	115	137
rect	114	142	115	143
rect	114	145	115	146
rect	114	148	115	149
rect	114	154	115	155
rect	114	157	115	158
rect	114	160	115	161
rect	114	163	115	164
rect	114	166	115	167
rect	114	169	115	170
rect	114	172	115	173
rect	114	175	115	176
rect	114	181	115	182
rect	114	184	115	185
rect	114	187	115	188
rect	114	196	115	197
rect	114	205	115	206
rect	114	208	115	209
rect	114	211	115	212
rect	114	214	115	215
rect	114	217	115	218
rect	114	226	115	227
rect	114	229	115	230
rect	114	232	115	233
rect	114	235	115	236
rect	114	238	115	239
rect	114	241	115	242
rect	114	244	115	245
rect	114	253	115	254
rect	114	265	115	266
rect	114	268	115	269
rect	114	271	115	272
rect	114	277	115	278
rect	114	289	115	290
rect	114	292	115	293
rect	114	307	115	308
rect	114	310	115	311
rect	115	13	116	14
rect	115	22	116	23
rect	115	25	116	26
rect	115	28	116	29
rect	115	31	116	32
rect	115	37	116	38
rect	115	40	116	41
rect	115	43	116	44
rect	115	46	116	47
rect	115	49	116	50
rect	115	58	116	59
rect	115	61	116	62
rect	115	64	116	65
rect	115	70	116	71
rect	115	73	116	74
rect	115	76	116	77
rect	115	85	116	86
rect	115	94	116	95
rect	115	106	116	107
rect	115	109	116	110
rect	115	118	116	119
rect	115	121	116	122
rect	115	127	116	128
rect	115	130	116	131
rect	115	133	116	134
rect	115	136	116	137
rect	115	142	116	143
rect	115	145	116	146
rect	115	148	116	149
rect	115	154	116	155
rect	115	157	116	158
rect	115	160	116	161
rect	115	163	116	164
rect	115	166	116	167
rect	115	169	116	170
rect	115	172	116	173
rect	115	175	116	176
rect	115	181	116	182
rect	115	184	116	185
rect	115	187	116	188
rect	115	196	116	197
rect	115	205	116	206
rect	115	208	116	209
rect	115	211	116	212
rect	115	214	116	215
rect	115	217	116	218
rect	115	226	116	227
rect	115	229	116	230
rect	115	232	116	233
rect	115	238	116	239
rect	115	241	116	242
rect	115	244	116	245
rect	115	253	116	254
rect	115	265	116	266
rect	115	268	116	269
rect	115	271	116	272
rect	115	277	116	278
rect	115	289	116	290
rect	115	292	116	293
rect	115	307	116	308
rect	115	310	116	311
rect	116	13	117	14
rect	116	22	117	23
rect	116	25	117	26
rect	116	28	117	29
rect	116	31	117	32
rect	116	37	117	38
rect	116	40	117	41
rect	116	43	117	44
rect	116	46	117	47
rect	116	49	117	50
rect	116	58	117	59
rect	116	61	117	62
rect	116	64	117	65
rect	116	70	117	71
rect	116	73	117	74
rect	116	76	117	77
rect	116	85	117	86
rect	116	94	117	95
rect	116	103	117	104
rect	116	106	117	107
rect	116	109	117	110
rect	116	118	117	119
rect	116	121	117	122
rect	116	127	117	128
rect	116	130	117	131
rect	116	133	117	134
rect	116	136	117	137
rect	116	142	117	143
rect	116	145	117	146
rect	116	148	117	149
rect	116	154	117	155
rect	116	157	117	158
rect	116	160	117	161
rect	116	163	117	164
rect	116	166	117	167
rect	116	169	117	170
rect	116	172	117	173
rect	116	175	117	176
rect	116	181	117	182
rect	116	184	117	185
rect	116	187	117	188
rect	116	196	117	197
rect	116	205	117	206
rect	116	208	117	209
rect	116	211	117	212
rect	116	214	117	215
rect	116	217	117	218
rect	116	226	117	227
rect	116	229	117	230
rect	116	232	117	233
rect	116	238	117	239
rect	116	241	117	242
rect	116	244	117	245
rect	116	250	117	251
rect	116	253	117	254
rect	116	265	117	266
rect	116	268	117	269
rect	116	271	117	272
rect	116	277	117	278
rect	116	289	117	290
rect	116	292	117	293
rect	116	307	117	308
rect	116	310	117	311
rect	117	13	118	14
rect	117	22	118	23
rect	117	25	118	26
rect	117	28	118	29
rect	117	31	118	32
rect	117	37	118	38
rect	117	40	118	41
rect	117	43	118	44
rect	117	46	118	47
rect	117	49	118	50
rect	117	58	118	59
rect	117	61	118	62
rect	117	64	118	65
rect	117	70	118	71
rect	117	73	118	74
rect	117	76	118	77
rect	117	85	118	86
rect	117	94	118	95
rect	117	103	118	104
rect	117	106	118	107
rect	117	109	118	110
rect	117	118	118	119
rect	117	121	118	122
rect	117	127	118	128
rect	117	130	118	131
rect	117	133	118	134
rect	117	136	118	137
rect	117	142	118	143
rect	117	145	118	146
rect	117	148	118	149
rect	117	154	118	155
rect	117	157	118	158
rect	117	160	118	161
rect	117	163	118	164
rect	117	166	118	167
rect	117	169	118	170
rect	117	172	118	173
rect	117	181	118	182
rect	117	184	118	185
rect	117	187	118	188
rect	117	196	118	197
rect	117	205	118	206
rect	117	208	118	209
rect	117	211	118	212
rect	117	214	118	215
rect	117	226	118	227
rect	117	229	118	230
rect	117	232	118	233
rect	117	238	118	239
rect	117	241	118	242
rect	117	244	118	245
rect	117	250	118	251
rect	117	253	118	254
rect	117	265	118	266
rect	117	268	118	269
rect	117	271	118	272
rect	117	289	118	290
rect	117	292	118	293
rect	117	307	118	308
rect	117	310	118	311
rect	118	13	119	14
rect	118	22	119	23
rect	118	25	119	26
rect	118	28	119	29
rect	118	31	119	32
rect	118	37	119	38
rect	118	40	119	41
rect	118	43	119	44
rect	118	46	119	47
rect	118	49	119	50
rect	118	58	119	59
rect	118	61	119	62
rect	118	64	119	65
rect	118	70	119	71
rect	118	73	119	74
rect	118	76	119	77
rect	118	85	119	86
rect	118	94	119	95
rect	118	103	119	104
rect	118	106	119	107
rect	118	109	119	110
rect	118	112	119	113
rect	118	118	119	119
rect	118	121	119	122
rect	118	127	119	128
rect	118	130	119	131
rect	118	133	119	134
rect	118	136	119	137
rect	118	142	119	143
rect	118	145	119	146
rect	118	148	119	149
rect	118	154	119	155
rect	118	157	119	158
rect	118	160	119	161
rect	118	163	119	164
rect	118	166	119	167
rect	118	169	119	170
rect	118	172	119	173
rect	118	181	119	182
rect	118	184	119	185
rect	118	187	119	188
rect	118	196	119	197
rect	118	205	119	206
rect	118	208	119	209
rect	118	211	119	212
rect	118	214	119	215
rect	118	226	119	227
rect	118	229	119	230
rect	118	232	119	233
rect	118	235	119	236
rect	118	238	119	239
rect	118	241	119	242
rect	118	244	119	245
rect	118	250	119	251
rect	118	253	119	254
rect	118	265	119	266
rect	118	268	119	269
rect	118	271	119	272
rect	118	274	119	275
rect	118	289	119	290
rect	118	292	119	293
rect	118	307	119	308
rect	118	310	119	311
rect	119	13	120	14
rect	119	22	120	23
rect	119	25	120	26
rect	119	28	120	29
rect	119	31	120	32
rect	119	37	120	38
rect	119	40	120	41
rect	119	43	120	44
rect	119	46	120	47
rect	119	49	120	50
rect	119	61	120	62
rect	119	64	120	65
rect	119	70	120	71
rect	119	73	120	74
rect	119	76	120	77
rect	119	85	120	86
rect	119	94	120	95
rect	119	103	120	104
rect	119	106	120	107
rect	119	109	120	110
rect	119	112	120	113
rect	119	118	120	119
rect	119	121	120	122
rect	119	127	120	128
rect	119	130	120	131
rect	119	133	120	134
rect	119	136	120	137
rect	119	142	120	143
rect	119	145	120	146
rect	119	148	120	149
rect	119	154	120	155
rect	119	157	120	158
rect	119	160	120	161
rect	119	163	120	164
rect	119	169	120	170
rect	119	172	120	173
rect	119	181	120	182
rect	119	184	120	185
rect	119	187	120	188
rect	119	196	120	197
rect	119	208	120	209
rect	119	211	120	212
rect	119	214	120	215
rect	119	226	120	227
rect	119	229	120	230
rect	119	232	120	233
rect	119	235	120	236
rect	119	238	120	239
rect	119	241	120	242
rect	119	244	120	245
rect	119	250	120	251
rect	119	265	120	266
rect	119	268	120	269
rect	119	271	120	272
rect	119	274	120	275
rect	119	289	120	290
rect	119	292	120	293
rect	119	307	120	308
rect	119	310	120	311
rect	120	13	121	14
rect	120	22	121	23
rect	120	25	121	26
rect	120	28	121	29
rect	120	31	121	32
rect	120	37	121	38
rect	120	40	121	41
rect	120	43	121	44
rect	120	46	121	47
rect	120	49	121	50
rect	120	61	121	62
rect	120	64	121	65
rect	120	70	121	71
rect	120	73	121	74
rect	120	76	121	77
rect	120	85	121	86
rect	120	94	121	95
rect	120	103	121	104
rect	120	106	121	107
rect	120	109	121	110
rect	120	112	121	113
rect	120	118	121	119
rect	120	121	121	122
rect	120	127	121	128
rect	120	130	121	131
rect	120	133	121	134
rect	120	136	121	137
rect	120	142	121	143
rect	120	145	121	146
rect	120	148	121	149
rect	120	154	121	155
rect	120	157	121	158
rect	120	160	121	161
rect	120	163	121	164
rect	120	169	121	170
rect	120	172	121	173
rect	120	181	121	182
rect	120	184	121	185
rect	120	187	121	188
rect	120	196	121	197
rect	120	208	121	209
rect	120	211	121	212
rect	120	214	121	215
rect	120	217	121	218
rect	120	226	121	227
rect	120	229	121	230
rect	120	232	121	233
rect	120	235	121	236
rect	120	238	121	239
rect	120	241	121	242
rect	120	244	121	245
rect	120	250	121	251
rect	120	265	121	266
rect	120	268	121	269
rect	120	271	121	272
rect	120	274	121	275
rect	120	277	121	278
rect	120	289	121	290
rect	120	292	121	293
rect	120	307	121	308
rect	120	310	121	311
rect	121	13	122	14
rect	121	22	122	23
rect	121	25	122	26
rect	121	28	122	29
rect	121	31	122	32
rect	121	37	122	38
rect	121	40	122	41
rect	121	43	122	44
rect	121	46	122	47
rect	121	49	122	50
rect	121	61	122	62
rect	121	64	122	65
rect	121	70	122	71
rect	121	73	122	74
rect	121	76	122	77
rect	121	85	122	86
rect	121	94	122	95
rect	121	103	122	104
rect	121	106	122	107
rect	121	112	122	113
rect	121	118	122	119
rect	121	121	122	122
rect	121	127	122	128
rect	121	130	122	131
rect	121	133	122	134
rect	121	136	122	137
rect	121	142	122	143
rect	121	148	122	149
rect	121	154	122	155
rect	121	160	122	161
rect	121	163	122	164
rect	121	169	122	170
rect	121	172	122	173
rect	121	184	122	185
rect	121	187	122	188
rect	121	196	122	197
rect	121	208	122	209
rect	121	211	122	212
rect	121	214	122	215
rect	121	217	122	218
rect	121	226	122	227
rect	121	229	122	230
rect	121	232	122	233
rect	121	235	122	236
rect	121	238	122	239
rect	121	241	122	242
rect	121	244	122	245
rect	121	250	122	251
rect	121	265	122	266
rect	121	268	122	269
rect	121	274	122	275
rect	121	277	122	278
rect	121	289	122	290
rect	121	292	122	293
rect	121	307	122	308
rect	121	310	122	311
rect	122	13	123	14
rect	122	22	123	23
rect	122	25	123	26
rect	122	28	123	29
rect	122	31	123	32
rect	122	37	123	38
rect	122	40	123	41
rect	122	43	123	44
rect	122	46	123	47
rect	122	49	123	50
rect	122	61	123	62
rect	122	64	123	65
rect	122	70	123	71
rect	122	73	123	74
rect	122	76	123	77
rect	122	85	123	86
rect	122	94	123	95
rect	122	103	123	104
rect	122	106	123	107
rect	122	112	123	113
rect	122	115	123	116
rect	122	118	123	119
rect	122	121	123	122
rect	122	127	123	128
rect	122	130	123	131
rect	122	133	123	134
rect	122	136	123	137
rect	122	142	123	143
rect	122	148	123	149
rect	122	151	123	152
rect	122	154	123	155
rect	122	160	123	161
rect	122	163	123	164
rect	122	166	123	167
rect	122	169	123	170
rect	122	172	123	173
rect	122	184	123	185
rect	122	187	123	188
rect	122	196	123	197
rect	122	205	123	206
rect	122	208	123	209
rect	122	211	123	212
rect	122	214	123	215
rect	122	217	123	218
rect	122	226	123	227
rect	122	229	123	230
rect	122	232	123	233
rect	122	235	123	236
rect	122	238	123	239
rect	122	241	123	242
rect	122	244	123	245
rect	122	247	123	248
rect	122	250	123	251
rect	122	265	123	266
rect	122	268	123	269
rect	122	274	123	275
rect	122	277	123	278
rect	122	289	123	290
rect	122	292	123	293
rect	122	307	123	308
rect	122	310	123	311
rect	123	13	124	14
rect	123	22	124	23
rect	123	25	124	26
rect	123	28	124	29
rect	123	31	124	32
rect	123	37	124	38
rect	123	40	124	41
rect	123	43	124	44
rect	123	46	124	47
rect	123	49	124	50
rect	123	61	124	62
rect	123	64	124	65
rect	123	70	124	71
rect	123	73	124	74
rect	123	76	124	77
rect	123	94	124	95
rect	123	103	124	104
rect	123	106	124	107
rect	123	112	124	113
rect	123	115	124	116
rect	123	121	124	122
rect	123	127	124	128
rect	123	130	124	131
rect	123	133	124	134
rect	123	142	124	143
rect	123	148	124	149
rect	123	151	124	152
rect	123	154	124	155
rect	123	160	124	161
rect	123	163	124	164
rect	123	166	124	167
rect	123	169	124	170
rect	123	184	124	185
rect	123	187	124	188
rect	123	196	124	197
rect	123	205	124	206
rect	123	211	124	212
rect	123	214	124	215
rect	123	217	124	218
rect	123	226	124	227
rect	123	229	124	230
rect	123	235	124	236
rect	123	238	124	239
rect	123	241	124	242
rect	123	244	124	245
rect	123	247	124	248
rect	123	250	124	251
rect	123	265	124	266
rect	123	268	124	269
rect	123	274	124	275
rect	123	277	124	278
rect	123	289	124	290
rect	123	292	124	293
rect	123	307	124	308
rect	123	310	124	311
rect	124	13	125	14
rect	124	22	125	23
rect	124	25	125	26
rect	124	28	125	29
rect	124	31	125	32
rect	124	37	125	38
rect	124	40	125	41
rect	124	43	125	44
rect	124	46	125	47
rect	124	49	125	50
rect	124	61	125	62
rect	124	64	125	65
rect	124	70	125	71
rect	124	73	125	74
rect	124	76	125	77
rect	124	91	125	92
rect	124	94	125	95
rect	124	103	125	104
rect	124	106	125	107
rect	124	109	125	110
rect	124	112	125	113
rect	124	115	125	116
rect	124	121	125	122
rect	124	127	125	128
rect	124	130	125	131
rect	124	133	125	134
rect	124	142	125	143
rect	124	148	125	149
rect	124	151	125	152
rect	124	154	125	155
rect	124	157	125	158
rect	124	160	125	161
rect	124	163	125	164
rect	124	166	125	167
rect	124	169	125	170
rect	124	181	125	182
rect	124	184	125	185
rect	124	187	125	188
rect	124	196	125	197
rect	124	205	125	206
rect	124	211	125	212
rect	124	214	125	215
rect	124	217	125	218
rect	124	223	125	224
rect	124	226	125	227
rect	124	229	125	230
rect	124	235	125	236
rect	124	238	125	239
rect	124	241	125	242
rect	124	244	125	245
rect	124	247	125	248
rect	124	250	125	251
rect	124	256	125	257
rect	124	265	125	266
rect	124	268	125	269
rect	124	274	125	275
rect	124	277	125	278
rect	124	289	125	290
rect	124	292	125	293
rect	124	307	125	308
rect	124	310	125	311
rect	125	13	126	14
rect	125	22	126	23
rect	125	25	126	26
rect	125	28	126	29
rect	125	31	126	32
rect	125	37	126	38
rect	125	40	126	41
rect	125	43	126	44
rect	125	46	126	47
rect	125	49	126	50
rect	125	61	126	62
rect	125	70	126	71
rect	125	76	126	77
rect	125	91	126	92
rect	125	94	126	95
rect	125	103	126	104
rect	125	109	126	110
rect	125	112	126	113
rect	125	115	126	116
rect	125	121	126	122
rect	125	127	126	128
rect	125	130	126	131
rect	125	142	126	143
rect	125	148	126	149
rect	125	151	126	152
rect	125	154	126	155
rect	125	157	126	158
rect	125	160	126	161
rect	125	163	126	164
rect	125	166	126	167
rect	125	181	126	182
rect	125	184	126	185
rect	125	187	126	188
rect	125	196	126	197
rect	125	205	126	206
rect	125	211	126	212
rect	125	217	126	218
rect	125	223	126	224
rect	125	226	126	227
rect	125	229	126	230
rect	125	235	126	236
rect	125	238	126	239
rect	125	244	126	245
rect	125	247	126	248
rect	125	250	126	251
rect	125	256	126	257
rect	125	265	126	266
rect	125	268	126	269
rect	125	274	126	275
rect	125	277	126	278
rect	125	289	126	290
rect	125	292	126	293
rect	125	307	126	308
rect	125	310	126	311
rect	126	13	127	14
rect	126	22	127	23
rect	126	25	127	26
rect	126	28	127	29
rect	126	31	127	32
rect	126	37	127	38
rect	126	40	127	41
rect	126	43	127	44
rect	126	46	127	47
rect	126	49	127	50
rect	126	55	127	56
rect	126	61	127	62
rect	126	70	127	71
rect	126	76	127	77
rect	126	85	127	86
rect	126	91	127	92
rect	126	94	127	95
rect	126	103	127	104
rect	126	109	127	110
rect	126	112	127	113
rect	126	115	127	116
rect	126	118	127	119
rect	126	121	127	122
rect	126	127	127	128
rect	126	130	127	131
rect	126	142	127	143
rect	126	145	127	146
rect	126	148	127	149
rect	126	151	127	152
rect	126	154	127	155
rect	126	157	127	158
rect	126	160	127	161
rect	126	163	127	164
rect	126	166	127	167
rect	126	181	127	182
rect	126	184	127	185
rect	126	187	127	188
rect	126	196	127	197
rect	126	205	127	206
rect	126	208	127	209
rect	126	211	127	212
rect	126	217	127	218
rect	126	223	127	224
rect	126	226	127	227
rect	126	229	127	230
rect	126	232	127	233
rect	126	235	127	236
rect	126	238	127	239
rect	126	244	127	245
rect	126	247	127	248
rect	126	250	127	251
rect	126	256	127	257
rect	126	262	127	263
rect	126	265	127	266
rect	126	268	127	269
rect	126	274	127	275
rect	126	277	127	278
rect	126	289	127	290
rect	126	292	127	293
rect	126	307	127	308
rect	126	310	127	311
rect	127	13	128	14
rect	127	22	128	23
rect	127	25	128	26
rect	127	28	128	29
rect	127	31	128	32
rect	127	37	128	38
rect	127	40	128	41
rect	127	43	128	44
rect	127	46	128	47
rect	127	55	128	56
rect	127	61	128	62
rect	127	76	128	77
rect	127	85	128	86
rect	127	91	128	92
rect	127	94	128	95
rect	127	103	128	104
rect	127	109	128	110
rect	127	112	128	113
rect	127	115	128	116
rect	127	118	128	119
rect	127	121	128	122
rect	127	127	128	128
rect	127	130	128	131
rect	127	142	128	143
rect	127	145	128	146
rect	127	148	128	149
rect	127	151	128	152
rect	127	154	128	155
rect	127	157	128	158
rect	127	160	128	161
rect	127	163	128	164
rect	127	166	128	167
rect	127	181	128	182
rect	127	184	128	185
rect	127	187	128	188
rect	127	196	128	197
rect	127	205	128	206
rect	127	208	128	209
rect	127	211	128	212
rect	127	217	128	218
rect	127	223	128	224
rect	127	226	128	227
rect	127	229	128	230
rect	127	232	128	233
rect	127	235	128	236
rect	127	238	128	239
rect	127	244	128	245
rect	127	247	128	248
rect	127	250	128	251
rect	127	256	128	257
rect	127	262	128	263
rect	127	265	128	266
rect	127	268	128	269
rect	127	274	128	275
rect	127	277	128	278
rect	127	289	128	290
rect	127	307	128	308
rect	127	310	128	311
rect	128	13	129	14
rect	128	22	129	23
rect	128	25	129	26
rect	128	28	129	29
rect	128	31	129	32
rect	128	37	129	38
rect	128	40	129	41
rect	128	43	129	44
rect	128	46	129	47
rect	128	55	129	56
rect	128	58	129	59
rect	128	61	129	62
rect	128	76	129	77
rect	128	85	129	86
rect	128	91	129	92
rect	128	94	129	95
rect	128	103	129	104
rect	128	109	129	110
rect	128	112	129	113
rect	128	115	129	116
rect	128	118	129	119
rect	128	121	129	122
rect	128	127	129	128
rect	128	130	129	131
rect	128	142	129	143
rect	128	145	129	146
rect	128	148	129	149
rect	128	151	129	152
rect	128	154	129	155
rect	128	157	129	158
rect	128	160	129	161
rect	128	163	129	164
rect	128	166	129	167
rect	128	181	129	182
rect	128	184	129	185
rect	128	187	129	188
rect	128	196	129	197
rect	128	205	129	206
rect	128	208	129	209
rect	128	211	129	212
rect	128	217	129	218
rect	128	223	129	224
rect	128	226	129	227
rect	128	229	129	230
rect	128	232	129	233
rect	128	235	129	236
rect	128	238	129	239
rect	128	244	129	245
rect	128	247	129	248
rect	128	250	129	251
rect	128	256	129	257
rect	128	262	129	263
rect	128	265	129	266
rect	128	268	129	269
rect	128	274	129	275
rect	128	277	129	278
rect	128	289	129	290
rect	128	307	129	308
rect	128	310	129	311
rect	129	13	130	14
rect	129	22	130	23
rect	129	25	130	26
rect	129	28	130	29
rect	129	31	130	32
rect	129	40	130	41
rect	129	43	130	44
rect	129	46	130	47
rect	129	55	130	56
rect	129	58	130	59
rect	129	61	130	62
rect	129	76	130	77
rect	129	85	130	86
rect	129	91	130	92
rect	129	103	130	104
rect	129	109	130	110
rect	129	112	130	113
rect	129	115	130	116
rect	129	118	130	119
rect	129	121	130	122
rect	129	127	130	128
rect	129	142	130	143
rect	129	145	130	146
rect	129	148	130	149
rect	129	151	130	152
rect	129	154	130	155
rect	129	157	130	158
rect	129	160	130	161
rect	129	166	130	167
rect	129	181	130	182
rect	129	184	130	185
rect	129	187	130	188
rect	129	196	130	197
rect	129	205	130	206
rect	129	208	130	209
rect	129	211	130	212
rect	129	217	130	218
rect	129	223	130	224
rect	129	229	130	230
rect	129	232	130	233
rect	129	235	130	236
rect	129	244	130	245
rect	129	247	130	248
rect	129	250	130	251
rect	129	256	130	257
rect	129	262	130	263
rect	129	265	130	266
rect	129	268	130	269
rect	129	274	130	275
rect	129	277	130	278
rect	129	289	130	290
rect	129	307	130	308
rect	129	310	130	311
rect	130	13	131	14
rect	130	22	131	23
rect	130	25	131	26
rect	130	28	131	29
rect	130	31	131	32
rect	130	40	131	41
rect	130	43	131	44
rect	130	46	131	47
rect	130	55	131	56
rect	130	58	131	59
rect	130	61	131	62
rect	130	76	131	77
rect	130	85	131	86
rect	130	88	131	89
rect	130	91	131	92
rect	130	103	131	104
rect	130	106	131	107
rect	130	109	131	110
rect	130	112	131	113
rect	130	115	131	116
rect	130	118	131	119
rect	130	121	131	122
rect	130	127	131	128
rect	130	139	131	140
rect	130	142	131	143
rect	130	145	131	146
rect	130	148	131	149
rect	130	151	131	152
rect	130	154	131	155
rect	130	157	131	158
rect	130	160	131	161
rect	130	166	131	167
rect	130	175	131	176
rect	130	181	131	182
rect	130	184	131	185
rect	130	187	131	188
rect	130	196	131	197
rect	130	205	131	206
rect	130	208	131	209
rect	130	211	131	212
rect	130	214	131	215
rect	130	217	131	218
rect	130	223	131	224
rect	130	229	131	230
rect	130	232	131	233
rect	130	235	131	236
rect	130	244	131	245
rect	130	247	131	248
rect	130	250	131	251
rect	130	256	131	257
rect	130	259	131	260
rect	130	262	131	263
rect	130	265	131	266
rect	130	268	131	269
rect	130	274	131	275
rect	130	277	131	278
rect	130	289	131	290
rect	130	307	131	308
rect	130	310	131	311
rect	131	13	132	14
rect	131	22	132	23
rect	131	25	132	26
rect	131	28	132	29
rect	131	40	132	41
rect	131	43	132	44
rect	131	55	132	56
rect	131	58	132	59
rect	131	61	132	62
rect	131	76	132	77
rect	131	85	132	86
rect	131	88	132	89
rect	131	91	132	92
rect	131	103	132	104
rect	131	106	132	107
rect	131	109	132	110
rect	131	112	132	113
rect	131	115	132	116
rect	131	118	132	119
rect	131	121	132	122
rect	131	127	132	128
rect	131	139	132	140
rect	131	142	132	143
rect	131	145	132	146
rect	131	148	132	149
rect	131	151	132	152
rect	131	154	132	155
rect	131	157	132	158
rect	131	160	132	161
rect	131	166	132	167
rect	131	175	132	176
rect	131	181	132	182
rect	131	184	132	185
rect	131	187	132	188
rect	131	196	132	197
rect	131	205	132	206
rect	131	208	132	209
rect	131	211	132	212
rect	131	214	132	215
rect	131	217	132	218
rect	131	223	132	224
rect	131	229	132	230
rect	131	232	132	233
rect	131	235	132	236
rect	131	244	132	245
rect	131	247	132	248
rect	131	250	132	251
rect	131	256	132	257
rect	131	259	132	260
rect	131	262	132	263
rect	131	265	132	266
rect	131	268	132	269
rect	131	274	132	275
rect	131	277	132	278
rect	131	289	132	290
rect	131	307	132	308
rect	131	310	132	311
rect	132	13	133	14
rect	132	22	133	23
rect	132	25	133	26
rect	132	28	133	29
rect	132	37	133	38
rect	132	40	133	41
rect	132	43	133	44
rect	132	52	133	53
rect	132	55	133	56
rect	132	58	133	59
rect	132	61	133	62
rect	132	64	133	65
rect	132	76	133	77
rect	132	85	133	86
rect	132	88	133	89
rect	132	91	133	92
rect	132	103	133	104
rect	132	106	133	107
rect	132	109	133	110
rect	132	112	133	113
rect	132	115	133	116
rect	132	118	133	119
rect	132	121	133	122
rect	132	127	133	128
rect	132	139	133	140
rect	132	142	133	143
rect	132	145	133	146
rect	132	148	133	149
rect	132	151	133	152
rect	132	154	133	155
rect	132	157	133	158
rect	132	160	133	161
rect	132	166	133	167
rect	132	175	133	176
rect	132	181	133	182
rect	132	184	133	185
rect	132	187	133	188
rect	132	196	133	197
rect	132	205	133	206
rect	132	208	133	209
rect	132	211	133	212
rect	132	214	133	215
rect	132	217	133	218
rect	132	223	133	224
rect	132	229	133	230
rect	132	232	133	233
rect	132	235	133	236
rect	132	244	133	245
rect	132	247	133	248
rect	132	250	133	251
rect	132	256	133	257
rect	132	259	133	260
rect	132	262	133	263
rect	132	265	133	266
rect	132	268	133	269
rect	132	274	133	275
rect	132	277	133	278
rect	132	286	133	287
rect	132	289	133	290
rect	132	307	133	308
rect	132	310	133	311
rect	133	13	134	14
rect	133	22	134	23
rect	133	25	134	26
rect	133	37	134	38
rect	133	40	134	41
rect	133	52	134	53
rect	133	55	134	56
rect	133	58	134	59
rect	133	64	134	65
rect	133	76	134	77
rect	133	85	134	86
rect	133	88	134	89
rect	133	91	134	92
rect	133	103	134	104
rect	133	106	134	107
rect	133	109	134	110
rect	133	112	134	113
rect	133	115	134	116
rect	133	118	134	119
rect	133	121	134	122
rect	133	139	134	140
rect	133	142	134	143
rect	133	145	134	146
rect	133	148	134	149
rect	133	151	134	152
rect	133	154	134	155
rect	133	157	134	158
rect	133	166	134	167
rect	133	175	134	176
rect	133	181	134	182
rect	133	184	134	185
rect	133	187	134	188
rect	133	196	134	197
rect	133	205	134	206
rect	133	208	134	209
rect	133	214	134	215
rect	133	217	134	218
rect	133	223	134	224
rect	133	232	134	233
rect	133	235	134	236
rect	133	244	134	245
rect	133	247	134	248
rect	133	250	134	251
rect	133	256	134	257
rect	133	259	134	260
rect	133	262	134	263
rect	133	265	134	266
rect	133	268	134	269
rect	133	274	134	275
rect	133	277	134	278
rect	133	286	134	287
rect	133	289	134	290
rect	133	307	134	308
rect	134	13	135	14
rect	134	22	135	23
rect	134	25	135	26
rect	134	34	135	35
rect	134	37	135	38
rect	134	40	135	41
rect	134	49	135	50
rect	134	52	135	53
rect	134	55	135	56
rect	134	58	135	59
rect	134	64	135	65
rect	134	73	135	74
rect	134	76	135	77
rect	134	85	135	86
rect	134	88	135	89
rect	134	91	135	92
rect	134	94	135	95
rect	134	97	135	98
rect	134	103	135	104
rect	134	106	135	107
rect	134	109	135	110
rect	134	112	135	113
rect	134	115	135	116
rect	134	118	135	119
rect	134	121	135	122
rect	134	136	135	137
rect	134	139	135	140
rect	134	142	135	143
rect	134	145	135	146
rect	134	148	135	149
rect	134	151	135	152
rect	134	154	135	155
rect	134	157	135	158
rect	134	166	135	167
rect	134	175	135	176
rect	134	178	135	179
rect	134	181	135	182
rect	134	184	135	185
rect	134	187	135	188
rect	134	196	135	197
rect	134	205	135	206
rect	134	208	135	209
rect	134	214	135	215
rect	134	217	135	218
rect	134	220	135	221
rect	134	223	135	224
rect	134	232	135	233
rect	134	235	135	236
rect	134	244	135	245
rect	134	247	135	248
rect	134	250	135	251
rect	134	253	135	254
rect	134	256	135	257
rect	134	259	135	260
rect	134	262	135	263
rect	134	265	135	266
rect	134	268	135	269
rect	134	274	135	275
rect	134	277	135	278
rect	134	286	135	287
rect	134	289	135	290
rect	134	307	135	308
rect	134	316	135	317
rect	135	22	136	23
rect	135	34	136	35
rect	135	37	136	38
rect	135	49	136	50
rect	135	52	136	53
rect	135	55	136	56
rect	135	58	136	59
rect	135	64	136	65
rect	135	73	136	74
rect	135	76	136	77
rect	135	85	136	86
rect	135	88	136	89
rect	135	91	136	92
rect	135	94	136	95
rect	135	97	136	98
rect	135	103	136	104
rect	135	106	136	107
rect	135	109	136	110
rect	135	112	136	113
rect	135	115	136	116
rect	135	118	136	119
rect	135	121	136	122
rect	135	136	136	137
rect	135	139	136	140
rect	135	142	136	143
rect	135	145	136	146
rect	135	148	136	149
rect	135	151	136	152
rect	135	154	136	155
rect	135	157	136	158
rect	135	166	136	167
rect	135	175	136	176
rect	135	178	136	179
rect	135	181	136	182
rect	135	184	136	185
rect	135	187	136	188
rect	135	196	136	197
rect	135	205	136	206
rect	135	208	136	209
rect	135	214	136	215
rect	135	217	136	218
rect	135	220	136	221
rect	135	223	136	224
rect	135	232	136	233
rect	135	235	136	236
rect	135	244	136	245
rect	135	247	136	248
rect	135	250	136	251
rect	135	253	136	254
rect	135	256	136	257
rect	135	259	136	260
rect	135	262	136	263
rect	135	265	136	266
rect	135	268	136	269
rect	135	274	136	275
rect	135	277	136	278
rect	135	286	136	287
rect	135	289	136	290
rect	135	316	136	317
rect	136	16	137	17
rect	136	22	137	23
rect	136	31	137	32
rect	136	34	137	35
rect	136	37	137	38
rect	136	46	137	47
rect	136	49	137	50
rect	136	52	137	53
rect	136	55	137	56
rect	136	58	137	59
rect	136	61	137	62
rect	136	64	137	65
rect	136	73	137	74
rect	136	76	137	77
rect	136	85	137	86
rect	136	88	137	89
rect	136	91	137	92
rect	136	94	137	95
rect	136	97	137	98
rect	136	103	137	104
rect	136	106	137	107
rect	136	109	137	110
rect	136	112	137	113
rect	136	115	137	116
rect	136	118	137	119
rect	136	121	137	122
rect	136	136	137	137
rect	136	139	137	140
rect	136	142	137	143
rect	136	145	137	146
rect	136	148	137	149
rect	136	151	137	152
rect	136	154	137	155
rect	136	157	137	158
rect	136	166	137	167
rect	136	175	137	176
rect	136	178	137	179
rect	136	181	137	182
rect	136	184	137	185
rect	136	187	137	188
rect	136	196	137	197
rect	136	205	137	206
rect	136	208	137	209
rect	136	214	137	215
rect	136	217	137	218
rect	136	220	137	221
rect	136	223	137	224
rect	136	232	137	233
rect	136	235	137	236
rect	136	244	137	245
rect	136	247	137	248
rect	136	250	137	251
rect	136	253	137	254
rect	136	256	137	257
rect	136	259	137	260
rect	136	262	137	263
rect	136	265	137	266
rect	136	268	137	269
rect	136	271	137	272
rect	136	274	137	275
rect	136	277	137	278
rect	136	286	137	287
rect	136	289	137	290
rect	136	298	137	299
rect	136	301	137	302
rect	136	313	137	314
rect	136	316	137	317
rect	137	16	138	17
rect	137	31	138	32
rect	137	34	138	35
rect	137	37	138	38
rect	137	46	138	47
rect	137	49	138	50
rect	137	52	138	53
rect	137	55	138	56
rect	137	58	138	59
rect	137	61	138	62
rect	137	64	138	65
rect	137	73	138	74
rect	137	76	138	77
rect	137	85	138	86
rect	137	88	138	89
rect	137	91	138	92
rect	137	94	138	95
rect	137	97	138	98
rect	137	103	138	104
rect	137	106	138	107
rect	137	109	138	110
rect	137	112	138	113
rect	137	115	138	116
rect	137	118	138	119
rect	137	121	138	122
rect	137	136	138	137
rect	137	139	138	140
rect	137	142	138	143
rect	137	145	138	146
rect	137	148	138	149
rect	137	151	138	152
rect	137	154	138	155
rect	137	157	138	158
rect	137	166	138	167
rect	137	175	138	176
rect	137	178	138	179
rect	137	181	138	182
rect	137	184	138	185
rect	137	187	138	188
rect	137	196	138	197
rect	137	205	138	206
rect	137	208	138	209
rect	137	214	138	215
rect	137	217	138	218
rect	137	220	138	221
rect	137	223	138	224
rect	137	232	138	233
rect	137	235	138	236
rect	137	244	138	245
rect	137	247	138	248
rect	137	250	138	251
rect	137	253	138	254
rect	137	256	138	257
rect	137	259	138	260
rect	137	262	138	263
rect	137	268	138	269
rect	137	271	138	272
rect	137	274	138	275
rect	137	277	138	278
rect	137	286	138	287
rect	137	289	138	290
rect	137	298	138	299
rect	137	301	138	302
rect	137	313	138	314
rect	137	316	138	317
rect	138	10	139	11
rect	138	13	139	14
rect	138	16	139	17
rect	138	31	139	32
rect	138	34	139	35
rect	138	37	139	38
rect	138	46	139	47
rect	138	49	139	50
rect	138	52	139	53
rect	138	55	139	56
rect	138	58	139	59
rect	138	61	139	62
rect	138	64	139	65
rect	138	73	139	74
rect	138	76	139	77
rect	138	85	139	86
rect	138	88	139	89
rect	138	91	139	92
rect	138	94	139	95
rect	138	97	139	98
rect	138	103	139	104
rect	138	106	139	107
rect	138	109	139	110
rect	138	112	139	113
rect	138	115	139	116
rect	138	118	139	119
rect	138	121	139	122
rect	138	136	139	137
rect	138	139	139	140
rect	138	142	139	143
rect	138	145	139	146
rect	138	148	139	149
rect	138	151	139	152
rect	138	154	139	155
rect	138	157	139	158
rect	138	166	139	167
rect	138	175	139	176
rect	138	178	139	179
rect	138	181	139	182
rect	138	184	139	185
rect	138	187	139	188
rect	138	196	139	197
rect	138	205	139	206
rect	138	208	139	209
rect	138	214	139	215
rect	138	217	139	218
rect	138	220	139	221
rect	138	223	139	224
rect	138	232	139	233
rect	138	235	139	236
rect	138	244	139	245
rect	138	247	139	248
rect	138	250	139	251
rect	138	253	139	254
rect	138	256	139	257
rect	138	259	139	260
rect	138	262	139	263
rect	138	268	139	269
rect	138	271	139	272
rect	138	274	139	275
rect	138	277	139	278
rect	138	286	139	287
rect	138	289	139	290
rect	138	292	139	293
rect	138	298	139	299
rect	138	301	139	302
rect	138	310	139	311
rect	138	313	139	314
rect	138	316	139	317
rect	145	10	146	11
rect	145	13	146	14
rect	145	16	146	17
rect	145	19	146	20
rect	145	25	146	26
rect	145	31	146	32
rect	145	34	146	35
rect	145	37	146	38
rect	145	46	146	47
rect	145	49	146	50
rect	145	52	146	53
rect	145	55	146	56
rect	145	58	146	59
rect	145	61	146	62
rect	145	73	146	74
rect	145	76	146	77
rect	145	85	146	86
rect	145	88	146	89
rect	145	91	146	92
rect	145	94	146	95
rect	145	103	146	104
rect	145	106	146	107
rect	145	109	146	110
rect	145	118	146	119
rect	145	121	146	122
rect	145	127	146	128
rect	145	136	146	137
rect	145	139	146	140
rect	145	142	146	143
rect	145	145	146	146
rect	145	148	146	149
rect	145	151	146	152
rect	145	154	146	155
rect	145	157	146	158
rect	145	166	146	167
rect	145	175	146	176
rect	145	178	146	179
rect	145	181	146	182
rect	145	184	146	185
rect	145	187	146	188
rect	145	196	146	197
rect	145	199	146	200
rect	145	205	146	206
rect	145	208	146	209
rect	145	214	146	215
rect	145	217	146	218
rect	145	220	146	221
rect	145	223	146	224
rect	145	232	146	233
rect	145	235	146	236
rect	145	244	146	245
rect	145	247	146	248
rect	145	250	146	251
rect	145	253	146	254
rect	145	256	146	257
rect	145	259	146	260
rect	145	262	146	263
rect	145	271	146	272
rect	145	274	146	275
rect	145	277	146	278
rect	145	283	146	284
rect	145	286	146	287
rect	145	289	146	290
rect	145	292	146	293
rect	145	298	146	299
rect	145	307	146	308
rect	145	310	146	311
rect	145	313	146	314
rect	145	316	146	317
rect	146	10	147	11
rect	146	13	147	14
rect	146	16	147	17
rect	146	19	147	20
rect	146	25	147	26
rect	146	31	147	32
rect	146	34	147	35
rect	146	37	147	38
rect	146	46	147	47
rect	146	49	147	50
rect	146	52	147	53
rect	146	55	147	56
rect	146	58	147	59
rect	146	61	147	62
rect	146	73	147	74
rect	146	76	147	77
rect	146	85	147	86
rect	146	88	147	89
rect	146	91	147	92
rect	146	94	147	95
rect	146	103	147	104
rect	146	106	147	107
rect	146	109	147	110
rect	146	118	147	119
rect	146	121	147	122
rect	146	127	147	128
rect	146	136	147	137
rect	146	139	147	140
rect	146	142	147	143
rect	146	145	147	146
rect	146	148	147	149
rect	146	151	147	152
rect	146	154	147	155
rect	146	166	147	167
rect	146	175	147	176
rect	146	178	147	179
rect	146	181	147	182
rect	146	184	147	185
rect	146	187	147	188
rect	146	196	147	197
rect	146	199	147	200
rect	146	205	147	206
rect	146	208	147	209
rect	146	214	147	215
rect	146	217	147	218
rect	146	220	147	221
rect	146	223	147	224
rect	146	232	147	233
rect	146	235	147	236
rect	146	244	147	245
rect	146	247	147	248
rect	146	250	147	251
rect	146	253	147	254
rect	146	256	147	257
rect	146	259	147	260
rect	146	262	147	263
rect	146	271	147	272
rect	146	274	147	275
rect	146	277	147	278
rect	146	283	147	284
rect	146	286	147	287
rect	146	289	147	290
rect	146	292	147	293
rect	146	298	147	299
rect	146	307	147	308
rect	146	310	147	311
rect	146	313	147	314
rect	146	316	147	317
rect	147	10	148	11
rect	147	13	148	14
rect	147	16	148	17
rect	147	19	148	20
rect	147	25	148	26
rect	147	31	148	32
rect	147	34	148	35
rect	147	37	148	38
rect	147	46	148	47
rect	147	49	148	50
rect	147	52	148	53
rect	147	55	148	56
rect	147	58	148	59
rect	147	61	148	62
rect	147	73	148	74
rect	147	76	148	77
rect	147	85	148	86
rect	147	88	148	89
rect	147	91	148	92
rect	147	94	148	95
rect	147	103	148	104
rect	147	106	148	107
rect	147	109	148	110
rect	147	118	148	119
rect	147	121	148	122
rect	147	127	148	128
rect	147	130	148	131
rect	147	136	148	137
rect	147	139	148	140
rect	147	142	148	143
rect	147	145	148	146
rect	147	148	148	149
rect	147	151	148	152
rect	147	154	148	155
rect	147	166	148	167
rect	147	175	148	176
rect	147	178	148	179
rect	147	181	148	182
rect	147	184	148	185
rect	147	187	148	188
rect	147	196	148	197
rect	147	199	148	200
rect	147	205	148	206
rect	147	208	148	209
rect	147	214	148	215
rect	147	217	148	218
rect	147	220	148	221
rect	147	223	148	224
rect	147	232	148	233
rect	147	235	148	236
rect	147	244	148	245
rect	147	247	148	248
rect	147	250	148	251
rect	147	253	148	254
rect	147	256	148	257
rect	147	259	148	260
rect	147	262	148	263
rect	147	271	148	272
rect	147	274	148	275
rect	147	277	148	278
rect	147	283	148	284
rect	147	286	148	287
rect	147	289	148	290
rect	147	292	148	293
rect	147	298	148	299
rect	147	307	148	308
rect	147	310	148	311
rect	147	313	148	314
rect	147	316	148	317
rect	148	10	149	11
rect	148	13	149	14
rect	148	16	149	17
rect	148	19	149	20
rect	148	25	149	26
rect	148	31	149	32
rect	148	34	149	35
rect	148	37	149	38
rect	148	46	149	47
rect	148	49	149	50
rect	148	52	149	53
rect	148	55	149	56
rect	148	58	149	59
rect	148	61	149	62
rect	148	73	149	74
rect	148	76	149	77
rect	148	85	149	86
rect	148	88	149	89
rect	148	91	149	92
rect	148	94	149	95
rect	148	103	149	104
rect	148	106	149	107
rect	148	109	149	110
rect	148	118	149	119
rect	148	121	149	122
rect	148	127	149	128
rect	148	130	149	131
rect	148	136	149	137
rect	148	139	149	140
rect	148	142	149	143
rect	148	145	149	146
rect	148	148	149	149
rect	148	154	149	155
rect	148	166	149	167
rect	148	175	149	176
rect	148	178	149	179
rect	148	181	149	182
rect	148	184	149	185
rect	148	187	149	188
rect	148	196	149	197
rect	148	199	149	200
rect	148	205	149	206
rect	148	208	149	209
rect	148	214	149	215
rect	148	217	149	218
rect	148	220	149	221
rect	148	223	149	224
rect	148	232	149	233
rect	148	235	149	236
rect	148	244	149	245
rect	148	247	149	248
rect	148	250	149	251
rect	148	253	149	254
rect	148	256	149	257
rect	148	259	149	260
rect	148	262	149	263
rect	148	271	149	272
rect	148	274	149	275
rect	148	277	149	278
rect	148	283	149	284
rect	148	286	149	287
rect	148	289	149	290
rect	148	292	149	293
rect	148	298	149	299
rect	148	307	149	308
rect	148	310	149	311
rect	148	313	149	314
rect	148	316	149	317
rect	149	10	150	11
rect	149	13	150	14
rect	149	16	150	17
rect	149	19	150	20
rect	149	25	150	26
rect	149	31	150	32
rect	149	34	150	35
rect	149	37	150	38
rect	149	46	150	47
rect	149	49	150	50
rect	149	52	150	53
rect	149	55	150	56
rect	149	58	150	59
rect	149	61	150	62
rect	149	73	150	74
rect	149	76	150	77
rect	149	85	150	86
rect	149	88	150	89
rect	149	91	150	92
rect	149	94	150	95
rect	149	103	150	104
rect	149	106	150	107
rect	149	109	150	110
rect	149	118	150	119
rect	149	121	150	122
rect	149	127	150	128
rect	149	130	150	131
rect	149	136	150	137
rect	149	139	150	140
rect	149	142	150	143
rect	149	145	150	146
rect	149	148	150	149
rect	149	154	150	155
rect	149	157	150	158
rect	149	166	150	167
rect	149	175	150	176
rect	149	178	150	179
rect	149	181	150	182
rect	149	184	150	185
rect	149	187	150	188
rect	149	196	150	197
rect	149	199	150	200
rect	149	205	150	206
rect	149	208	150	209
rect	149	214	150	215
rect	149	217	150	218
rect	149	220	150	221
rect	149	223	150	224
rect	149	232	150	233
rect	149	235	150	236
rect	149	244	150	245
rect	149	247	150	248
rect	149	250	150	251
rect	149	253	150	254
rect	149	256	150	257
rect	149	259	150	260
rect	149	262	150	263
rect	149	271	150	272
rect	149	274	150	275
rect	149	277	150	278
rect	149	283	150	284
rect	149	286	150	287
rect	149	289	150	290
rect	149	292	150	293
rect	149	298	150	299
rect	149	307	150	308
rect	149	310	150	311
rect	149	313	150	314
rect	149	316	150	317
rect	150	10	151	11
rect	150	13	151	14
rect	150	16	151	17
rect	150	19	151	20
rect	150	25	151	26
rect	150	31	151	32
rect	150	34	151	35
rect	150	37	151	38
rect	150	46	151	47
rect	150	49	151	50
rect	150	52	151	53
rect	150	55	151	56
rect	150	58	151	59
rect	150	61	151	62
rect	150	73	151	74
rect	150	76	151	77
rect	150	85	151	86
rect	150	88	151	89
rect	150	91	151	92
rect	150	94	151	95
rect	150	103	151	104
rect	150	106	151	107
rect	150	109	151	110
rect	150	118	151	119
rect	150	121	151	122
rect	150	127	151	128
rect	150	130	151	131
rect	150	136	151	137
rect	150	139	151	140
rect	150	145	151	146
rect	150	148	151	149
rect	150	154	151	155
rect	150	157	151	158
rect	150	166	151	167
rect	150	175	151	176
rect	150	178	151	179
rect	150	181	151	182
rect	150	184	151	185
rect	150	187	151	188
rect	150	196	151	197
rect	150	199	151	200
rect	150	205	151	206
rect	150	208	151	209
rect	150	214	151	215
rect	150	217	151	218
rect	150	220	151	221
rect	150	223	151	224
rect	150	232	151	233
rect	150	235	151	236
rect	150	244	151	245
rect	150	247	151	248
rect	150	250	151	251
rect	150	253	151	254
rect	150	256	151	257
rect	150	259	151	260
rect	150	262	151	263
rect	150	271	151	272
rect	150	274	151	275
rect	150	277	151	278
rect	150	283	151	284
rect	150	286	151	287
rect	150	289	151	290
rect	150	292	151	293
rect	150	298	151	299
rect	150	307	151	308
rect	150	310	151	311
rect	150	313	151	314
rect	150	316	151	317
rect	151	10	152	11
rect	151	13	152	14
rect	151	16	152	17
rect	151	19	152	20
rect	151	25	152	26
rect	151	31	152	32
rect	151	34	152	35
rect	151	37	152	38
rect	151	46	152	47
rect	151	49	152	50
rect	151	52	152	53
rect	151	55	152	56
rect	151	58	152	59
rect	151	61	152	62
rect	151	73	152	74
rect	151	76	152	77
rect	151	85	152	86
rect	151	88	152	89
rect	151	91	152	92
rect	151	94	152	95
rect	151	103	152	104
rect	151	106	152	107
rect	151	109	152	110
rect	151	118	152	119
rect	151	121	152	122
rect	151	127	152	128
rect	151	130	152	131
rect	151	136	152	137
rect	151	139	152	140
rect	151	145	152	146
rect	151	148	152	149
rect	151	151	152	152
rect	151	154	152	155
rect	151	157	152	158
rect	151	166	152	167
rect	151	175	152	176
rect	151	178	152	179
rect	151	181	152	182
rect	151	184	152	185
rect	151	187	152	188
rect	151	196	152	197
rect	151	199	152	200
rect	151	205	152	206
rect	151	208	152	209
rect	151	214	152	215
rect	151	217	152	218
rect	151	220	152	221
rect	151	223	152	224
rect	151	232	152	233
rect	151	235	152	236
rect	151	244	152	245
rect	151	247	152	248
rect	151	250	152	251
rect	151	253	152	254
rect	151	256	152	257
rect	151	259	152	260
rect	151	262	152	263
rect	151	271	152	272
rect	151	274	152	275
rect	151	277	152	278
rect	151	283	152	284
rect	151	286	152	287
rect	151	289	152	290
rect	151	292	152	293
rect	151	298	152	299
rect	151	307	152	308
rect	151	310	152	311
rect	151	313	152	314
rect	151	316	152	317
rect	152	10	153	11
rect	152	13	153	14
rect	152	16	153	17
rect	152	19	153	20
rect	152	25	153	26
rect	152	31	153	32
rect	152	34	153	35
rect	152	37	153	38
rect	152	46	153	47
rect	152	49	153	50
rect	152	52	153	53
rect	152	55	153	56
rect	152	58	153	59
rect	152	61	153	62
rect	152	73	153	74
rect	152	76	153	77
rect	152	85	153	86
rect	152	88	153	89
rect	152	91	153	92
rect	152	94	153	95
rect	152	103	153	104
rect	152	106	153	107
rect	152	109	153	110
rect	152	118	153	119
rect	152	121	153	122
rect	152	130	153	131
rect	152	136	153	137
rect	152	139	153	140
rect	152	145	153	146
rect	152	148	153	149
rect	152	151	153	152
rect	152	154	153	155
rect	152	157	153	158
rect	152	166	153	167
rect	152	175	153	176
rect	152	178	153	179
rect	152	181	153	182
rect	152	184	153	185
rect	152	187	153	188
rect	152	196	153	197
rect	152	199	153	200
rect	152	205	153	206
rect	152	208	153	209
rect	152	214	153	215
rect	152	217	153	218
rect	152	220	153	221
rect	152	223	153	224
rect	152	232	153	233
rect	152	235	153	236
rect	152	244	153	245
rect	152	247	153	248
rect	152	250	153	251
rect	152	253	153	254
rect	152	256	153	257
rect	152	259	153	260
rect	152	262	153	263
rect	152	271	153	272
rect	152	274	153	275
rect	152	277	153	278
rect	152	283	153	284
rect	152	289	153	290
rect	152	298	153	299
rect	152	307	153	308
rect	152	310	153	311
rect	152	313	153	314
rect	152	316	153	317
rect	153	10	154	11
rect	153	13	154	14
rect	153	16	154	17
rect	153	19	154	20
rect	153	25	154	26
rect	153	31	154	32
rect	153	34	154	35
rect	153	37	154	38
rect	153	46	154	47
rect	153	49	154	50
rect	153	52	154	53
rect	153	55	154	56
rect	153	58	154	59
rect	153	61	154	62
rect	153	73	154	74
rect	153	76	154	77
rect	153	85	154	86
rect	153	88	154	89
rect	153	91	154	92
rect	153	94	154	95
rect	153	103	154	104
rect	153	106	154	107
rect	153	109	154	110
rect	153	118	154	119
rect	153	121	154	122
rect	153	130	154	131
rect	153	136	154	137
rect	153	139	154	140
rect	153	142	154	143
rect	153	145	154	146
rect	153	148	154	149
rect	153	151	154	152
rect	153	154	154	155
rect	153	157	154	158
rect	153	166	154	167
rect	153	175	154	176
rect	153	178	154	179
rect	153	181	154	182
rect	153	184	154	185
rect	153	187	154	188
rect	153	196	154	197
rect	153	199	154	200
rect	153	205	154	206
rect	153	208	154	209
rect	153	214	154	215
rect	153	217	154	218
rect	153	220	154	221
rect	153	223	154	224
rect	153	232	154	233
rect	153	235	154	236
rect	153	244	154	245
rect	153	247	154	248
rect	153	250	154	251
rect	153	253	154	254
rect	153	256	154	257
rect	153	259	154	260
rect	153	262	154	263
rect	153	271	154	272
rect	153	274	154	275
rect	153	277	154	278
rect	153	283	154	284
rect	153	289	154	290
rect	153	298	154	299
rect	153	307	154	308
rect	153	310	154	311
rect	153	313	154	314
rect	153	316	154	317
rect	154	10	155	11
rect	154	13	155	14
rect	154	16	155	17
rect	154	19	155	20
rect	154	25	155	26
rect	154	31	155	32
rect	154	34	155	35
rect	154	37	155	38
rect	154	46	155	47
rect	154	49	155	50
rect	154	52	155	53
rect	154	55	155	56
rect	154	58	155	59
rect	154	73	155	74
rect	154	76	155	77
rect	154	85	155	86
rect	154	88	155	89
rect	154	91	155	92
rect	154	94	155	95
rect	154	103	155	104
rect	154	109	155	110
rect	154	118	155	119
rect	154	121	155	122
rect	154	130	155	131
rect	154	136	155	137
rect	154	139	155	140
rect	154	142	155	143
rect	154	145	155	146
rect	154	148	155	149
rect	154	151	155	152
rect	154	154	155	155
rect	154	157	155	158
rect	154	166	155	167
rect	154	175	155	176
rect	154	178	155	179
rect	154	181	155	182
rect	154	184	155	185
rect	154	187	155	188
rect	154	196	155	197
rect	154	199	155	200
rect	154	205	155	206
rect	154	208	155	209
rect	154	214	155	215
rect	154	217	155	218
rect	154	220	155	221
rect	154	223	155	224
rect	154	232	155	233
rect	154	235	155	236
rect	154	244	155	245
rect	154	247	155	248
rect	154	250	155	251
rect	154	253	155	254
rect	154	256	155	257
rect	154	259	155	260
rect	154	262	155	263
rect	154	271	155	272
rect	154	274	155	275
rect	154	283	155	284
rect	154	289	155	290
rect	154	298	155	299
rect	154	307	155	308
rect	154	310	155	311
rect	154	313	155	314
rect	154	316	155	317
rect	155	10	156	11
rect	155	13	156	14
rect	155	16	156	17
rect	155	19	156	20
rect	155	25	156	26
rect	155	31	156	32
rect	155	34	156	35
rect	155	37	156	38
rect	155	46	156	47
rect	155	49	156	50
rect	155	52	156	53
rect	155	55	156	56
rect	155	58	156	59
rect	155	70	156	71
rect	155	73	156	74
rect	155	76	156	77
rect	155	85	156	86
rect	155	88	156	89
rect	155	91	156	92
rect	155	94	156	95
rect	155	103	156	104
rect	155	109	156	110
rect	155	118	156	119
rect	155	121	156	122
rect	155	127	156	128
rect	155	130	156	131
rect	155	136	156	137
rect	155	139	156	140
rect	155	142	156	143
rect	155	145	156	146
rect	155	148	156	149
rect	155	151	156	152
rect	155	154	156	155
rect	155	157	156	158
rect	155	166	156	167
rect	155	175	156	176
rect	155	178	156	179
rect	155	181	156	182
rect	155	184	156	185
rect	155	187	156	188
rect	155	196	156	197
rect	155	199	156	200
rect	155	205	156	206
rect	155	208	156	209
rect	155	214	156	215
rect	155	217	156	218
rect	155	220	156	221
rect	155	223	156	224
rect	155	232	156	233
rect	155	235	156	236
rect	155	244	156	245
rect	155	247	156	248
rect	155	250	156	251
rect	155	253	156	254
rect	155	256	156	257
rect	155	259	156	260
rect	155	262	156	263
rect	155	271	156	272
rect	155	274	156	275
rect	155	283	156	284
rect	155	289	156	290
rect	155	292	156	293
rect	155	298	156	299
rect	155	307	156	308
rect	155	310	156	311
rect	155	313	156	314
rect	155	316	156	317
rect	156	10	157	11
rect	156	13	157	14
rect	156	16	157	17
rect	156	19	157	20
rect	156	25	157	26
rect	156	31	157	32
rect	156	34	157	35
rect	156	37	157	38
rect	156	46	157	47
rect	156	49	157	50
rect	156	52	157	53
rect	156	55	157	56
rect	156	70	157	71
rect	156	73	157	74
rect	156	76	157	77
rect	156	85	157	86
rect	156	88	157	89
rect	156	94	157	95
rect	156	103	157	104
rect	156	109	157	110
rect	156	118	157	119
rect	156	121	157	122
rect	156	127	157	128
rect	156	130	157	131
rect	156	136	157	137
rect	156	139	157	140
rect	156	142	157	143
rect	156	145	157	146
rect	156	148	157	149
rect	156	151	157	152
rect	156	154	157	155
rect	156	157	157	158
rect	156	166	157	167
rect	156	175	157	176
rect	156	178	157	179
rect	156	181	157	182
rect	156	184	157	185
rect	156	187	157	188
rect	156	196	157	197
rect	156	199	157	200
rect	156	205	157	206
rect	156	208	157	209
rect	156	214	157	215
rect	156	217	157	218
rect	156	220	157	221
rect	156	223	157	224
rect	156	232	157	233
rect	156	235	157	236
rect	156	244	157	245
rect	156	247	157	248
rect	156	250	157	251
rect	156	253	157	254
rect	156	256	157	257
rect	156	262	157	263
rect	156	271	157	272
rect	156	274	157	275
rect	156	283	157	284
rect	156	289	157	290
rect	156	292	157	293
rect	156	298	157	299
rect	156	307	157	308
rect	156	310	157	311
rect	156	313	157	314
rect	156	316	157	317
rect	157	10	158	11
rect	157	13	158	14
rect	157	16	158	17
rect	157	19	158	20
rect	157	25	158	26
rect	157	31	158	32
rect	157	34	158	35
rect	157	37	158	38
rect	157	46	158	47
rect	157	49	158	50
rect	157	52	158	53
rect	157	55	158	56
rect	157	61	158	62
rect	157	70	158	71
rect	157	73	158	74
rect	157	76	158	77
rect	157	85	158	86
rect	157	88	158	89
rect	157	94	158	95
rect	157	103	158	104
rect	157	106	158	107
rect	157	109	158	110
rect	157	118	158	119
rect	157	121	158	122
rect	157	127	158	128
rect	157	130	158	131
rect	157	136	158	137
rect	157	139	158	140
rect	157	142	158	143
rect	157	145	158	146
rect	157	148	158	149
rect	157	151	158	152
rect	157	154	158	155
rect	157	157	158	158
rect	157	166	158	167
rect	157	175	158	176
rect	157	178	158	179
rect	157	181	158	182
rect	157	184	158	185
rect	157	187	158	188
rect	157	196	158	197
rect	157	199	158	200
rect	157	205	158	206
rect	157	208	158	209
rect	157	214	158	215
rect	157	217	158	218
rect	157	220	158	221
rect	157	223	158	224
rect	157	232	158	233
rect	157	235	158	236
rect	157	244	158	245
rect	157	247	158	248
rect	157	250	158	251
rect	157	253	158	254
rect	157	256	158	257
rect	157	262	158	263
rect	157	271	158	272
rect	157	274	158	275
rect	157	277	158	278
rect	157	283	158	284
rect	157	289	158	290
rect	157	292	158	293
rect	157	298	158	299
rect	157	307	158	308
rect	157	310	158	311
rect	157	313	158	314
rect	157	316	158	317
rect	158	10	159	11
rect	158	13	159	14
rect	158	16	159	17
rect	158	19	159	20
rect	158	25	159	26
rect	158	31	159	32
rect	158	34	159	35
rect	158	37	159	38
rect	158	46	159	47
rect	158	49	159	50
rect	158	55	159	56
rect	158	61	159	62
rect	158	70	159	71
rect	158	76	159	77
rect	158	85	159	86
rect	158	88	159	89
rect	158	94	159	95
rect	158	103	159	104
rect	158	106	159	107
rect	158	109	159	110
rect	158	118	159	119
rect	158	121	159	122
rect	158	127	159	128
rect	158	130	159	131
rect	158	136	159	137
rect	158	139	159	140
rect	158	142	159	143
rect	158	145	159	146
rect	158	148	159	149
rect	158	151	159	152
rect	158	157	159	158
rect	158	166	159	167
rect	158	175	159	176
rect	158	178	159	179
rect	158	181	159	182
rect	158	184	159	185
rect	158	187	159	188
rect	158	196	159	197
rect	158	199	159	200
rect	158	205	159	206
rect	158	208	159	209
rect	158	220	159	221
rect	158	223	159	224
rect	158	232	159	233
rect	158	235	159	236
rect	158	244	159	245
rect	158	247	159	248
rect	158	250	159	251
rect	158	256	159	257
rect	158	262	159	263
rect	158	271	159	272
rect	158	274	159	275
rect	158	277	159	278
rect	158	283	159	284
rect	158	289	159	290
rect	158	292	159	293
rect	158	298	159	299
rect	158	307	159	308
rect	158	310	159	311
rect	158	313	159	314
rect	158	316	159	317
rect	159	10	160	11
rect	159	13	160	14
rect	159	16	160	17
rect	159	19	160	20
rect	159	25	160	26
rect	159	31	160	32
rect	159	34	160	35
rect	159	37	160	38
rect	159	46	160	47
rect	159	49	160	50
rect	159	55	160	56
rect	159	58	160	59
rect	159	61	160	62
rect	159	70	160	71
rect	159	76	160	77
rect	159	85	160	86
rect	159	88	160	89
rect	159	91	160	92
rect	159	94	160	95
rect	159	103	160	104
rect	159	106	160	107
rect	159	109	160	110
rect	159	118	160	119
rect	159	121	160	122
rect	159	127	160	128
rect	159	130	160	131
rect	159	136	160	137
rect	159	139	160	140
rect	159	142	160	143
rect	159	145	160	146
rect	159	148	160	149
rect	159	151	160	152
rect	159	157	160	158
rect	159	160	160	161
rect	159	166	160	167
rect	159	175	160	176
rect	159	178	160	179
rect	159	181	160	182
rect	159	184	160	185
rect	159	187	160	188
rect	159	196	160	197
rect	159	199	160	200
rect	159	205	160	206
rect	159	208	160	209
rect	159	220	160	221
rect	159	223	160	224
rect	159	232	160	233
rect	159	235	160	236
rect	159	244	160	245
rect	159	247	160	248
rect	159	250	160	251
rect	159	256	160	257
rect	159	259	160	260
rect	159	262	160	263
rect	159	271	160	272
rect	159	274	160	275
rect	159	277	160	278
rect	159	283	160	284
rect	159	289	160	290
rect	159	292	160	293
rect	159	298	160	299
rect	159	307	160	308
rect	159	310	160	311
rect	159	313	160	314
rect	159	316	160	317
rect	160	10	161	11
rect	160	13	161	14
rect	160	16	161	17
rect	160	19	161	20
rect	160	25	161	26
rect	160	31	161	32
rect	160	37	161	38
rect	160	46	161	47
rect	160	49	161	50
rect	160	58	161	59
rect	160	61	161	62
rect	160	70	161	71
rect	160	85	161	86
rect	160	91	161	92
rect	160	94	161	95
rect	160	103	161	104
rect	160	106	161	107
rect	160	109	161	110
rect	160	118	161	119
rect	160	121	161	122
rect	160	127	161	128
rect	160	130	161	131
rect	160	136	161	137
rect	160	139	161	140
rect	160	142	161	143
rect	160	145	161	146
rect	160	151	161	152
rect	160	157	161	158
rect	160	160	161	161
rect	160	166	161	167
rect	160	178	161	179
rect	160	181	161	182
rect	160	184	161	185
rect	160	187	161	188
rect	160	196	161	197
rect	160	199	161	200
rect	160	208	161	209
rect	160	220	161	221
rect	160	223	161	224
rect	160	232	161	233
rect	160	235	161	236
rect	160	245	161	246
rect	160	246	161	247
rect	160	247	161	248
rect	160	248	161	249
rect	160	249	161	250
rect	160	250	161	251
rect	160	251	161	252
rect	160	252	161	253
rect	160	256	161	257
rect	160	259	161	260
rect	160	262	161	263
rect	160	271	161	272
rect	160	274	161	275
rect	160	277	161	278
rect	160	283	161	284
rect	160	289	161	290
rect	160	292	161	293
rect	160	298	161	299
rect	160	307	161	308
rect	160	310	161	311
rect	160	313	161	314
rect	160	316	161	317
rect	161	10	162	11
rect	161	13	162	14
rect	161	16	162	17
rect	161	19	162	20
rect	161	25	162	26
rect	161	31	162	32
rect	161	37	162	38
rect	161	40	162	41
rect	161	46	162	47
rect	161	49	162	50
rect	161	52	162	53
rect	161	58	162	59
rect	161	61	162	62
rect	161	70	162	71
rect	161	73	162	74
rect	161	83	162	84
rect	161	85	162	86
rect	161	91	162	92
rect	161	94	162	95
rect	161	103	162	104
rect	161	106	162	107
rect	161	109	162	110
rect	161	118	162	119
rect	161	121	162	122
rect	161	127	162	128
rect	161	130	162	131
rect	161	136	162	137
rect	161	139	162	140
rect	161	142	162	143
rect	161	145	162	146
rect	161	151	162	152
rect	161	154	162	155
rect	161	157	162	158
rect	161	160	162	161
rect	161	166	162	167
rect	161	172	162	173
rect	161	178	162	179
rect	161	181	162	182
rect	161	184	162	185
rect	161	187	162	188
rect	161	196	162	197
rect	161	199	162	200
rect	161	208	162	209
rect	161	214	162	215
rect	161	220	162	221
rect	161	223	162	224
rect	161	232	162	233
rect	161	235	162	236
rect	161	247	162	248
rect	161	250	162	251
rect	161	253	162	254
rect	161	256	162	257
rect	161	259	162	260
rect	161	262	162	263
rect	161	271	162	272
rect	161	274	162	275
rect	161	277	162	278
rect	161	283	162	284
rect	161	289	162	290
rect	161	292	162	293
rect	161	298	162	299
rect	161	307	162	308
rect	161	310	162	311
rect	161	313	162	314
rect	161	316	162	317
rect	162	10	163	11
rect	162	13	163	14
rect	162	16	163	17
rect	162	19	163	20
rect	162	25	163	26
rect	162	31	163	32
rect	162	37	163	38
rect	162	40	163	41
rect	162	46	163	47
rect	162	49	163	50
rect	162	52	163	53
rect	162	58	163	59
rect	162	61	163	62
rect	162	70	163	71
rect	162	73	163	74
rect	162	83	163	84
rect	162	85	163	86
rect	162	91	163	92
rect	162	94	163	95
rect	162	103	163	104
rect	162	106	163	107
rect	162	109	163	110
rect	162	118	163	119
rect	162	121	163	122
rect	162	127	163	128
rect	162	130	163	131
rect	162	136	163	137
rect	162	139	163	140
rect	162	142	163	143
rect	162	145	163	146
rect	162	151	163	152
rect	162	154	163	155
rect	162	157	163	158
rect	162	160	163	161
rect	162	172	163	173
rect	162	181	163	182
rect	162	184	163	185
rect	162	187	163	188
rect	162	196	163	197
rect	162	199	163	200
rect	162	208	163	209
rect	162	214	163	215
rect	162	223	163	224
rect	162	232	163	233
rect	162	235	163	236
rect	162	250	163	251
rect	162	253	163	254
rect	162	256	163	257
rect	162	259	163	260
rect	162	262	163	263
rect	162	271	163	272
rect	162	274	163	275
rect	162	277	163	278
rect	162	283	163	284
rect	162	289	163	290
rect	162	292	163	293
rect	162	298	163	299
rect	162	307	163	308
rect	162	310	163	311
rect	162	313	163	314
rect	162	316	163	317
rect	163	10	164	11
rect	163	13	164	14
rect	163	16	164	17
rect	163	19	164	20
rect	163	25	164	26
rect	163	31	164	32
rect	163	34	164	35
rect	163	37	164	38
rect	163	40	164	41
rect	163	46	164	47
rect	163	49	164	50
rect	163	52	164	53
rect	163	58	164	59
rect	163	61	164	62
rect	163	70	164	71
rect	163	73	164	74
rect	163	83	164	84
rect	163	85	164	86
rect	163	91	164	92
rect	163	94	164	95
rect	163	103	164	104
rect	163	106	164	107
rect	163	109	164	110
rect	163	118	164	119
rect	163	121	164	122
rect	163	127	164	128
rect	163	130	164	131
rect	163	136	164	137
rect	163	139	164	140
rect	163	142	164	143
rect	163	145	164	146
rect	163	151	164	152
rect	163	154	164	155
rect	163	157	164	158
rect	163	160	164	161
rect	163	163	164	164
rect	163	172	164	173
rect	163	175	164	176
rect	163	181	164	182
rect	163	184	164	185
rect	163	187	164	188
rect	163	196	164	197
rect	163	199	164	200
rect	163	205	164	206
rect	163	208	164	209
rect	163	214	164	215
rect	163	217	164	218
rect	163	223	164	224
rect	163	232	164	233
rect	163	235	164	236
rect	163	241	164	242
rect	163	250	164	251
rect	163	253	164	254
rect	163	256	164	257
rect	163	259	164	260
rect	163	262	164	263
rect	163	271	164	272
rect	163	274	164	275
rect	163	277	164	278
rect	163	283	164	284
rect	163	289	164	290
rect	163	292	164	293
rect	163	298	164	299
rect	163	307	164	308
rect	163	310	164	311
rect	163	313	164	314
rect	163	316	164	317
rect	164	10	165	11
rect	164	13	165	14
rect	164	16	165	17
rect	164	25	165	26
rect	164	31	165	32
rect	164	34	165	35
rect	164	37	165	38
rect	164	40	165	41
rect	164	46	165	47
rect	164	49	165	50
rect	164	52	165	53
rect	164	58	165	59
rect	164	61	165	62
rect	164	70	165	71
rect	164	73	165	74
rect	164	83	165	84
rect	164	85	165	86
rect	164	91	165	92
rect	164	94	165	95
rect	164	106	165	107
rect	164	109	165	110
rect	164	118	165	119
rect	164	121	165	122
rect	164	127	165	128
rect	164	130	165	131
rect	164	136	165	137
rect	164	142	165	143
rect	164	145	165	146
rect	164	151	165	152
rect	164	154	165	155
rect	164	157	165	158
rect	164	160	165	161
rect	164	163	165	164
rect	164	172	165	173
rect	164	175	165	176
rect	164	181	165	182
rect	164	184	165	185
rect	164	187	165	188
rect	164	196	165	197
rect	164	199	165	200
rect	164	205	165	206
rect	164	208	165	209
rect	164	214	165	215
rect	164	217	165	218
rect	164	223	165	224
rect	164	232	165	233
rect	164	235	165	236
rect	164	241	165	242
rect	164	250	165	251
rect	164	253	165	254
rect	164	256	165	257
rect	164	259	165	260
rect	164	262	165	263
rect	164	271	165	272
rect	164	274	165	275
rect	164	277	165	278
rect	164	283	165	284
rect	164	289	165	290
rect	164	292	165	293
rect	164	298	165	299
rect	164	310	165	311
rect	164	313	165	314
rect	164	316	165	317
rect	165	10	166	11
rect	165	13	166	14
rect	165	16	166	17
rect	165	25	166	26
rect	165	31	166	32
rect	165	34	166	35
rect	165	37	166	38
rect	165	40	166	41
rect	165	46	166	47
rect	165	49	166	50
rect	165	52	166	53
rect	165	58	166	59
rect	165	61	166	62
rect	165	70	166	71
rect	165	73	166	74
rect	165	76	166	77
rect	165	83	166	84
rect	165	85	166	86
rect	165	88	166	89
rect	165	91	166	92
rect	165	94	166	95
rect	165	106	166	107
rect	165	109	166	110
rect	165	118	166	119
rect	165	121	166	122
rect	165	127	166	128
rect	165	130	166	131
rect	165	136	166	137
rect	165	142	166	143
rect	165	145	166	146
rect	165	151	166	152
rect	165	154	166	155
rect	165	157	166	158
rect	165	160	166	161
rect	165	163	166	164
rect	165	172	166	173
rect	165	175	166	176
rect	165	181	166	182
rect	165	184	166	185
rect	165	187	166	188
rect	165	196	166	197
rect	165	199	166	200
rect	165	205	166	206
rect	165	208	166	209
rect	165	214	166	215
rect	165	217	166	218
rect	165	223	166	224
rect	165	232	166	233
rect	165	235	166	236
rect	165	241	166	242
rect	165	250	166	251
rect	165	253	166	254
rect	165	256	166	257
rect	165	259	166	260
rect	165	262	166	263
rect	165	271	166	272
rect	165	274	166	275
rect	165	277	166	278
rect	165	283	166	284
rect	165	289	166	290
rect	165	292	166	293
rect	165	298	166	299
rect	165	310	166	311
rect	165	313	166	314
rect	165	316	166	317
rect	166	10	167	11
rect	166	13	167	14
rect	166	25	167	26
rect	166	34	167	35
rect	166	37	167	38
rect	166	40	167	41
rect	166	46	167	47
rect	166	49	167	50
rect	166	52	167	53
rect	166	58	167	59
rect	166	61	167	62
rect	166	70	167	71
rect	166	73	167	74
rect	166	76	167	77
rect	166	83	167	84
rect	166	85	167	86
rect	166	88	167	89
rect	166	91	167	92
rect	166	94	167	95
rect	166	106	167	107
rect	166	109	167	110
rect	166	118	167	119
rect	166	121	167	122
rect	166	127	167	128
rect	166	130	167	131
rect	166	136	167	137
rect	166	142	167	143
rect	166	145	167	146
rect	166	151	167	152
rect	166	154	167	155
rect	166	157	167	158
rect	166	160	167	161
rect	166	163	167	164
rect	166	172	167	173
rect	166	175	167	176
rect	166	181	167	182
rect	166	184	167	185
rect	166	187	167	188
rect	166	196	167	197
rect	166	205	167	206
rect	166	214	167	215
rect	166	217	167	218
rect	166	223	167	224
rect	166	235	167	236
rect	166	241	167	242
rect	166	250	167	251
rect	166	253	167	254
rect	166	256	167	257
rect	166	259	167	260
rect	166	262	167	263
rect	166	271	167	272
rect	166	274	167	275
rect	166	277	167	278
rect	166	283	167	284
rect	166	292	167	293
rect	166	298	167	299
rect	166	310	167	311
rect	166	316	167	317
rect	167	10	168	11
rect	167	13	168	14
rect	167	19	168	20
rect	167	25	168	26
rect	167	34	168	35
rect	167	37	168	38
rect	167	40	168	41
rect	167	46	168	47
rect	167	49	168	50
rect	167	52	168	53
rect	167	58	168	59
rect	167	61	168	62
rect	167	70	168	71
rect	167	73	168	74
rect	167	76	168	77
rect	167	83	168	84
rect	167	85	168	86
rect	167	88	168	89
rect	167	91	168	92
rect	167	94	168	95
rect	167	106	168	107
rect	167	109	168	110
rect	167	118	168	119
rect	167	121	168	122
rect	167	127	168	128
rect	167	130	168	131
rect	167	136	168	137
rect	167	142	168	143
rect	167	145	168	146
rect	167	151	168	152
rect	167	154	168	155
rect	167	157	168	158
rect	167	160	168	161
rect	167	163	168	164
rect	167	172	168	173
rect	167	175	168	176
rect	167	181	168	182
rect	167	184	168	185
rect	167	187	168	188
rect	167	196	168	197
rect	167	205	168	206
rect	167	214	168	215
rect	167	217	168	218
rect	167	220	168	221
rect	167	223	168	224
rect	167	235	168	236
rect	167	241	168	242
rect	167	250	168	251
rect	167	253	168	254
rect	167	256	168	257
rect	167	259	168	260
rect	167	262	168	263
rect	167	265	168	266
rect	167	271	168	272
rect	167	274	168	275
rect	167	277	168	278
rect	167	283	168	284
rect	167	292	168	293
rect	167	298	168	299
rect	167	304	168	305
rect	167	310	168	311
rect	167	316	168	317
rect	167	322	168	323
rect	168	10	169	11
rect	168	19	169	20
rect	168	25	169	26
rect	168	34	169	35
rect	168	40	169	41
rect	168	46	169	47
rect	168	52	169	53
rect	168	58	169	59
rect	168	61	169	62
rect	168	70	169	71
rect	168	73	169	74
rect	168	76	169	77
rect	168	85	169	86
rect	168	88	169	89
rect	168	91	169	92
rect	168	94	169	95
rect	168	106	169	107
rect	168	109	169	110
rect	168	118	169	119
rect	168	121	169	122
rect	168	127	169	128
rect	168	130	169	131
rect	168	142	169	143
rect	168	145	169	146
rect	168	151	169	152
rect	168	154	169	155
rect	168	157	169	158
rect	168	160	169	161
rect	168	163	169	164
rect	168	172	169	173
rect	168	175	169	176
rect	168	184	169	185
rect	168	187	169	188
rect	168	196	169	197
rect	168	205	169	206
rect	168	214	169	215
rect	168	217	169	218
rect	168	220	169	221
rect	168	223	169	224
rect	168	235	169	236
rect	168	241	169	242
rect	168	253	169	254
rect	168	256	169	257
rect	168	259	169	260
rect	168	265	169	266
rect	168	271	169	272
rect	168	274	169	275
rect	168	277	169	278
rect	168	283	169	284
rect	168	292	169	293
rect	168	298	169	299
rect	168	304	169	305
rect	168	316	169	317
rect	168	322	169	323
rect	169	10	170	11
rect	169	16	170	17
rect	169	19	170	20
rect	169	25	170	26
rect	169	28	170	29
rect	169	34	170	35
rect	169	40	170	41
rect	169	46	170	47
rect	169	52	170	53
rect	169	55	170	56
rect	169	58	170	59
rect	169	61	170	62
rect	169	70	170	71
rect	169	73	170	74
rect	169	76	170	77
rect	169	85	170	86
rect	169	88	170	89
rect	169	91	170	92
rect	169	94	170	95
rect	169	103	170	104
rect	169	106	170	107
rect	169	109	170	110
rect	169	112	170	113
rect	169	115	170	116
rect	169	118	170	119
rect	169	121	170	122
rect	169	127	170	128
rect	169	130	170	131
rect	169	142	170	143
rect	169	145	170	146
rect	169	151	170	152
rect	169	154	170	155
rect	169	157	170	158
rect	169	160	170	161
rect	169	163	170	164
rect	169	172	170	173
rect	169	175	170	176
rect	169	178	170	179
rect	169	184	170	185
rect	169	187	170	188
rect	169	196	170	197
rect	169	205	170	206
rect	169	208	170	209
rect	169	214	170	215
rect	169	217	170	218
rect	169	220	170	221
rect	169	223	170	224
rect	169	229	170	230
rect	169	235	170	236
rect	169	241	170	242
rect	169	253	170	254
rect	169	256	170	257
rect	169	259	170	260
rect	169	265	170	266
rect	169	271	170	272
rect	169	274	170	275
rect	169	277	170	278
rect	169	283	170	284
rect	169	289	170	290
rect	169	292	170	293
rect	169	295	170	296
rect	169	298	170	299
rect	169	301	170	302
rect	169	304	170	305
rect	169	316	170	317
rect	169	322	170	323
rect	169	328	170	329
rect	170	16	171	17
rect	170	19	171	20
rect	170	28	171	29
rect	170	34	171	35
rect	170	40	171	41
rect	170	52	171	53
rect	170	55	171	56
rect	170	58	171	59
rect	170	61	171	62
rect	170	70	171	71
rect	170	73	171	74
rect	170	76	171	77
rect	170	85	171	86
rect	170	88	171	89
rect	170	91	171	92
rect	170	94	171	95
rect	170	103	171	104
rect	170	106	171	107
rect	170	109	171	110
rect	170	112	171	113
rect	170	115	171	116
rect	170	127	171	128
rect	170	130	171	131
rect	170	142	171	143
rect	170	151	171	152
rect	170	154	171	155
rect	170	157	171	158
rect	170	160	171	161
rect	170	163	171	164
rect	170	172	171	173
rect	170	175	171	176
rect	170	178	171	179
rect	170	184	171	185
rect	170	187	171	188
rect	170	196	171	197
rect	170	205	171	206
rect	170	208	171	209
rect	170	214	171	215
rect	170	217	171	218
rect	170	220	171	221
rect	170	229	171	230
rect	170	241	171	242
rect	170	253	171	254
rect	170	259	171	260
rect	170	265	171	266
rect	170	274	171	275
rect	170	277	171	278
rect	170	289	171	290
rect	170	292	171	293
rect	170	295	171	296
rect	170	301	171	302
rect	170	304	171	305
rect	170	322	171	323
rect	170	328	171	329
rect	171	13	172	14
rect	171	16	172	17
rect	171	19	172	20
rect	171	28	172	29
rect	171	34	172	35
rect	171	37	172	38
rect	171	40	172	41
rect	171	49	172	50
rect	171	52	172	53
rect	171	55	172	56
rect	171	58	172	59
rect	171	61	172	62
rect	171	70	172	71
rect	171	73	172	74
rect	171	76	172	77
rect	171	85	172	86
rect	171	88	172	89
rect	171	91	172	92
rect	171	94	172	95
rect	171	97	172	98
rect	171	103	172	104
rect	171	106	172	107
rect	171	109	172	110
rect	171	112	172	113
rect	171	115	172	116
rect	171	127	172	128
rect	171	130	172	131
rect	171	139	172	140
rect	171	142	172	143
rect	171	151	172	152
rect	171	154	172	155
rect	171	157	172	158
rect	171	160	172	161
rect	171	163	172	164
rect	171	172	172	173
rect	171	175	172	176
rect	171	178	172	179
rect	171	181	172	182
rect	171	184	172	185
rect	171	187	172	188
rect	171	196	172	197
rect	171	205	172	206
rect	171	208	172	209
rect	171	214	172	215
rect	171	217	172	218
rect	171	220	172	221
rect	171	229	172	230
rect	171	232	172	233
rect	171	241	172	242
rect	171	244	172	245
rect	171	253	172	254
rect	171	259	172	260
rect	171	262	172	263
rect	171	265	172	266
rect	171	274	172	275
rect	171	277	172	278
rect	171	286	172	287
rect	171	289	172	290
rect	171	292	172	293
rect	171	295	172	296
rect	171	301	172	302
rect	171	304	172	305
rect	171	307	172	308
rect	171	313	172	314
rect	171	322	172	323
rect	171	325	172	326
rect	171	328	172	329
rect	178	13	179	14
rect	178	16	179	17
rect	178	19	179	20
rect	178	28	179	29
rect	178	31	179	32
rect	178	37	179	38
rect	178	40	179	41
rect	178	49	179	50
rect	178	52	179	53
rect	178	55	179	56
rect	178	58	179	59
rect	178	61	179	62
rect	178	70	179	71
rect	178	73	179	74
rect	178	76	179	77
rect	178	82	179	83
rect	178	85	179	86
rect	178	88	179	89
rect	178	91	179	92
rect	178	94	179	95
rect	178	100	179	101
rect	178	103	179	104
rect	178	106	179	107
rect	178	109	179	110
rect	178	112	179	113
rect	178	127	179	128
rect	178	130	179	131
rect	178	136	179	137
rect	178	139	179	140
rect	178	142	179	143
rect	178	151	179	152
rect	178	154	179	155
rect	178	157	179	158
rect	178	160	179	161
rect	178	163	179	164
rect	178	172	179	173
rect	178	175	179	176
rect	178	178	179	179
rect	178	181	179	182
rect	178	184	179	185
rect	178	187	179	188
rect	178	196	179	197
rect	178	205	179	206
rect	178	214	179	215
rect	178	217	179	218
rect	178	220	179	221
rect	178	223	179	224
rect	178	229	179	230
rect	178	232	179	233
rect	178	235	179	236
rect	178	241	179	242
rect	178	244	179	245
rect	178	259	179	260
rect	178	262	179	263
rect	178	265	179	266
rect	178	268	179	269
rect	178	274	179	275
rect	178	277	179	278
rect	178	286	179	287
rect	178	289	179	290
rect	178	292	179	293
rect	178	301	179	302
rect	178	304	179	305
rect	178	313	179	314
rect	178	322	179	323
rect	178	325	179	326
rect	178	328	179	329
rect	179	13	180	14
rect	179	16	180	17
rect	179	19	180	20
rect	179	28	180	29
rect	179	31	180	32
rect	179	37	180	38
rect	179	40	180	41
rect	179	49	180	50
rect	179	52	180	53
rect	179	55	180	56
rect	179	58	180	59
rect	179	61	180	62
rect	179	70	180	71
rect	179	73	180	74
rect	179	76	180	77
rect	179	82	180	83
rect	179	85	180	86
rect	179	88	180	89
rect	179	91	180	92
rect	179	94	180	95
rect	179	100	180	101
rect	179	103	180	104
rect	179	106	180	107
rect	179	109	180	110
rect	179	112	180	113
rect	179	127	180	128
rect	179	130	180	131
rect	179	136	180	137
rect	179	139	180	140
rect	179	142	180	143
rect	179	151	180	152
rect	179	154	180	155
rect	179	157	180	158
rect	179	160	180	161
rect	179	163	180	164
rect	179	172	180	173
rect	179	175	180	176
rect	179	178	180	179
rect	179	184	180	185
rect	179	187	180	188
rect	179	196	180	197
rect	179	205	180	206
rect	179	214	180	215
rect	179	217	180	218
rect	179	220	180	221
rect	179	223	180	224
rect	179	229	180	230
rect	179	232	180	233
rect	179	235	180	236
rect	179	241	180	242
rect	179	244	180	245
rect	179	259	180	260
rect	179	262	180	263
rect	179	265	180	266
rect	179	268	180	269
rect	179	274	180	275
rect	179	277	180	278
rect	179	286	180	287
rect	179	289	180	290
rect	179	292	180	293
rect	179	301	180	302
rect	179	304	180	305
rect	179	313	180	314
rect	179	322	180	323
rect	179	325	180	326
rect	179	328	180	329
rect	180	13	181	14
rect	180	16	181	17
rect	180	19	181	20
rect	180	28	181	29
rect	180	31	181	32
rect	180	37	181	38
rect	180	40	181	41
rect	180	49	181	50
rect	180	52	181	53
rect	180	55	181	56
rect	180	58	181	59
rect	180	61	181	62
rect	180	70	181	71
rect	180	73	181	74
rect	180	76	181	77
rect	180	82	181	83
rect	180	85	181	86
rect	180	88	181	89
rect	180	91	181	92
rect	180	94	181	95
rect	180	100	181	101
rect	180	103	181	104
rect	180	106	181	107
rect	180	109	181	110
rect	180	112	181	113
rect	180	127	181	128
rect	180	130	181	131
rect	180	136	181	137
rect	180	139	181	140
rect	180	142	181	143
rect	180	151	181	152
rect	180	154	181	155
rect	180	157	181	158
rect	180	160	181	161
rect	180	163	181	164
rect	180	172	181	173
rect	180	175	181	176
rect	180	178	181	179
rect	180	184	181	185
rect	180	187	181	188
rect	180	196	181	197
rect	180	199	181	200
rect	180	205	181	206
rect	180	214	181	215
rect	180	217	181	218
rect	180	220	181	221
rect	180	223	181	224
rect	180	229	181	230
rect	180	232	181	233
rect	180	235	181	236
rect	180	241	181	242
rect	180	244	181	245
rect	180	259	181	260
rect	180	262	181	263
rect	180	265	181	266
rect	180	268	181	269
rect	180	274	181	275
rect	180	277	181	278
rect	180	286	181	287
rect	180	289	181	290
rect	180	292	181	293
rect	180	301	181	302
rect	180	304	181	305
rect	180	313	181	314
rect	180	322	181	323
rect	180	325	181	326
rect	180	328	181	329
rect	181	13	182	14
rect	181	16	182	17
rect	181	19	182	20
rect	181	28	182	29
rect	181	31	182	32
rect	181	37	182	38
rect	181	40	182	41
rect	181	49	182	50
rect	181	52	182	53
rect	181	55	182	56
rect	181	58	182	59
rect	181	61	182	62
rect	181	70	182	71
rect	181	73	182	74
rect	181	76	182	77
rect	181	82	182	83
rect	181	88	182	89
rect	181	91	182	92
rect	181	94	182	95
rect	181	103	182	104
rect	181	106	182	107
rect	181	109	182	110
rect	181	112	182	113
rect	181	127	182	128
rect	181	130	182	131
rect	181	136	182	137
rect	181	139	182	140
rect	181	142	182	143
rect	181	151	182	152
rect	181	154	182	155
rect	181	157	182	158
rect	181	163	182	164
rect	181	172	182	173
rect	181	175	182	176
rect	181	178	182	179
rect	181	184	182	185
rect	181	187	182	188
rect	181	196	182	197
rect	181	199	182	200
rect	181	205	182	206
rect	181	214	182	215
rect	181	217	182	218
rect	181	220	182	221
rect	181	223	182	224
rect	181	229	182	230
rect	181	232	182	233
rect	181	235	182	236
rect	181	241	182	242
rect	181	244	182	245
rect	181	259	182	260
rect	181	262	182	263
rect	181	265	182	266
rect	181	268	182	269
rect	181	274	182	275
rect	181	277	182	278
rect	181	286	182	287
rect	181	289	182	290
rect	181	292	182	293
rect	181	301	182	302
rect	181	304	182	305
rect	181	322	182	323
rect	181	325	182	326
rect	181	328	182	329
rect	182	13	183	14
rect	182	16	183	17
rect	182	19	183	20
rect	182	28	183	29
rect	182	31	183	32
rect	182	37	183	38
rect	182	40	183	41
rect	182	49	183	50
rect	182	52	183	53
rect	182	55	183	56
rect	182	58	183	59
rect	182	61	183	62
rect	182	70	183	71
rect	182	73	183	74
rect	182	76	183	77
rect	182	82	183	83
rect	182	88	183	89
rect	182	91	183	92
rect	182	94	183	95
rect	182	103	183	104
rect	182	106	183	107
rect	182	109	183	110
rect	182	112	183	113
rect	182	127	183	128
rect	182	130	183	131
rect	182	136	183	137
rect	182	139	183	140
rect	182	142	183	143
rect	182	151	183	152
rect	182	154	183	155
rect	182	157	183	158
rect	182	163	183	164
rect	182	172	183	173
rect	182	175	183	176
rect	182	178	183	179
rect	182	181	183	182
rect	182	184	183	185
rect	182	187	183	188
rect	182	196	183	197
rect	182	199	183	200
rect	182	205	183	206
rect	182	214	183	215
rect	182	217	183	218
rect	182	220	183	221
rect	182	223	183	224
rect	182	229	183	230
rect	182	232	183	233
rect	182	235	183	236
rect	182	241	183	242
rect	182	244	183	245
rect	182	259	183	260
rect	182	262	183	263
rect	182	265	183	266
rect	182	268	183	269
rect	182	274	183	275
rect	182	277	183	278
rect	182	286	183	287
rect	182	289	183	290
rect	182	292	183	293
rect	182	301	183	302
rect	182	304	183	305
rect	182	319	183	320
rect	182	322	183	323
rect	182	325	183	326
rect	182	328	183	329
rect	183	13	184	14
rect	183	19	184	20
rect	183	28	184	29
rect	183	31	184	32
rect	183	37	184	38
rect	183	40	184	41
rect	183	49	184	50
rect	183	52	184	53
rect	183	55	184	56
rect	183	58	184	59
rect	183	61	184	62
rect	183	70	184	71
rect	183	73	184	74
rect	183	76	184	77
rect	183	82	184	83
rect	183	88	184	89
rect	183	91	184	92
rect	183	94	184	95
rect	183	103	184	104
rect	183	106	184	107
rect	183	109	184	110
rect	183	112	184	113
rect	183	127	184	128
rect	183	130	184	131
rect	183	136	184	137
rect	183	139	184	140
rect	183	142	184	143
rect	183	151	184	152
rect	183	154	184	155
rect	183	157	184	158
rect	183	163	184	164
rect	183	172	184	173
rect	183	175	184	176
rect	183	178	184	179
rect	183	181	184	182
rect	183	184	184	185
rect	183	187	184	188
rect	183	196	184	197
rect	183	199	184	200
rect	183	205	184	206
rect	183	214	184	215
rect	183	217	184	218
rect	183	220	184	221
rect	183	223	184	224
rect	183	229	184	230
rect	183	232	184	233
rect	183	235	184	236
rect	183	241	184	242
rect	183	244	184	245
rect	183	259	184	260
rect	183	262	184	263
rect	183	265	184	266
rect	183	274	184	275
rect	183	277	184	278
rect	183	286	184	287
rect	183	289	184	290
rect	183	292	184	293
rect	183	301	184	302
rect	183	319	184	320
rect	183	322	184	323
rect	183	325	184	326
rect	183	328	184	329
rect	184	13	185	14
rect	184	19	185	20
rect	184	28	185	29
rect	184	31	185	32
rect	184	37	185	38
rect	184	40	185	41
rect	184	49	185	50
rect	184	52	185	53
rect	184	55	185	56
rect	184	58	185	59
rect	184	61	185	62
rect	184	70	185	71
rect	184	73	185	74
rect	184	76	185	77
rect	184	82	185	83
rect	184	88	185	89
rect	184	91	185	92
rect	184	94	185	95
rect	184	103	185	104
rect	184	106	185	107
rect	184	109	185	110
rect	184	112	185	113
rect	184	127	185	128
rect	184	130	185	131
rect	184	136	185	137
rect	184	139	185	140
rect	184	142	185	143
rect	184	151	185	152
rect	184	154	185	155
rect	184	157	185	158
rect	184	163	185	164
rect	184	172	185	173
rect	184	175	185	176
rect	184	178	185	179
rect	184	181	185	182
rect	184	184	185	185
rect	184	187	185	188
rect	184	196	185	197
rect	184	199	185	200
rect	184	205	185	206
rect	184	214	185	215
rect	184	217	185	218
rect	184	220	185	221
rect	184	223	185	224
rect	184	229	185	230
rect	184	232	185	233
rect	184	235	185	236
rect	184	241	185	242
rect	184	244	185	245
rect	184	259	185	260
rect	184	262	185	263
rect	184	265	185	266
rect	184	274	185	275
rect	184	277	185	278
rect	184	286	185	287
rect	184	289	185	290
rect	184	292	185	293
rect	184	301	185	302
rect	184	316	185	317
rect	184	319	185	320
rect	184	322	185	323
rect	184	325	185	326
rect	184	328	185	329
rect	185	13	186	14
rect	185	19	186	20
rect	185	28	186	29
rect	185	31	186	32
rect	185	37	186	38
rect	185	40	186	41
rect	185	49	186	50
rect	185	52	186	53
rect	185	55	186	56
rect	185	58	186	59
rect	185	61	186	62
rect	185	70	186	71
rect	185	73	186	74
rect	185	76	186	77
rect	185	82	186	83
rect	185	88	186	89
rect	185	94	186	95
rect	185	103	186	104
rect	185	109	186	110
rect	185	112	186	113
rect	185	127	186	128
rect	185	130	186	131
rect	185	136	186	137
rect	185	139	186	140
rect	185	142	186	143
rect	185	151	186	152
rect	185	154	186	155
rect	185	163	186	164
rect	185	172	186	173
rect	185	175	186	176
rect	185	178	186	179
rect	185	181	186	182
rect	185	184	186	185
rect	185	187	186	188
rect	185	196	186	197
rect	185	199	186	200
rect	185	205	186	206
rect	185	214	186	215
rect	185	217	186	218
rect	185	220	186	221
rect	185	223	186	224
rect	185	229	186	230
rect	185	232	186	233
rect	185	235	186	236
rect	185	241	186	242
rect	185	244	186	245
rect	185	259	186	260
rect	185	262	186	263
rect	185	265	186	266
rect	185	277	186	278
rect	185	286	186	287
rect	185	289	186	290
rect	185	292	186	293
rect	185	316	186	317
rect	185	319	186	320
rect	185	322	186	323
rect	185	325	186	326
rect	185	328	186	329
rect	186	13	187	14
rect	186	19	187	20
rect	186	28	187	29
rect	186	31	187	32
rect	186	37	187	38
rect	186	40	187	41
rect	186	49	187	50
rect	186	52	187	53
rect	186	55	187	56
rect	186	58	187	59
rect	186	61	187	62
rect	186	70	187	71
rect	186	73	187	74
rect	186	76	187	77
rect	186	82	187	83
rect	186	88	187	89
rect	186	94	187	95
rect	186	100	187	101
rect	186	103	187	104
rect	186	109	187	110
rect	186	112	187	113
rect	186	124	187	125
rect	186	127	187	128
rect	186	130	187	131
rect	186	136	187	137
rect	186	139	187	140
rect	186	142	187	143
rect	186	151	187	152
rect	186	154	187	155
rect	186	160	187	161
rect	186	163	187	164
rect	186	172	187	173
rect	186	175	187	176
rect	186	178	187	179
rect	186	181	187	182
rect	186	184	187	185
rect	186	187	187	188
rect	186	196	187	197
rect	186	199	187	200
rect	186	205	187	206
rect	186	214	187	215
rect	186	217	187	218
rect	186	220	187	221
rect	186	223	187	224
rect	186	229	187	230
rect	186	232	187	233
rect	186	235	187	236
rect	186	241	187	242
rect	186	244	187	245
rect	186	259	187	260
rect	186	262	187	263
rect	186	265	187	266
rect	186	268	187	269
rect	186	277	187	278
rect	186	286	187	287
rect	186	289	187	290
rect	186	292	187	293
rect	186	313	187	314
rect	186	316	187	317
rect	186	319	187	320
rect	186	322	187	323
rect	186	325	187	326
rect	186	328	187	329
rect	187	13	188	14
rect	187	19	188	20
rect	187	28	188	29
rect	187	31	188	32
rect	187	37	188	38
rect	187	40	188	41
rect	187	52	188	53
rect	187	55	188	56
rect	187	58	188	59
rect	187	61	188	62
rect	187	70	188	71
rect	187	73	188	74
rect	187	76	188	77
rect	187	88	188	89
rect	187	94	188	95
rect	187	100	188	101
rect	187	103	188	104
rect	187	109	188	110
rect	187	112	188	113
rect	187	124	188	125
rect	187	127	188	128
rect	187	130	188	131
rect	187	136	188	137
rect	187	139	188	140
rect	187	142	188	143
rect	187	151	188	152
rect	187	154	188	155
rect	187	160	188	161
rect	187	163	188	164
rect	187	172	188	173
rect	187	175	188	176
rect	187	178	188	179
rect	187	181	188	182
rect	187	184	188	185
rect	187	187	188	188
rect	187	196	188	197
rect	187	199	188	200
rect	187	205	188	206
rect	187	214	188	215
rect	187	217	188	218
rect	187	220	188	221
rect	187	223	188	224
rect	187	229	188	230
rect	187	232	188	233
rect	187	235	188	236
rect	187	241	188	242
rect	187	244	188	245
rect	187	259	188	260
rect	187	262	188	263
rect	187	265	188	266
rect	187	268	188	269
rect	187	277	188	278
rect	187	286	188	287
rect	187	289	188	290
rect	187	292	188	293
rect	187	313	188	314
rect	187	316	188	317
rect	187	319	188	320
rect	187	322	188	323
rect	187	325	188	326
rect	187	328	188	329
rect	188	13	189	14
rect	188	19	189	20
rect	188	28	189	29
rect	188	31	189	32
rect	188	37	189	38
rect	188	40	189	41
rect	188	44	189	45
rect	188	52	189	53
rect	188	55	189	56
rect	188	58	189	59
rect	188	61	189	62
rect	188	70	189	71
rect	188	73	189	74
rect	188	76	189	77
rect	188	88	189	89
rect	188	94	189	95
rect	188	100	189	101
rect	188	103	189	104
rect	188	109	189	110
rect	188	112	189	113
rect	188	124	189	125
rect	188	127	189	128
rect	188	130	189	131
rect	188	136	189	137
rect	188	139	189	140
rect	188	142	189	143
rect	188	151	189	152
rect	188	154	189	155
rect	188	160	189	161
rect	188	163	189	164
rect	188	172	189	173
rect	188	175	189	176
rect	188	178	189	179
rect	188	181	189	182
rect	188	184	189	185
rect	188	187	189	188
rect	188	196	189	197
rect	188	199	189	200
rect	188	205	189	206
rect	188	214	189	215
rect	188	217	189	218
rect	188	220	189	221
rect	188	223	189	224
rect	188	229	189	230
rect	188	232	189	233
rect	188	235	189	236
rect	188	241	189	242
rect	188	244	189	245
rect	188	259	189	260
rect	188	262	189	263
rect	188	265	189	266
rect	188	268	189	269
rect	188	277	189	278
rect	188	286	189	287
rect	188	289	189	290
rect	188	292	189	293
rect	188	304	189	305
rect	188	313	189	314
rect	188	316	189	317
rect	188	319	189	320
rect	188	322	189	323
rect	188	325	189	326
rect	188	328	189	329
rect	189	13	190	14
rect	189	19	190	20
rect	189	28	190	29
rect	189	31	190	32
rect	189	40	190	41
rect	189	44	190	45
rect	189	52	190	53
rect	189	55	190	56
rect	189	58	190	59
rect	189	70	190	71
rect	189	73	190	74
rect	189	88	190	89
rect	189	94	190	95
rect	189	100	190	101
rect	189	103	190	104
rect	189	109	190	110
rect	189	124	190	125
rect	189	127	190	128
rect	189	130	190	131
rect	189	136	190	137
rect	189	142	190	143
rect	189	151	190	152
rect	189	154	190	155
rect	189	160	190	161
rect	189	163	190	164
rect	189	172	190	173
rect	189	178	190	179
rect	189	181	190	182
rect	189	184	190	185
rect	189	187	190	188
rect	189	196	190	197
rect	189	199	190	200
rect	189	205	190	206
rect	189	214	190	215
rect	189	217	190	218
rect	189	220	190	221
rect	189	223	190	224
rect	189	229	190	230
rect	189	232	190	233
rect	189	235	190	236
rect	189	241	190	242
rect	189	244	190	245
rect	189	259	190	260
rect	189	262	190	263
rect	189	265	190	266
rect	189	268	190	269
rect	189	286	190	287
rect	189	289	190	290
rect	189	304	190	305
rect	189	313	190	314
rect	189	316	190	317
rect	189	319	190	320
rect	189	322	190	323
rect	189	325	190	326
rect	189	328	190	329
rect	190	13	191	14
rect	190	19	191	20
rect	190	28	191	29
rect	190	31	191	32
rect	190	40	191	41
rect	190	44	191	45
rect	190	46	191	47
rect	190	52	191	53
rect	190	55	191	56
rect	190	58	191	59
rect	190	67	191	68
rect	190	70	191	71
rect	190	73	191	74
rect	190	88	191	89
rect	190	91	191	92
rect	190	94	191	95
rect	190	100	191	101
rect	190	103	191	104
rect	190	106	191	107
rect	190	109	191	110
rect	190	124	191	125
rect	190	127	191	128
rect	190	130	191	131
rect	190	136	191	137
rect	190	142	191	143
rect	190	151	191	152
rect	190	154	191	155
rect	190	157	191	158
rect	190	160	191	161
rect	190	163	191	164
rect	190	172	191	173
rect	190	178	191	179
rect	190	181	191	182
rect	190	184	191	185
rect	190	187	191	188
rect	190	193	191	194
rect	190	196	191	197
rect	190	199	191	200
rect	190	205	191	206
rect	190	211	191	212
rect	190	214	191	215
rect	190	217	191	218
rect	190	220	191	221
rect	190	223	191	224
rect	190	229	191	230
rect	190	232	191	233
rect	190	235	191	236
rect	190	241	191	242
rect	190	244	191	245
rect	190	259	191	260
rect	190	262	191	263
rect	190	265	191	266
rect	190	268	191	269
rect	190	286	191	287
rect	190	289	191	290
rect	190	301	191	302
rect	190	304	191	305
rect	190	313	191	314
rect	190	316	191	317
rect	190	319	191	320
rect	190	322	191	323
rect	190	325	191	326
rect	190	328	191	329
rect	191	13	192	14
rect	191	28	192	29
rect	191	40	192	41
rect	191	44	192	45
rect	191	46	192	47
rect	191	52	192	53
rect	191	55	192	56
rect	191	58	192	59
rect	191	67	192	68
rect	191	70	192	71
rect	191	73	192	74
rect	191	88	192	89
rect	191	91	192	92
rect	191	94	192	95
rect	191	100	192	101
rect	191	103	192	104
rect	191	106	192	107
rect	191	109	192	110
rect	191	124	192	125
rect	191	130	192	131
rect	191	136	192	137
rect	191	142	192	143
rect	191	151	192	152
rect	191	154	192	155
rect	191	157	192	158
rect	191	160	192	161
rect	191	163	192	164
rect	191	172	192	173
rect	191	178	192	179
rect	191	181	192	182
rect	191	184	192	185
rect	191	193	192	194
rect	191	199	192	200
rect	191	205	192	206
rect	191	211	192	212
rect	191	217	192	218
rect	191	220	192	221
rect	191	223	192	224
rect	191	229	192	230
rect	191	232	192	233
rect	191	235	192	236
rect	191	241	192	242
rect	191	244	192	245
rect	191	259	192	260
rect	191	262	192	263
rect	191	268	192	269
rect	191	286	192	287
rect	191	301	192	302
rect	191	304	192	305
rect	191	313	192	314
rect	191	316	192	317
rect	191	319	192	320
rect	191	322	192	323
rect	191	325	192	326
rect	192	13	193	14
rect	192	25	193	26
rect	192	28	193	29
rect	192	40	193	41
rect	192	44	193	45
rect	192	46	193	47
rect	192	52	193	53
rect	192	55	193	56
rect	192	58	193	59
rect	192	67	193	68
rect	192	70	193	71
rect	192	73	193	74
rect	192	88	193	89
rect	192	91	193	92
rect	192	94	193	95
rect	192	100	193	101
rect	192	103	193	104
rect	192	106	193	107
rect	192	109	193	110
rect	192	121	193	122
rect	192	124	193	125
rect	192	130	193	131
rect	192	136	193	137
rect	192	139	193	140
rect	192	142	193	143
rect	192	151	193	152
rect	192	154	193	155
rect	192	157	193	158
rect	192	160	193	161
rect	192	163	193	164
rect	192	166	193	167
rect	192	172	193	173
rect	192	178	193	179
rect	192	181	193	182
rect	192	184	193	185
rect	192	190	193	191
rect	192	193	193	194
rect	192	199	193	200
rect	192	205	193	206
rect	192	211	193	212
rect	192	217	193	218
rect	192	220	193	221
rect	192	223	193	224
rect	192	226	193	227
rect	192	229	193	230
rect	192	232	193	233
rect	192	235	193	236
rect	192	241	193	242
rect	192	244	193	245
rect	192	259	193	260
rect	192	262	193	263
rect	192	268	193	269
rect	192	277	193	278
rect	192	286	193	287
rect	192	298	193	299
rect	192	301	193	302
rect	192	304	193	305
rect	192	313	193	314
rect	192	316	193	317
rect	192	319	193	320
rect	192	322	193	323
rect	192	325	193	326
rect	192	334	193	335
rect	193	13	194	14
rect	193	25	194	26
rect	193	40	194	41
rect	193	44	194	45
rect	193	46	194	47
rect	193	55	194	56
rect	193	67	194	68
rect	193	70	194	71
rect	193	91	194	92
rect	193	94	194	95
rect	193	100	194	101
rect	193	106	194	107
rect	193	109	194	110
rect	193	121	194	122
rect	193	124	194	125
rect	193	130	194	131
rect	193	139	194	140
rect	193	142	194	143
rect	193	151	194	152
rect	193	157	194	158
rect	193	160	194	161
rect	193	163	194	164
rect	193	166	194	167
rect	193	172	194	173
rect	193	181	194	182
rect	193	184	194	185
rect	193	190	194	191
rect	193	193	194	194
rect	193	199	194	200
rect	193	205	194	206
rect	193	211	194	212
rect	193	220	194	221
rect	193	226	194	227
rect	193	232	194	233
rect	193	235	194	236
rect	193	244	194	245
rect	193	262	194	263
rect	193	268	194	269
rect	193	277	194	278
rect	193	298	194	299
rect	193	301	194	302
rect	193	304	194	305
rect	193	313	194	314
rect	193	316	194	317
rect	193	319	194	320
rect	193	322	194	323
rect	193	334	194	335
rect	194	13	195	14
rect	194	16	195	17
rect	194	19	195	20
rect	194	25	195	26
rect	194	37	195	38
rect	194	40	195	41
rect	194	44	195	45
rect	194	46	195	47
rect	194	49	195	50
rect	194	55	195	56
rect	194	64	195	65
rect	194	67	195	68
rect	194	70	195	71
rect	194	79	195	80
rect	194	82	195	83
rect	194	91	195	92
rect	194	94	195	95
rect	194	100	195	101
rect	194	106	195	107
rect	194	109	195	110
rect	194	115	195	116
rect	194	118	195	119
rect	194	121	195	122
rect	194	124	195	125
rect	194	130	195	131
rect	194	139	195	140
rect	194	142	195	143
rect	194	151	195	152
rect	194	157	195	158
rect	194	160	195	161
rect	194	163	195	164
rect	194	166	195	167
rect	194	172	195	173
rect	194	175	195	176
rect	194	181	195	182
rect	194	184	195	185
rect	194	190	195	191
rect	194	193	195	194
rect	194	196	195	197
rect	194	199	195	200
rect	194	205	195	206
rect	194	211	195	212
rect	194	214	195	215
rect	194	220	195	221
rect	194	226	195	227
rect	194	232	195	233
rect	194	235	195	236
rect	194	238	195	239
rect	194	244	195	245
rect	194	262	195	263
rect	194	268	195	269
rect	194	271	195	272
rect	194	277	195	278
rect	194	295	195	296
rect	194	298	195	299
rect	194	301	195	302
rect	194	304	195	305
rect	194	313	195	314
rect	194	316	195	317
rect	194	319	195	320
rect	194	322	195	323
rect	194	331	195	332
rect	194	334	195	335
rect	195	16	196	17
rect	195	19	196	20
rect	195	25	196	26
rect	195	37	196	38
rect	195	46	196	47
rect	195	49	196	50
rect	195	64	196	65
rect	195	67	196	68
rect	195	79	196	80
rect	195	82	196	83
rect	195	91	196	92
rect	195	100	196	101
rect	195	106	196	107
rect	195	115	196	116
rect	195	118	196	119
rect	195	121	196	122
rect	195	124	196	125
rect	195	139	196	140
rect	195	142	196	143
rect	195	157	196	158
rect	195	160	196	161
rect	195	163	196	164
rect	195	166	196	167
rect	195	175	196	176
rect	195	181	196	182
rect	195	190	196	191
rect	195	193	196	194
rect	195	196	196	197
rect	195	199	196	200
rect	195	211	196	212
rect	195	214	196	215
rect	195	220	196	221
rect	195	226	196	227
rect	195	238	196	239
rect	195	244	196	245
rect	195	268	196	269
rect	195	271	196	272
rect	195	277	196	278
rect	195	295	196	296
rect	195	298	196	299
rect	195	301	196	302
rect	195	304	196	305
rect	195	313	196	314
rect	195	316	196	317
rect	195	319	196	320
rect	195	331	196	332
rect	195	334	196	335
rect	196	16	197	17
rect	196	19	197	20
rect	196	22	197	23
rect	196	25	197	26
rect	196	28	197	29
rect	196	37	197	38
rect	196	46	197	47
rect	196	49	197	50
rect	196	52	197	53
rect	196	61	197	62
rect	196	64	197	65
rect	196	67	197	68
rect	196	76	197	77
rect	196	79	197	80
rect	196	82	197	83
rect	196	88	197	89
rect	196	91	197	92
rect	196	100	197	101
rect	196	103	197	104
rect	196	106	197	107
rect	196	115	197	116
rect	196	118	197	119
rect	196	121	197	122
rect	196	124	197	125
rect	196	127	197	128
rect	196	133	197	134
rect	196	136	197	137
rect	196	139	197	140
rect	196	142	197	143
rect	196	145	197	146
rect	196	154	197	155
rect	196	157	197	158
rect	196	160	197	161
rect	196	163	197	164
rect	196	166	197	167
rect	196	175	197	176
rect	196	178	197	179
rect	196	181	197	182
rect	196	190	197	191
rect	196	193	197	194
rect	196	196	197	197
rect	196	199	197	200
rect	196	211	197	212
rect	196	214	197	215
rect	196	217	197	218
rect	196	220	197	221
rect	196	226	197	227
rect	196	229	197	230
rect	196	238	197	239
rect	196	241	197	242
rect	196	244	197	245
rect	196	253	197	254
rect	196	259	197	260
rect	196	268	197	269
rect	196	271	197	272
rect	196	274	197	275
rect	196	277	197	278
rect	196	286	197	287
rect	196	292	197	293
rect	196	295	197	296
rect	196	298	197	299
rect	196	301	197	302
rect	196	304	197	305
rect	196	313	197	314
rect	196	316	197	317
rect	196	319	197	320
rect	196	328	197	329
rect	196	331	197	332
rect	196	334	197	335
rect	203	10	204	11
rect	203	19	204	20
rect	203	22	204	23
rect	203	25	204	26
rect	203	28	204	29
rect	203	37	204	38
rect	203	46	204	47
rect	203	49	204	50
rect	203	52	204	53
rect	203	61	204	62
rect	203	64	204	65
rect	203	67	204	68
rect	203	70	204	71
rect	203	76	204	77
rect	203	79	204	80
rect	203	88	204	89
rect	203	91	204	92
rect	203	100	204	101
rect	203	103	204	104
rect	203	106	204	107
rect	203	115	204	116
rect	203	118	204	119
rect	203	121	204	122
rect	203	124	204	125
rect	203	127	204	128
rect	203	136	204	137
rect	203	139	204	140
rect	203	142	204	143
rect	203	145	204	146
rect	203	154	204	155
rect	203	157	204	158
rect	203	160	204	161
rect	203	163	204	164
rect	203	166	204	167
rect	203	175	204	176
rect	203	178	204	179
rect	203	181	204	182
rect	203	190	204	191
rect	203	193	204	194
rect	203	196	204	197
rect	203	199	204	200
rect	203	214	204	215
rect	203	217	204	218
rect	203	220	204	221
rect	203	229	204	230
rect	203	232	204	233
rect	203	238	204	239
rect	203	241	204	242
rect	203	244	204	245
rect	203	253	204	254
rect	203	256	204	257
rect	203	259	204	260
rect	203	262	204	263
rect	203	265	204	266
rect	203	268	204	269
rect	203	271	204	272
rect	203	274	204	275
rect	203	277	204	278
rect	203	286	204	287
rect	203	295	204	296
rect	203	298	204	299
rect	203	301	204	302
rect	203	304	204	305
rect	203	313	204	314
rect	203	316	204	317
rect	203	319	204	320
rect	203	328	204	329
rect	203	331	204	332
rect	203	334	204	335
rect	204	10	205	11
rect	204	19	205	20
rect	204	22	205	23
rect	204	25	205	26
rect	204	28	205	29
rect	204	37	205	38
rect	204	46	205	47
rect	204	49	205	50
rect	204	52	205	53
rect	204	61	205	62
rect	204	64	205	65
rect	204	67	205	68
rect	204	70	205	71
rect	204	76	205	77
rect	204	79	205	80
rect	204	88	205	89
rect	204	91	205	92
rect	204	100	205	101
rect	204	103	205	104
rect	204	106	205	107
rect	204	115	205	116
rect	204	118	205	119
rect	204	121	205	122
rect	204	124	205	125
rect	204	127	205	128
rect	204	136	205	137
rect	204	139	205	140
rect	204	145	205	146
rect	204	154	205	155
rect	204	157	205	158
rect	204	160	205	161
rect	204	163	205	164
rect	204	166	205	167
rect	204	175	205	176
rect	204	178	205	179
rect	204	181	205	182
rect	204	190	205	191
rect	204	193	205	194
rect	204	196	205	197
rect	204	199	205	200
rect	204	214	205	215
rect	204	217	205	218
rect	204	220	205	221
rect	204	229	205	230
rect	204	232	205	233
rect	204	238	205	239
rect	204	241	205	242
rect	204	244	205	245
rect	204	253	205	254
rect	204	256	205	257
rect	204	259	205	260
rect	204	262	205	263
rect	204	265	205	266
rect	204	268	205	269
rect	204	271	205	272
rect	204	274	205	275
rect	204	277	205	278
rect	204	286	205	287
rect	204	295	205	296
rect	204	298	205	299
rect	204	301	205	302
rect	204	304	205	305
rect	204	313	205	314
rect	204	316	205	317
rect	204	319	205	320
rect	204	328	205	329
rect	204	331	205	332
rect	204	334	205	335
rect	205	10	206	11
rect	205	19	206	20
rect	205	22	206	23
rect	205	25	206	26
rect	205	28	206	29
rect	205	37	206	38
rect	205	46	206	47
rect	205	49	206	50
rect	205	52	206	53
rect	205	61	206	62
rect	205	64	206	65
rect	205	67	206	68
rect	205	70	206	71
rect	205	76	206	77
rect	205	79	206	80
rect	205	88	206	89
rect	205	91	206	92
rect	205	100	206	101
rect	205	103	206	104
rect	205	106	206	107
rect	205	115	206	116
rect	205	118	206	119
rect	205	121	206	122
rect	205	124	206	125
rect	205	127	206	128
rect	205	136	206	137
rect	205	139	206	140
rect	205	145	206	146
rect	205	151	206	152
rect	205	154	206	155
rect	205	157	206	158
rect	205	160	206	161
rect	205	163	206	164
rect	205	166	206	167
rect	205	175	206	176
rect	205	178	206	179
rect	205	181	206	182
rect	205	190	206	191
rect	205	193	206	194
rect	205	196	206	197
rect	205	199	206	200
rect	205	214	206	215
rect	205	217	206	218
rect	205	220	206	221
rect	205	229	206	230
rect	205	232	206	233
rect	205	238	206	239
rect	205	241	206	242
rect	205	244	206	245
rect	205	253	206	254
rect	205	256	206	257
rect	205	259	206	260
rect	205	262	206	263
rect	205	265	206	266
rect	205	268	206	269
rect	205	271	206	272
rect	205	274	206	275
rect	205	277	206	278
rect	205	286	206	287
rect	205	295	206	296
rect	205	298	206	299
rect	205	301	206	302
rect	205	304	206	305
rect	205	313	206	314
rect	205	316	206	317
rect	205	319	206	320
rect	205	328	206	329
rect	205	331	206	332
rect	205	334	206	335
rect	206	10	207	11
rect	206	19	207	20
rect	206	22	207	23
rect	206	25	207	26
rect	206	28	207	29
rect	206	37	207	38
rect	206	46	207	47
rect	206	49	207	50
rect	206	52	207	53
rect	206	61	207	62
rect	206	64	207	65
rect	206	67	207	68
rect	206	70	207	71
rect	206	76	207	77
rect	206	79	207	80
rect	206	88	207	89
rect	206	91	207	92
rect	206	100	207	101
rect	206	103	207	104
rect	206	106	207	107
rect	206	115	207	116
rect	206	118	207	119
rect	206	121	207	122
rect	206	124	207	125
rect	206	136	207	137
rect	206	139	207	140
rect	206	145	207	146
rect	206	151	207	152
rect	206	154	207	155
rect	206	157	207	158
rect	206	160	207	161
rect	206	163	207	164
rect	206	166	207	167
rect	206	175	207	176
rect	206	178	207	179
rect	206	181	207	182
rect	206	190	207	191
rect	206	193	207	194
rect	206	196	207	197
rect	206	199	207	200
rect	206	214	207	215
rect	206	217	207	218
rect	206	220	207	221
rect	206	229	207	230
rect	206	232	207	233
rect	206	238	207	239
rect	206	241	207	242
rect	206	244	207	245
rect	206	253	207	254
rect	206	256	207	257
rect	206	259	207	260
rect	206	262	207	263
rect	206	265	207	266
rect	206	268	207	269
rect	206	271	207	272
rect	206	274	207	275
rect	206	277	207	278
rect	206	286	207	287
rect	206	295	207	296
rect	206	298	207	299
rect	206	301	207	302
rect	206	304	207	305
rect	206	313	207	314
rect	206	316	207	317
rect	206	319	207	320
rect	206	328	207	329
rect	206	331	207	332
rect	206	334	207	335
rect	207	10	208	11
rect	207	19	208	20
rect	207	22	208	23
rect	207	25	208	26
rect	207	28	208	29
rect	207	37	208	38
rect	207	46	208	47
rect	207	49	208	50
rect	207	52	208	53
rect	207	61	208	62
rect	207	64	208	65
rect	207	67	208	68
rect	207	70	208	71
rect	207	76	208	77
rect	207	79	208	80
rect	207	88	208	89
rect	207	91	208	92
rect	207	100	208	101
rect	207	103	208	104
rect	207	106	208	107
rect	207	115	208	116
rect	207	118	208	119
rect	207	121	208	122
rect	207	124	208	125
rect	207	136	208	137
rect	207	139	208	140
rect	207	142	208	143
rect	207	145	208	146
rect	207	151	208	152
rect	207	154	208	155
rect	207	157	208	158
rect	207	160	208	161
rect	207	163	208	164
rect	207	166	208	167
rect	207	175	208	176
rect	207	178	208	179
rect	207	181	208	182
rect	207	190	208	191
rect	207	193	208	194
rect	207	196	208	197
rect	207	199	208	200
rect	207	214	208	215
rect	207	217	208	218
rect	207	220	208	221
rect	207	229	208	230
rect	207	232	208	233
rect	207	238	208	239
rect	207	241	208	242
rect	207	244	208	245
rect	207	253	208	254
rect	207	256	208	257
rect	207	259	208	260
rect	207	262	208	263
rect	207	265	208	266
rect	207	268	208	269
rect	207	271	208	272
rect	207	274	208	275
rect	207	277	208	278
rect	207	286	208	287
rect	207	295	208	296
rect	207	298	208	299
rect	207	301	208	302
rect	207	304	208	305
rect	207	313	208	314
rect	207	316	208	317
rect	207	319	208	320
rect	207	328	208	329
rect	207	331	208	332
rect	207	334	208	335
rect	208	10	209	11
rect	208	19	209	20
rect	208	22	209	23
rect	208	25	209	26
rect	208	28	209	29
rect	208	37	209	38
rect	208	46	209	47
rect	208	49	209	50
rect	208	52	209	53
rect	208	61	209	62
rect	208	64	209	65
rect	208	67	209	68
rect	208	70	209	71
rect	208	76	209	77
rect	208	79	209	80
rect	208	88	209	89
rect	208	91	209	92
rect	208	103	209	104
rect	208	106	209	107
rect	208	115	209	116
rect	208	118	209	119
rect	208	121	209	122
rect	208	136	209	137
rect	208	139	209	140
rect	208	142	209	143
rect	208	145	209	146
rect	208	151	209	152
rect	208	154	209	155
rect	208	157	209	158
rect	208	160	209	161
rect	208	163	209	164
rect	208	166	209	167
rect	208	175	209	176
rect	208	178	209	179
rect	208	181	209	182
rect	208	190	209	191
rect	208	193	209	194
rect	208	196	209	197
rect	208	214	209	215
rect	208	217	209	218
rect	208	220	209	221
rect	208	229	209	230
rect	208	232	209	233
rect	208	238	209	239
rect	208	241	209	242
rect	208	244	209	245
rect	208	253	209	254
rect	208	256	209	257
rect	208	259	209	260
rect	208	262	209	263
rect	208	265	209	266
rect	208	268	209	269
rect	208	271	209	272
rect	208	274	209	275
rect	208	277	209	278
rect	208	286	209	287
rect	208	295	209	296
rect	208	298	209	299
rect	208	301	209	302
rect	208	304	209	305
rect	208	313	209	314
rect	208	316	209	317
rect	208	319	209	320
rect	208	328	209	329
rect	208	331	209	332
rect	208	334	209	335
rect	209	10	210	11
rect	209	19	210	20
rect	209	22	210	23
rect	209	25	210	26
rect	209	28	210	29
rect	209	37	210	38
rect	209	46	210	47
rect	209	49	210	50
rect	209	52	210	53
rect	209	61	210	62
rect	209	64	210	65
rect	209	67	210	68
rect	209	70	210	71
rect	209	76	210	77
rect	209	79	210	80
rect	209	88	210	89
rect	209	91	210	92
rect	209	94	210	95
rect	209	103	210	104
rect	209	106	210	107
rect	209	115	210	116
rect	209	118	210	119
rect	209	121	210	122
rect	209	127	210	128
rect	209	136	210	137
rect	209	139	210	140
rect	209	142	210	143
rect	209	145	210	146
rect	209	151	210	152
rect	209	154	210	155
rect	209	157	210	158
rect	209	160	210	161
rect	209	163	210	164
rect	209	166	210	167
rect	209	175	210	176
rect	209	178	210	179
rect	209	181	210	182
rect	209	190	210	191
rect	209	193	210	194
rect	209	196	210	197
rect	209	205	210	206
rect	209	214	210	215
rect	209	217	210	218
rect	209	220	210	221
rect	209	229	210	230
rect	209	232	210	233
rect	209	238	210	239
rect	209	241	210	242
rect	209	244	210	245
rect	209	253	210	254
rect	209	256	210	257
rect	209	259	210	260
rect	209	262	210	263
rect	209	265	210	266
rect	209	268	210	269
rect	209	271	210	272
rect	209	274	210	275
rect	209	277	210	278
rect	209	286	210	287
rect	209	295	210	296
rect	209	298	210	299
rect	209	301	210	302
rect	209	304	210	305
rect	209	313	210	314
rect	209	316	210	317
rect	209	319	210	320
rect	209	328	210	329
rect	209	331	210	332
rect	209	334	210	335
rect	210	10	211	11
rect	210	19	211	20
rect	210	22	211	23
rect	210	25	211	26
rect	210	28	211	29
rect	210	37	211	38
rect	210	46	211	47
rect	210	49	211	50
rect	210	52	211	53
rect	210	61	211	62
rect	210	64	211	65
rect	210	67	211	68
rect	210	70	211	71
rect	210	76	211	77
rect	210	79	211	80
rect	210	88	211	89
rect	210	94	211	95
rect	210	103	211	104
rect	210	106	211	107
rect	210	115	211	116
rect	210	118	211	119
rect	210	127	211	128
rect	210	136	211	137
rect	210	139	211	140
rect	210	142	211	143
rect	210	145	211	146
rect	210	151	211	152
rect	210	154	211	155
rect	210	157	211	158
rect	210	160	211	161
rect	210	163	211	164
rect	210	166	211	167
rect	210	175	211	176
rect	210	178	211	179
rect	210	190	211	191
rect	210	193	211	194
rect	210	205	211	206
rect	210	214	211	215
rect	210	217	211	218
rect	210	220	211	221
rect	210	229	211	230
rect	210	232	211	233
rect	210	238	211	239
rect	210	241	211	242
rect	210	244	211	245
rect	210	253	211	254
rect	210	256	211	257
rect	210	259	211	260
rect	210	262	211	263
rect	210	265	211	266
rect	210	268	211	269
rect	210	271	211	272
rect	210	274	211	275
rect	210	277	211	278
rect	210	286	211	287
rect	210	295	211	296
rect	210	298	211	299
rect	210	301	211	302
rect	210	304	211	305
rect	210	313	211	314
rect	210	316	211	317
rect	210	319	211	320
rect	210	328	211	329
rect	210	331	211	332
rect	210	334	211	335
rect	211	10	212	11
rect	211	19	212	20
rect	211	22	212	23
rect	211	25	212	26
rect	211	28	212	29
rect	211	37	212	38
rect	211	46	212	47
rect	211	49	212	50
rect	211	52	212	53
rect	211	61	212	62
rect	211	64	212	65
rect	211	67	212	68
rect	211	70	212	71
rect	211	76	212	77
rect	211	79	212	80
rect	211	88	212	89
rect	211	94	212	95
rect	211	100	212	101
rect	211	103	212	104
rect	211	106	212	107
rect	211	115	212	116
rect	211	118	212	119
rect	211	124	212	125
rect	211	127	212	128
rect	211	136	212	137
rect	211	139	212	140
rect	211	142	212	143
rect	211	145	212	146
rect	211	151	212	152
rect	211	154	212	155
rect	211	157	212	158
rect	211	160	212	161
rect	211	163	212	164
rect	211	166	212	167
rect	211	175	212	176
rect	211	178	212	179
rect	211	187	212	188
rect	211	190	212	191
rect	211	193	212	194
rect	211	202	212	203
rect	211	205	212	206
rect	211	214	212	215
rect	211	217	212	218
rect	211	220	212	221
rect	211	229	212	230
rect	211	232	212	233
rect	211	238	212	239
rect	211	241	212	242
rect	211	244	212	245
rect	211	253	212	254
rect	211	256	212	257
rect	211	259	212	260
rect	211	262	212	263
rect	211	265	212	266
rect	211	268	212	269
rect	211	271	212	272
rect	211	274	212	275
rect	211	277	212	278
rect	211	286	212	287
rect	211	295	212	296
rect	211	298	212	299
rect	211	301	212	302
rect	211	304	212	305
rect	211	313	212	314
rect	211	316	212	317
rect	211	319	212	320
rect	211	328	212	329
rect	211	331	212	332
rect	211	334	212	335
rect	212	10	213	11
rect	212	19	213	20
rect	212	22	213	23
rect	212	25	213	26
rect	212	28	213	29
rect	212	37	213	38
rect	212	46	213	47
rect	212	49	213	50
rect	212	52	213	53
rect	212	64	213	65
rect	212	67	213	68
rect	212	70	213	71
rect	212	76	213	77
rect	212	79	213	80
rect	212	88	213	89
rect	212	94	213	95
rect	212	100	213	101
rect	212	103	213	104
rect	212	106	213	107
rect	212	115	213	116
rect	212	118	213	119
rect	212	124	213	125
rect	212	127	213	128
rect	212	136	213	137
rect	212	139	213	140
rect	212	142	213	143
rect	212	145	213	146
rect	212	151	213	152
rect	212	154	213	155
rect	212	157	213	158
rect	212	160	213	161
rect	212	163	213	164
rect	212	166	213	167
rect	212	175	213	176
rect	212	178	213	179
rect	212	187	213	188
rect	212	190	213	191
rect	212	193	213	194
rect	212	202	213	203
rect	212	205	213	206
rect	212	214	213	215
rect	212	217	213	218
rect	212	220	213	221
rect	212	229	213	230
rect	212	232	213	233
rect	212	238	213	239
rect	212	241	213	242
rect	212	244	213	245
rect	212	253	213	254
rect	212	259	213	260
rect	212	262	213	263
rect	212	265	213	266
rect	212	268	213	269
rect	212	271	213	272
rect	212	274	213	275
rect	212	277	213	278
rect	212	286	213	287
rect	212	295	213	296
rect	212	298	213	299
rect	212	301	213	302
rect	212	304	213	305
rect	212	313	213	314
rect	212	316	213	317
rect	212	319	213	320
rect	212	328	213	329
rect	212	331	213	332
rect	212	334	213	335
rect	213	10	214	11
rect	213	19	214	20
rect	213	22	214	23
rect	213	25	214	26
rect	213	28	214	29
rect	213	37	214	38
rect	213	46	214	47
rect	213	49	214	50
rect	213	52	214	53
rect	213	64	214	65
rect	213	67	214	68
rect	213	70	214	71
rect	213	76	214	77
rect	213	79	214	80
rect	213	88	214	89
rect	213	94	214	95
rect	213	100	214	101
rect	213	103	214	104
rect	213	106	214	107
rect	213	115	214	116
rect	213	118	214	119
rect	213	124	214	125
rect	213	127	214	128
rect	213	136	214	137
rect	213	139	214	140
rect	213	142	214	143
rect	213	145	214	146
rect	213	151	214	152
rect	213	154	214	155
rect	213	157	214	158
rect	213	160	214	161
rect	213	163	214	164
rect	213	166	214	167
rect	213	175	214	176
rect	213	178	214	179
rect	213	187	214	188
rect	213	190	214	191
rect	213	193	214	194
rect	213	202	214	203
rect	213	205	214	206
rect	213	214	214	215
rect	213	217	214	218
rect	213	220	214	221
rect	213	229	214	230
rect	213	232	214	233
rect	213	238	214	239
rect	213	241	214	242
rect	213	244	214	245
rect	213	253	214	254
rect	213	259	214	260
rect	213	262	214	263
rect	213	265	214	266
rect	213	268	214	269
rect	213	271	214	272
rect	213	274	214	275
rect	213	277	214	278
rect	213	286	214	287
rect	213	295	214	296
rect	213	298	214	299
rect	213	301	214	302
rect	213	304	214	305
rect	213	313	214	314
rect	213	316	214	317
rect	213	319	214	320
rect	213	328	214	329
rect	213	331	214	332
rect	213	334	214	335
rect	214	10	215	11
rect	214	19	215	20
rect	214	22	215	23
rect	214	25	215	26
rect	214	28	215	29
rect	214	37	215	38
rect	214	46	215	47
rect	214	49	215	50
rect	214	52	215	53
rect	214	64	215	65
rect	214	67	215	68
rect	214	70	215	71
rect	214	76	215	77
rect	214	79	215	80
rect	214	88	215	89
rect	214	94	215	95
rect	214	100	215	101
rect	214	103	215	104
rect	214	106	215	107
rect	214	115	215	116
rect	214	118	215	119
rect	214	124	215	125
rect	214	127	215	128
rect	214	136	215	137
rect	214	139	215	140
rect	214	142	215	143
rect	214	145	215	146
rect	214	151	215	152
rect	214	154	215	155
rect	214	157	215	158
rect	214	160	215	161
rect	214	163	215	164
rect	214	166	215	167
rect	214	175	215	176
rect	214	178	215	179
rect	214	187	215	188
rect	214	190	215	191
rect	214	193	215	194
rect	214	202	215	203
rect	214	205	215	206
rect	214	214	215	215
rect	214	217	215	218
rect	214	220	215	221
rect	214	232	215	233
rect	214	238	215	239
rect	214	241	215	242
rect	214	244	215	245
rect	214	253	215	254
rect	214	259	215	260
rect	214	262	215	263
rect	214	265	215	266
rect	214	268	215	269
rect	214	271	215	272
rect	214	274	215	275
rect	214	277	215	278
rect	214	286	215	287
rect	214	295	215	296
rect	214	298	215	299
rect	214	301	215	302
rect	214	304	215	305
rect	214	313	215	314
rect	214	316	215	317
rect	214	319	215	320
rect	214	328	215	329
rect	214	331	215	332
rect	214	334	215	335
rect	215	10	216	11
rect	215	19	216	20
rect	215	22	216	23
rect	215	25	216	26
rect	215	28	216	29
rect	215	37	216	38
rect	215	46	216	47
rect	215	49	216	50
rect	215	52	216	53
rect	215	61	216	62
rect	215	64	216	65
rect	215	67	216	68
rect	215	70	216	71
rect	215	76	216	77
rect	215	79	216	80
rect	215	88	216	89
rect	215	94	216	95
rect	215	100	216	101
rect	215	103	216	104
rect	215	106	216	107
rect	215	115	216	116
rect	215	118	216	119
rect	215	124	216	125
rect	215	127	216	128
rect	215	136	216	137
rect	215	139	216	140
rect	215	142	216	143
rect	215	145	216	146
rect	215	151	216	152
rect	215	154	216	155
rect	215	157	216	158
rect	215	160	216	161
rect	215	163	216	164
rect	215	166	216	167
rect	215	175	216	176
rect	215	178	216	179
rect	215	187	216	188
rect	215	190	216	191
rect	215	193	216	194
rect	215	202	216	203
rect	215	205	216	206
rect	215	214	216	215
rect	215	217	216	218
rect	215	220	216	221
rect	215	232	216	233
rect	215	238	216	239
rect	215	241	216	242
rect	215	244	216	245
rect	215	253	216	254
rect	215	259	216	260
rect	215	262	216	263
rect	215	265	216	266
rect	215	268	216	269
rect	215	271	216	272
rect	215	274	216	275
rect	215	277	216	278
rect	215	286	216	287
rect	215	295	216	296
rect	215	298	216	299
rect	215	301	216	302
rect	215	304	216	305
rect	215	313	216	314
rect	215	316	216	317
rect	215	319	216	320
rect	215	328	216	329
rect	215	331	216	332
rect	215	334	216	335
rect	216	10	217	11
rect	216	19	217	20
rect	216	25	217	26
rect	216	28	217	29
rect	216	37	217	38
rect	216	46	217	47
rect	216	49	217	50
rect	216	52	217	53
rect	216	61	217	62
rect	216	64	217	65
rect	216	67	217	68
rect	216	70	217	71
rect	216	76	217	77
rect	216	79	217	80
rect	216	88	217	89
rect	216	94	217	95
rect	216	100	217	101
rect	216	103	217	104
rect	216	106	217	107
rect	216	115	217	116
rect	216	118	217	119
rect	216	124	217	125
rect	216	127	217	128
rect	216	136	217	137
rect	216	139	217	140
rect	216	142	217	143
rect	216	145	217	146
rect	216	151	217	152
rect	216	154	217	155
rect	216	157	217	158
rect	216	160	217	161
rect	216	163	217	164
rect	216	166	217	167
rect	216	175	217	176
rect	216	178	217	179
rect	216	187	217	188
rect	216	190	217	191
rect	216	193	217	194
rect	216	202	217	203
rect	216	205	217	206
rect	216	214	217	215
rect	216	217	217	218
rect	216	220	217	221
rect	216	232	217	233
rect	216	238	217	239
rect	216	241	217	242
rect	216	244	217	245
rect	216	253	217	254
rect	216	259	217	260
rect	216	262	217	263
rect	216	268	217	269
rect	216	271	217	272
rect	216	274	217	275
rect	216	277	217	278
rect	216	286	217	287
rect	216	295	217	296
rect	216	298	217	299
rect	216	301	217	302
rect	216	304	217	305
rect	216	313	217	314
rect	216	316	217	317
rect	216	319	217	320
rect	216	328	217	329
rect	216	331	217	332
rect	216	334	217	335
rect	217	10	218	11
rect	217	19	218	20
rect	217	25	218	26
rect	217	28	218	29
rect	217	37	218	38
rect	217	46	218	47
rect	217	49	218	50
rect	217	52	218	53
rect	217	61	218	62
rect	217	64	218	65
rect	217	67	218	68
rect	217	70	218	71
rect	217	76	218	77
rect	217	79	218	80
rect	217	88	218	89
rect	217	94	218	95
rect	217	100	218	101
rect	217	103	218	104
rect	217	106	218	107
rect	217	115	218	116
rect	217	118	218	119
rect	217	124	218	125
rect	217	127	218	128
rect	217	136	218	137
rect	217	139	218	140
rect	217	142	218	143
rect	217	145	218	146
rect	217	151	218	152
rect	217	154	218	155
rect	217	157	218	158
rect	217	160	218	161
rect	217	163	218	164
rect	217	166	218	167
rect	217	175	218	176
rect	217	178	218	179
rect	217	187	218	188
rect	217	190	218	191
rect	217	193	218	194
rect	217	202	218	203
rect	217	205	218	206
rect	217	214	218	215
rect	217	217	218	218
rect	217	220	218	221
rect	217	232	218	233
rect	217	238	218	239
rect	217	241	218	242
rect	217	244	218	245
rect	217	253	218	254
rect	217	259	218	260
rect	217	262	218	263
rect	217	268	218	269
rect	217	271	218	272
rect	217	274	218	275
rect	217	277	218	278
rect	217	286	218	287
rect	217	295	218	296
rect	217	298	218	299
rect	217	301	218	302
rect	217	304	218	305
rect	217	313	218	314
rect	217	316	218	317
rect	217	319	218	320
rect	217	328	218	329
rect	217	331	218	332
rect	217	334	218	335
rect	218	10	219	11
rect	218	25	219	26
rect	218	28	219	29
rect	218	46	219	47
rect	218	49	219	50
rect	218	52	219	53
rect	218	61	219	62
rect	218	64	219	65
rect	218	67	219	68
rect	218	70	219	71
rect	218	76	219	77
rect	218	88	219	89
rect	218	94	219	95
rect	218	100	219	101
rect	218	115	219	116
rect	218	118	219	119
rect	218	124	219	125
rect	218	127	219	128
rect	218	136	219	137
rect	218	139	219	140
rect	218	142	219	143
rect	218	145	219	146
rect	218	151	219	152
rect	218	160	219	161
rect	218	163	219	164
rect	218	166	219	167
rect	218	175	219	176
rect	218	178	219	179
rect	218	187	219	188
rect	218	193	219	194
rect	218	202	219	203
rect	218	205	219	206
rect	218	220	219	221
rect	218	232	219	233
rect	218	238	219	239
rect	218	241	219	242
rect	218	253	219	254
rect	218	259	219	260
rect	218	262	219	263
rect	218	268	219	269
rect	218	271	219	272
rect	218	277	219	278
rect	218	286	219	287
rect	218	295	219	296
rect	218	298	219	299
rect	218	301	219	302
rect	218	304	219	305
rect	218	313	219	314
rect	218	316	219	317
rect	218	319	219	320
rect	218	328	219	329
rect	218	331	219	332
rect	218	334	219	335
rect	219	10	220	11
rect	219	25	220	26
rect	219	28	220	29
rect	219	31	220	32
rect	219	40	220	41
rect	219	46	220	47
rect	219	49	220	50
rect	219	52	220	53
rect	219	61	220	62
rect	219	64	220	65
rect	219	67	220	68
rect	219	70	220	71
rect	219	76	220	77
rect	219	82	220	83
rect	219	88	220	89
rect	219	91	220	92
rect	219	94	220	95
rect	219	100	220	101
rect	219	112	220	113
rect	219	115	220	116
rect	219	118	220	119
rect	219	121	220	122
rect	219	124	220	125
rect	219	127	220	128
rect	219	136	220	137
rect	219	139	220	140
rect	219	142	220	143
rect	219	145	220	146
rect	219	151	220	152
rect	219	160	220	161
rect	219	163	220	164
rect	219	166	220	167
rect	219	169	220	170
rect	219	175	220	176
rect	219	178	220	179
rect	219	181	220	182
rect	219	187	220	188
rect	219	193	220	194
rect	219	196	220	197
rect	219	202	220	203
rect	219	205	220	206
rect	219	220	220	221
rect	219	229	220	230
rect	219	232	220	233
rect	219	238	220	239
rect	219	241	220	242
rect	219	250	220	251
rect	219	253	220	254
rect	219	259	220	260
rect	219	262	220	263
rect	219	268	220	269
rect	219	271	220	272
rect	219	277	220	278
rect	219	280	220	281
rect	219	286	220	287
rect	219	295	220	296
rect	219	298	220	299
rect	219	301	220	302
rect	219	304	220	305
rect	219	313	220	314
rect	219	316	220	317
rect	219	319	220	320
rect	219	328	220	329
rect	219	331	220	332
rect	219	334	220	335
rect	220	10	221	11
rect	220	25	221	26
rect	220	31	221	32
rect	220	40	221	41
rect	220	46	221	47
rect	220	52	221	53
rect	220	61	221	62
rect	220	64	221	65
rect	220	70	221	71
rect	220	76	221	77
rect	220	82	221	83
rect	220	88	221	89
rect	220	91	221	92
rect	220	94	221	95
rect	220	100	221	101
rect	220	112	221	113
rect	220	115	221	116
rect	220	121	221	122
rect	220	124	221	125
rect	220	127	221	128
rect	220	136	221	137
rect	220	142	221	143
rect	220	145	221	146
rect	220	151	221	152
rect	220	166	221	167
rect	220	169	221	170
rect	220	175	221	176
rect	220	181	221	182
rect	220	187	221	188
rect	220	196	221	197
rect	220	202	221	203
rect	220	205	221	206
rect	220	220	221	221
rect	220	229	221	230
rect	220	232	221	233
rect	220	238	221	239
rect	220	250	221	251
rect	220	253	221	254
rect	220	259	221	260
rect	220	262	221	263
rect	220	271	221	272
rect	220	280	221	281
rect	220	286	221	287
rect	220	298	221	299
rect	220	301	221	302
rect	220	304	221	305
rect	220	313	221	314
rect	220	316	221	317
rect	220	319	221	320
rect	220	328	221	329
rect	220	331	221	332
rect	220	334	221	335
rect	221	10	222	11
rect	221	19	222	20
rect	221	25	222	26
rect	221	31	222	32
rect	221	34	222	35
rect	221	40	222	41
rect	221	46	222	47
rect	221	52	222	53
rect	221	61	222	62
rect	221	64	222	65
rect	221	70	222	71
rect	221	76	222	77
rect	221	82	222	83
rect	221	88	222	89
rect	221	91	222	92
rect	221	94	222	95
rect	221	100	222	101
rect	221	106	222	107
rect	221	109	222	110
rect	221	112	222	113
rect	221	115	222	116
rect	221	121	222	122
rect	221	124	222	125
rect	221	127	222	128
rect	221	136	222	137
rect	221	142	222	143
rect	221	145	222	146
rect	221	151	222	152
rect	221	154	222	155
rect	221	157	222	158
rect	221	166	222	167
rect	221	169	222	170
rect	221	172	222	173
rect	221	175	222	176
rect	221	181	222	182
rect	221	184	222	185
rect	221	187	222	188
rect	221	196	222	197
rect	221	202	222	203
rect	221	205	222	206
rect	221	217	222	218
rect	221	220	222	221
rect	221	229	222	230
rect	221	232	222	233
rect	221	238	222	239
rect	221	244	222	245
rect	221	247	222	248
rect	221	250	222	251
rect	221	253	222	254
rect	221	259	222	260
rect	221	262	222	263
rect	221	271	222	272
rect	221	274	222	275
rect	221	280	222	281
rect	221	286	222	287
rect	221	292	222	293
rect	221	298	222	299
rect	221	301	222	302
rect	221	304	222	305
rect	221	313	222	314
rect	221	316	222	317
rect	221	319	222	320
rect	221	328	222	329
rect	221	331	222	332
rect	221	334	222	335
rect	222	19	223	20
rect	222	25	223	26
rect	222	31	223	32
rect	222	34	223	35
rect	222	40	223	41
rect	222	46	223	47
rect	222	52	223	53
rect	222	61	223	62
rect	222	64	223	65
rect	222	70	223	71
rect	222	76	223	77
rect	222	82	223	83
rect	222	88	223	89
rect	222	91	223	92
rect	222	94	223	95
rect	222	100	223	101
rect	222	106	223	107
rect	222	109	223	110
rect	222	112	223	113
rect	222	115	223	116
rect	222	121	223	122
rect	222	124	223	125
rect	222	127	223	128
rect	222	136	223	137
rect	222	142	223	143
rect	222	145	223	146
rect	222	151	223	152
rect	222	154	223	155
rect	222	157	223	158
rect	222	166	223	167
rect	222	169	223	170
rect	222	172	223	173
rect	222	175	223	176
rect	222	181	223	182
rect	222	184	223	185
rect	222	187	223	188
rect	222	196	223	197
rect	222	202	223	203
rect	222	205	223	206
rect	222	217	223	218
rect	222	220	223	221
rect	222	229	223	230
rect	222	232	223	233
rect	222	244	223	245
rect	222	247	223	248
rect	222	250	223	251
rect	222	253	223	254
rect	222	259	223	260
rect	222	274	223	275
rect	222	280	223	281
rect	222	286	223	287
rect	222	292	223	293
rect	222	298	223	299
rect	222	301	223	302
rect	222	316	223	317
rect	222	319	223	320
rect	222	328	223	329
rect	222	331	223	332
rect	222	334	223	335
rect	223	19	224	20
rect	223	25	224	26
rect	223	31	224	32
rect	223	34	224	35
rect	223	40	224	41
rect	223	46	224	47
rect	223	52	224	53
rect	223	61	224	62
rect	223	64	224	65
rect	223	70	224	71
rect	223	76	224	77
rect	223	82	224	83
rect	223	88	224	89
rect	223	91	224	92
rect	223	94	224	95
rect	223	100	224	101
rect	223	106	224	107
rect	223	109	224	110
rect	223	112	224	113
rect	223	115	224	116
rect	223	121	224	122
rect	223	124	224	125
rect	223	127	224	128
rect	223	136	224	137
rect	223	142	224	143
rect	223	145	224	146
rect	223	151	224	152
rect	223	154	224	155
rect	223	157	224	158
rect	223	166	224	167
rect	223	169	224	170
rect	223	172	224	173
rect	223	175	224	176
rect	223	181	224	182
rect	223	184	224	185
rect	223	187	224	188
rect	223	196	224	197
rect	223	202	224	203
rect	223	205	224	206
rect	223	217	224	218
rect	223	220	224	221
rect	223	229	224	230
rect	223	232	224	233
rect	223	241	224	242
rect	223	244	224	245
rect	223	247	224	248
rect	223	250	224	251
rect	223	253	224	254
rect	223	259	224	260
rect	223	274	224	275
rect	223	277	224	278
rect	223	280	224	281
rect	223	283	224	284
rect	223	286	224	287
rect	223	289	224	290
rect	223	292	224	293
rect	223	295	224	296
rect	223	298	224	299
rect	223	301	224	302
rect	223	316	224	317
rect	223	319	224	320
rect	223	325	224	326
rect	223	328	224	329
rect	223	331	224	332
rect	223	334	224	335
rect	224	19	225	20
rect	224	25	225	26
rect	224	31	225	32
rect	224	34	225	35
rect	224	40	225	41
rect	224	46	225	47
rect	224	52	225	53
rect	224	61	225	62
rect	224	64	225	65
rect	224	70	225	71
rect	224	76	225	77
rect	224	82	225	83
rect	224	88	225	89
rect	224	91	225	92
rect	224	94	225	95
rect	224	100	225	101
rect	224	106	225	107
rect	224	109	225	110
rect	224	112	225	113
rect	224	115	225	116
rect	224	121	225	122
rect	224	124	225	125
rect	224	127	225	128
rect	224	136	225	137
rect	224	142	225	143
rect	224	145	225	146
rect	224	151	225	152
rect	224	154	225	155
rect	224	157	225	158
rect	224	166	225	167
rect	224	169	225	170
rect	224	172	225	173
rect	224	175	225	176
rect	224	181	225	182
rect	224	184	225	185
rect	224	187	225	188
rect	224	196	225	197
rect	224	202	225	203
rect	224	205	225	206
rect	224	217	225	218
rect	224	220	225	221
rect	224	229	225	230
rect	224	232	225	233
rect	224	241	225	242
rect	224	244	225	245
rect	224	247	225	248
rect	224	250	225	251
rect	224	274	225	275
rect	224	277	225	278
rect	224	280	225	281
rect	224	283	225	284
rect	224	286	225	287
rect	224	289	225	290
rect	224	292	225	293
rect	224	295	225	296
rect	224	301	225	302
rect	224	319	225	320
rect	224	325	225	326
rect	224	328	225	329
rect	224	331	225	332
rect	224	334	225	335
rect	225	19	226	20
rect	225	25	226	26
rect	225	28	226	29
rect	225	31	226	32
rect	225	34	226	35
rect	225	40	226	41
rect	225	46	226	47
rect	225	52	226	53
rect	225	61	226	62
rect	225	64	226	65
rect	225	70	226	71
rect	225	76	226	77
rect	225	82	226	83
rect	225	88	226	89
rect	225	91	226	92
rect	225	94	226	95
rect	225	100	226	101
rect	225	106	226	107
rect	225	109	226	110
rect	225	112	226	113
rect	225	115	226	116
rect	225	121	226	122
rect	225	124	226	125
rect	225	127	226	128
rect	225	136	226	137
rect	225	142	226	143
rect	225	145	226	146
rect	225	151	226	152
rect	225	154	226	155
rect	225	157	226	158
rect	225	166	226	167
rect	225	169	226	170
rect	225	172	226	173
rect	225	175	226	176
rect	225	181	226	182
rect	225	184	226	185
rect	225	187	226	188
rect	225	196	226	197
rect	225	202	226	203
rect	225	205	226	206
rect	225	211	226	212
rect	225	217	226	218
rect	225	220	226	221
rect	225	229	226	230
rect	225	232	226	233
rect	225	238	226	239
rect	225	241	226	242
rect	225	244	226	245
rect	225	247	226	248
rect	225	250	226	251
rect	225	265	226	266
rect	225	271	226	272
rect	225	274	226	275
rect	225	277	226	278
rect	225	280	226	281
rect	225	283	226	284
rect	225	286	226	287
rect	225	289	226	290
rect	225	292	226	293
rect	225	295	226	296
rect	225	301	226	302
rect	225	304	226	305
rect	225	319	226	320
rect	225	325	226	326
rect	225	328	226	329
rect	225	331	226	332
rect	225	334	226	335
rect	226	19	227	20
rect	226	28	227	29
rect	226	31	227	32
rect	226	34	227	35
rect	226	40	227	41
rect	226	61	227	62
rect	226	76	227	77
rect	226	82	227	83
rect	226	91	227	92
rect	226	94	227	95
rect	226	100	227	101
rect	226	106	227	107
rect	226	109	227	110
rect	226	112	227	113
rect	226	121	227	122
rect	226	124	227	125
rect	226	127	227	128
rect	226	136	227	137
rect	226	142	227	143
rect	226	151	227	152
rect	226	154	227	155
rect	226	157	227	158
rect	226	169	227	170
rect	226	172	227	173
rect	226	181	227	182
rect	226	184	227	185
rect	226	187	227	188
rect	226	196	227	197
rect	226	202	227	203
rect	226	205	227	206
rect	226	211	227	212
rect	226	217	227	218
rect	226	220	227	221
rect	226	229	227	230
rect	226	238	227	239
rect	226	241	227	242
rect	226	244	227	245
rect	226	247	227	248
rect	226	250	227	251
rect	226	265	227	266
rect	226	271	227	272
rect	226	274	227	275
rect	226	277	227	278
rect	226	280	227	281
rect	226	283	227	284
rect	226	289	227	290
rect	226	292	227	293
rect	226	295	227	296
rect	226	304	227	305
rect	226	319	227	320
rect	226	325	227	326
rect	226	328	227	329
rect	226	331	227	332
rect	226	334	227	335
rect	227	4	228	5
rect	227	7	228	8
rect	227	10	228	11
rect	227	16	228	17
rect	227	19	228	20
rect	227	28	228	29
rect	227	31	228	32
rect	227	34	228	35
rect	227	37	228	38
rect	227	40	228	41
rect	227	49	228	50
rect	227	58	228	59
rect	227	61	228	62
rect	227	67	228	68
rect	227	76	228	77
rect	227	79	228	80
rect	227	82	228	83
rect	227	91	228	92
rect	227	94	228	95
rect	227	97	228	98
rect	227	100	228	101
rect	227	106	228	107
rect	227	109	228	110
rect	227	112	228	113
rect	227	118	228	119
rect	227	121	228	122
rect	227	124	228	125
rect	227	127	228	128
rect	227	136	228	137
rect	227	139	228	140
rect	227	142	228	143
rect	227	151	228	152
rect	227	154	228	155
rect	227	157	228	158
rect	227	160	228	161
rect	227	169	228	170
rect	227	172	228	173
rect	227	181	228	182
rect	227	184	228	185
rect	227	187	228	188
rect	227	196	228	197
rect	227	199	228	200
rect	227	202	228	203
rect	227	205	228	206
rect	227	211	228	212
rect	227	217	228	218
rect	227	220	228	221
rect	227	229	228	230
rect	227	238	228	239
rect	227	241	228	242
rect	227	244	228	245
rect	227	247	228	248
rect	227	250	228	251
rect	227	253	228	254
rect	227	256	228	257
rect	227	262	228	263
rect	227	265	228	266
rect	227	268	228	269
rect	227	271	228	272
rect	227	274	228	275
rect	227	277	228	278
rect	227	280	228	281
rect	227	283	228	284
rect	227	289	228	290
rect	227	292	228	293
rect	227	295	228	296
rect	227	304	228	305
rect	227	313	228	314
rect	227	319	228	320
rect	227	325	228	326
rect	227	328	228	329
rect	227	331	228	332
rect	227	334	228	335
rect	234	1	235	2
rect	234	7	235	8
rect	234	10	235	11
rect	234	13	235	14
rect	234	16	235	17
rect	234	19	235	20
rect	234	28	235	29
rect	234	31	235	32
rect	234	34	235	35
rect	234	37	235	38
rect	234	40	235	41
rect	234	49	235	50
rect	234	58	235	59
rect	234	61	235	62
rect	234	67	235	68
rect	234	73	235	74
rect	234	76	235	77
rect	234	79	235	80
rect	234	82	235	83
rect	234	88	235	89
rect	234	91	235	92
rect	234	94	235	95
rect	234	97	235	98
rect	234	100	235	101
rect	234	103	235	104
rect	234	109	235	110
rect	234	112	235	113
rect	234	121	235	122
rect	234	124	235	125
rect	234	127	235	128
rect	234	136	235	137
rect	234	139	235	140
rect	234	142	235	143
rect	234	145	235	146
rect	234	151	235	152
rect	234	154	235	155
rect	234	157	235	158
rect	234	160	235	161
rect	234	169	235	170
rect	234	172	235	173
rect	234	181	235	182
rect	234	184	235	185
rect	234	187	235	188
rect	234	193	235	194
rect	234	196	235	197
rect	234	199	235	200
rect	234	202	235	203
rect	234	205	235	206
rect	234	214	235	215
rect	234	220	235	221
rect	234	229	235	230
rect	234	238	235	239
rect	234	241	235	242
rect	234	244	235	245
rect	234	247	235	248
rect	234	250	235	251
rect	234	253	235	254
rect	234	262	235	263
rect	234	265	235	266
rect	234	268	235	269
rect	234	271	235	272
rect	234	274	235	275
rect	234	277	235	278
rect	234	280	235	281
rect	234	289	235	290
rect	234	292	235	293
rect	234	295	235	296
rect	234	304	235	305
rect	234	319	235	320
rect	234	322	235	323
rect	234	328	235	329
rect	234	331	235	332
rect	234	334	235	335
rect	235	1	236	2
rect	235	7	236	8
rect	235	10	236	11
rect	235	13	236	14
rect	235	16	236	17
rect	235	19	236	20
rect	235	28	236	29
rect	235	31	236	32
rect	235	34	236	35
rect	235	37	236	38
rect	235	40	236	41
rect	235	49	236	50
rect	235	58	236	59
rect	235	61	236	62
rect	235	67	236	68
rect	235	73	236	74
rect	235	76	236	77
rect	235	79	236	80
rect	235	82	236	83
rect	235	88	236	89
rect	235	91	236	92
rect	235	97	236	98
rect	235	100	236	101
rect	235	103	236	104
rect	235	109	236	110
rect	235	112	236	113
rect	235	121	236	122
rect	235	124	236	125
rect	235	127	236	128
rect	235	136	236	137
rect	235	139	236	140
rect	235	142	236	143
rect	235	145	236	146
rect	235	151	236	152
rect	235	154	236	155
rect	235	157	236	158
rect	235	160	236	161
rect	235	169	236	170
rect	235	172	236	173
rect	235	181	236	182
rect	235	184	236	185
rect	235	187	236	188
rect	235	196	236	197
rect	235	199	236	200
rect	235	202	236	203
rect	235	205	236	206
rect	235	214	236	215
rect	235	220	236	221
rect	235	229	236	230
rect	235	238	236	239
rect	235	241	236	242
rect	235	244	236	245
rect	235	247	236	248
rect	235	250	236	251
rect	235	253	236	254
rect	235	262	236	263
rect	235	265	236	266
rect	235	268	236	269
rect	235	271	236	272
rect	235	274	236	275
rect	235	277	236	278
rect	235	280	236	281
rect	235	289	236	290
rect	235	292	236	293
rect	235	295	236	296
rect	235	304	236	305
rect	235	319	236	320
rect	235	322	236	323
rect	235	328	236	329
rect	235	331	236	332
rect	235	334	236	335
rect	236	1	237	2
rect	236	7	237	8
rect	236	10	237	11
rect	236	13	237	14
rect	236	16	237	17
rect	236	19	237	20
rect	236	28	237	29
rect	236	31	237	32
rect	236	34	237	35
rect	236	37	237	38
rect	236	40	237	41
rect	236	49	237	50
rect	236	58	237	59
rect	236	61	237	62
rect	236	67	237	68
rect	236	73	237	74
rect	236	76	237	77
rect	236	79	237	80
rect	236	82	237	83
rect	236	88	237	89
rect	236	91	237	92
rect	236	97	237	98
rect	236	100	237	101
rect	236	103	237	104
rect	236	109	237	110
rect	236	112	237	113
rect	236	118	237	119
rect	236	121	237	122
rect	236	124	237	125
rect	236	127	237	128
rect	236	136	237	137
rect	236	139	237	140
rect	236	142	237	143
rect	236	145	237	146
rect	236	151	237	152
rect	236	154	237	155
rect	236	157	237	158
rect	236	160	237	161
rect	236	169	237	170
rect	236	172	237	173
rect	236	181	237	182
rect	236	184	237	185
rect	236	187	237	188
rect	236	196	237	197
rect	236	199	237	200
rect	236	202	237	203
rect	236	205	237	206
rect	236	214	237	215
rect	236	217	237	218
rect	236	220	237	221
rect	236	229	237	230
rect	236	238	237	239
rect	236	241	237	242
rect	236	244	237	245
rect	236	247	237	248
rect	236	250	237	251
rect	236	253	237	254
rect	236	262	237	263
rect	236	265	237	266
rect	236	268	237	269
rect	236	271	237	272
rect	236	274	237	275
rect	236	277	237	278
rect	236	280	237	281
rect	236	289	237	290
rect	236	292	237	293
rect	236	295	237	296
rect	236	304	237	305
rect	236	319	237	320
rect	236	322	237	323
rect	236	328	237	329
rect	236	331	237	332
rect	236	334	237	335
rect	237	1	238	2
rect	237	7	238	8
rect	237	10	238	11
rect	237	13	238	14
rect	237	16	238	17
rect	237	28	238	29
rect	237	31	238	32
rect	237	34	238	35
rect	237	37	238	38
rect	237	40	238	41
rect	237	49	238	50
rect	237	58	238	59
rect	237	61	238	62
rect	237	67	238	68
rect	237	73	238	74
rect	237	79	238	80
rect	237	82	238	83
rect	237	88	238	89
rect	237	91	238	92
rect	237	97	238	98
rect	237	100	238	101
rect	237	103	238	104
rect	237	109	238	110
rect	237	112	238	113
rect	237	118	238	119
rect	237	121	238	122
rect	237	124	238	125
rect	237	127	238	128
rect	237	136	238	137
rect	237	139	238	140
rect	237	142	238	143
rect	237	145	238	146
rect	237	151	238	152
rect	237	154	238	155
rect	237	157	238	158
rect	237	160	238	161
rect	237	172	238	173
rect	237	181	238	182
rect	237	184	238	185
rect	237	187	238	188
rect	237	196	238	197
rect	237	199	238	200
rect	237	202	238	203
rect	237	205	238	206
rect	237	214	238	215
rect	237	217	238	218
rect	237	220	238	221
rect	237	229	238	230
rect	237	238	238	239
rect	237	241	238	242
rect	237	244	238	245
rect	237	247	238	248
rect	237	250	238	251
rect	237	253	238	254
rect	237	262	238	263
rect	237	265	238	266
rect	237	268	238	269
rect	237	271	238	272
rect	237	274	238	275
rect	237	277	238	278
rect	237	280	238	281
rect	237	289	238	290
rect	237	292	238	293
rect	237	295	238	296
rect	237	304	238	305
rect	237	319	238	320
rect	237	322	238	323
rect	237	328	238	329
rect	237	331	238	332
rect	237	334	238	335
rect	238	1	239	2
rect	238	5	239	6
rect	238	7	239	8
rect	238	10	239	11
rect	238	13	239	14
rect	238	16	239	17
rect	238	28	239	29
rect	238	31	239	32
rect	238	34	239	35
rect	238	37	239	38
rect	238	40	239	41
rect	238	49	239	50
rect	238	58	239	59
rect	238	61	239	62
rect	238	67	239	68
rect	238	73	239	74
rect	238	79	239	80
rect	238	82	239	83
rect	238	88	239	89
rect	238	91	239	92
rect	238	94	239	95
rect	238	97	239	98
rect	238	100	239	101
rect	238	103	239	104
rect	238	109	239	110
rect	238	112	239	113
rect	238	118	239	119
rect	238	121	239	122
rect	238	124	239	125
rect	238	127	239	128
rect	238	136	239	137
rect	238	139	239	140
rect	238	142	239	143
rect	238	145	239	146
rect	238	151	239	152
rect	238	154	239	155
rect	238	157	239	158
rect	238	160	239	161
rect	238	172	239	173
rect	238	181	239	182
rect	238	184	239	185
rect	238	187	239	188
rect	238	193	239	194
rect	238	196	239	197
rect	238	199	239	200
rect	238	202	239	203
rect	238	205	239	206
rect	238	214	239	215
rect	238	217	239	218
rect	238	220	239	221
rect	238	229	239	230
rect	238	238	239	239
rect	238	241	239	242
rect	238	244	239	245
rect	238	247	239	248
rect	238	250	239	251
rect	238	253	239	254
rect	238	262	239	263
rect	238	265	239	266
rect	238	268	239	269
rect	238	271	239	272
rect	238	274	239	275
rect	238	277	239	278
rect	238	280	239	281
rect	238	289	239	290
rect	238	292	239	293
rect	238	295	239	296
rect	238	304	239	305
rect	238	319	239	320
rect	238	322	239	323
rect	238	328	239	329
rect	238	331	239	332
rect	238	334	239	335
rect	239	1	240	2
rect	239	5	240	6
rect	239	7	240	8
rect	239	10	240	11
rect	239	13	240	14
rect	239	16	240	17
rect	239	28	240	29
rect	239	31	240	32
rect	239	34	240	35
rect	239	40	240	41
rect	239	49	240	50
rect	239	58	240	59
rect	239	61	240	62
rect	239	73	240	74
rect	239	79	240	80
rect	239	82	240	83
rect	239	88	240	89
rect	239	91	240	92
rect	239	94	240	95
rect	239	97	240	98
rect	239	100	240	101
rect	239	103	240	104
rect	239	109	240	110
rect	239	112	240	113
rect	239	118	240	119
rect	239	121	240	122
rect	239	124	240	125
rect	239	127	240	128
rect	239	136	240	137
rect	239	139	240	140
rect	239	142	240	143
rect	239	145	240	146
rect	239	151	240	152
rect	239	157	240	158
rect	239	160	240	161
rect	239	172	240	173
rect	239	181	240	182
rect	239	184	240	185
rect	239	187	240	188
rect	239	193	240	194
rect	239	196	240	197
rect	239	199	240	200
rect	239	202	240	203
rect	239	205	240	206
rect	239	214	240	215
rect	239	217	240	218
rect	239	220	240	221
rect	239	229	240	230
rect	239	238	240	239
rect	239	241	240	242
rect	239	244	240	245
rect	239	247	240	248
rect	239	250	240	251
rect	239	253	240	254
rect	239	262	240	263
rect	239	265	240	266
rect	239	268	240	269
rect	239	271	240	272
rect	239	274	240	275
rect	239	277	240	278
rect	239	280	240	281
rect	239	289	240	290
rect	239	292	240	293
rect	239	295	240	296
rect	239	304	240	305
rect	239	319	240	320
rect	239	322	240	323
rect	239	328	240	329
rect	239	331	240	332
rect	239	334	240	335
rect	240	1	241	2
rect	240	5	241	6
rect	240	7	241	8
rect	240	10	241	11
rect	240	13	241	14
rect	240	16	241	17
rect	240	19	241	20
rect	240	28	241	29
rect	240	31	241	32
rect	240	34	241	35
rect	240	40	241	41
rect	240	49	241	50
rect	240	58	241	59
rect	240	61	241	62
rect	240	73	241	74
rect	240	76	241	77
rect	240	79	241	80
rect	240	82	241	83
rect	240	88	241	89
rect	240	91	241	92
rect	240	94	241	95
rect	240	97	241	98
rect	240	100	241	101
rect	240	103	241	104
rect	240	109	241	110
rect	240	112	241	113
rect	240	118	241	119
rect	240	121	241	122
rect	240	124	241	125
rect	240	127	241	128
rect	240	136	241	137
rect	240	139	241	140
rect	240	142	241	143
rect	240	145	241	146
rect	240	151	241	152
rect	240	157	241	158
rect	240	160	241	161
rect	240	172	241	173
rect	240	175	241	176
rect	240	181	241	182
rect	240	184	241	185
rect	240	187	241	188
rect	240	193	241	194
rect	240	196	241	197
rect	240	199	241	200
rect	240	202	241	203
rect	240	205	241	206
rect	240	214	241	215
rect	240	217	241	218
rect	240	220	241	221
rect	240	229	241	230
rect	240	238	241	239
rect	240	241	241	242
rect	240	244	241	245
rect	240	247	241	248
rect	240	250	241	251
rect	240	253	241	254
rect	240	262	241	263
rect	240	265	241	266
rect	240	268	241	269
rect	240	271	241	272
rect	240	274	241	275
rect	240	277	241	278
rect	240	280	241	281
rect	240	289	241	290
rect	240	292	241	293
rect	240	295	241	296
rect	240	304	241	305
rect	240	319	241	320
rect	240	322	241	323
rect	240	328	241	329
rect	240	331	241	332
rect	240	334	241	335
rect	241	1	242	2
rect	241	5	242	6
rect	241	7	242	8
rect	241	10	242	11
rect	241	13	242	14
rect	241	19	242	20
rect	241	28	242	29
rect	241	31	242	32
rect	241	34	242	35
rect	241	40	242	41
rect	241	49	242	50
rect	241	58	242	59
rect	241	61	242	62
rect	241	76	242	77
rect	241	79	242	80
rect	241	82	242	83
rect	241	88	242	89
rect	241	91	242	92
rect	241	94	242	95
rect	241	97	242	98
rect	241	100	242	101
rect	241	103	242	104
rect	241	109	242	110
rect	241	112	242	113
rect	241	118	242	119
rect	241	121	242	122
rect	241	124	242	125
rect	241	127	242	128
rect	241	139	242	140
rect	241	142	242	143
rect	241	145	242	146
rect	241	151	242	152
rect	241	157	242	158
rect	241	160	242	161
rect	241	172	242	173
rect	241	175	242	176
rect	241	184	242	185
rect	241	187	242	188
rect	241	193	242	194
rect	241	196	242	197
rect	241	199	242	200
rect	241	202	242	203
rect	241	205	242	206
rect	241	214	242	215
rect	241	217	242	218
rect	241	220	242	221
rect	241	229	242	230
rect	241	238	242	239
rect	241	241	242	242
rect	241	244	242	245
rect	241	247	242	248
rect	241	250	242	251
rect	241	253	242	254
rect	241	262	242	263
rect	241	265	242	266
rect	241	268	242	269
rect	241	271	242	272
rect	241	274	242	275
rect	241	280	242	281
rect	241	292	242	293
rect	241	295	242	296
rect	241	304	242	305
rect	241	319	242	320
rect	241	322	242	323
rect	241	328	242	329
rect	241	331	242	332
rect	242	1	243	2
rect	242	5	243	6
rect	242	7	243	8
rect	242	10	243	11
rect	242	13	243	14
rect	242	19	243	20
rect	242	28	243	29
rect	242	31	243	32
rect	242	34	243	35
rect	242	37	243	38
rect	242	40	243	41
rect	242	49	243	50
rect	242	58	243	59
rect	242	61	243	62
rect	242	67	243	68
rect	242	76	243	77
rect	242	79	243	80
rect	242	82	243	83
rect	242	88	243	89
rect	242	91	243	92
rect	242	94	243	95
rect	242	97	243	98
rect	242	100	243	101
rect	242	103	243	104
rect	242	109	243	110
rect	242	112	243	113
rect	242	118	243	119
rect	242	121	243	122
rect	242	124	243	125
rect	242	127	243	128
rect	242	139	243	140
rect	242	142	243	143
rect	242	145	243	146
rect	242	151	243	152
rect	242	157	243	158
rect	242	160	243	161
rect	242	169	243	170
rect	242	172	243	173
rect	242	175	243	176
rect	242	184	243	185
rect	242	187	243	188
rect	242	190	243	191
rect	242	193	243	194
rect	242	196	243	197
rect	242	199	243	200
rect	242	202	243	203
rect	242	205	243	206
rect	242	214	243	215
rect	242	217	243	218
rect	242	220	243	221
rect	242	229	243	230
rect	242	238	243	239
rect	242	241	243	242
rect	242	244	243	245
rect	242	247	243	248
rect	242	250	243	251
rect	242	253	243	254
rect	242	262	243	263
rect	242	265	243	266
rect	242	268	243	269
rect	242	271	243	272
rect	242	274	243	275
rect	242	280	243	281
rect	242	283	243	284
rect	242	292	243	293
rect	242	295	243	296
rect	242	304	243	305
rect	242	310	243	311
rect	242	319	243	320
rect	242	322	243	323
rect	242	328	243	329
rect	242	331	243	332
rect	242	337	243	338
rect	243	1	244	2
rect	243	7	244	8
rect	243	10	244	11
rect	243	13	244	14
rect	243	19	244	20
rect	243	28	244	29
rect	243	31	244	32
rect	243	34	244	35
rect	243	37	244	38
rect	243	49	244	50
rect	243	58	244	59
rect	243	67	244	68
rect	243	76	244	77
rect	243	79	244	80
rect	243	82	244	83
rect	243	88	244	89
rect	243	91	244	92
rect	243	94	244	95
rect	243	97	244	98
rect	243	100	244	101
rect	243	109	244	110
rect	243	112	244	113
rect	243	118	244	119
rect	243	121	244	122
rect	243	124	244	125
rect	243	139	244	140
rect	243	142	244	143
rect	243	145	244	146
rect	243	151	244	152
rect	243	160	244	161
rect	243	169	244	170
rect	243	175	244	176
rect	243	184	244	185
rect	243	187	244	188
rect	243	190	244	191
rect	243	193	244	194
rect	243	196	244	197
rect	243	199	244	200
rect	243	202	244	203
rect	243	214	244	215
rect	243	217	244	218
rect	243	220	244	221
rect	243	238	244	239
rect	243	241	244	242
rect	243	244	244	245
rect	243	247	244	248
rect	243	250	244	251
rect	243	253	244	254
rect	243	265	244	266
rect	243	268	244	269
rect	243	271	244	272
rect	243	274	244	275
rect	243	280	244	281
rect	243	283	244	284
rect	243	292	244	293
rect	243	295	244	296
rect	243	304	244	305
rect	243	310	244	311
rect	243	319	244	320
rect	243	322	244	323
rect	243	328	244	329
rect	243	337	244	338
rect	244	1	245	2
rect	244	7	245	8
rect	244	10	245	11
rect	244	13	245	14
rect	244	16	245	17
rect	244	19	245	20
rect	244	22	245	23
rect	244	28	245	29
rect	244	31	245	32
rect	244	34	245	35
rect	244	37	245	38
rect	244	49	245	50
rect	244	58	245	59
rect	244	67	245	68
rect	244	73	245	74
rect	244	76	245	77
rect	244	79	245	80
rect	244	82	245	83
rect	244	88	245	89
rect	244	91	245	92
rect	244	94	245	95
rect	244	97	245	98
rect	244	100	245	101
rect	244	109	245	110
rect	244	112	245	113
rect	244	115	245	116
rect	244	118	245	119
rect	244	121	245	122
rect	244	124	245	125
rect	244	136	245	137
rect	244	139	245	140
rect	244	142	245	143
rect	244	145	245	146
rect	244	151	245	152
rect	244	154	245	155
rect	244	160	245	161
rect	244	169	245	170
rect	244	175	245	176
rect	244	181	245	182
rect	244	184	245	185
rect	244	187	245	188
rect	244	190	245	191
rect	244	193	245	194
rect	244	196	245	197
rect	244	199	245	200
rect	244	202	245	203
rect	244	208	245	209
rect	244	214	245	215
rect	244	217	245	218
rect	244	220	245	221
rect	244	232	245	233
rect	244	238	245	239
rect	244	241	245	242
rect	244	244	245	245
rect	244	247	245	248
rect	244	250	245	251
rect	244	253	245	254
rect	244	265	245	266
rect	244	268	245	269
rect	244	271	245	272
rect	244	274	245	275
rect	244	280	245	281
rect	244	283	245	284
rect	244	292	245	293
rect	244	295	245	296
rect	244	298	245	299
rect	244	304	245	305
rect	244	310	245	311
rect	244	319	245	320
rect	244	322	245	323
rect	244	328	245	329
rect	244	337	245	338
rect	244	355	245	356
rect	245	1	246	2
rect	245	7	246	8
rect	245	10	246	11
rect	245	16	246	17
rect	245	19	246	20
rect	245	22	246	23
rect	245	28	246	29
rect	245	31	246	32
rect	245	34	246	35
rect	245	37	246	38
rect	245	49	246	50
rect	245	58	246	59
rect	245	67	246	68
rect	245	73	246	74
rect	245	76	246	77
rect	245	79	246	80
rect	245	82	246	83
rect	245	88	246	89
rect	245	91	246	92
rect	245	94	246	95
rect	245	97	246	98
rect	245	100	246	101
rect	245	109	246	110
rect	245	112	246	113
rect	245	115	246	116
rect	245	118	246	119
rect	245	121	246	122
rect	245	124	246	125
rect	245	136	246	137
rect	245	139	246	140
rect	245	142	246	143
rect	245	145	246	146
rect	245	154	246	155
rect	245	160	246	161
rect	245	169	246	170
rect	245	175	246	176
rect	245	181	246	182
rect	245	184	246	185
rect	245	187	246	188
rect	245	190	246	191
rect	245	193	246	194
rect	245	196	246	197
rect	245	199	246	200
rect	245	208	246	209
rect	245	217	246	218
rect	245	232	246	233
rect	245	238	246	239
rect	245	241	246	242
rect	245	244	246	245
rect	245	247	246	248
rect	245	250	246	251
rect	245	265	246	266
rect	245	268	246	269
rect	245	271	246	272
rect	245	283	246	284
rect	245	292	246	293
rect	245	298	246	299
rect	245	304	246	305
rect	245	310	246	311
rect	245	319	246	320
rect	245	328	246	329
rect	245	337	246	338
rect	245	355	246	356
rect	246	1	247	2
rect	246	7	247	8
rect	246	10	247	11
rect	246	16	247	17
rect	246	19	247	20
rect	246	22	247	23
rect	246	28	247	29
rect	246	31	247	32
rect	246	34	247	35
rect	246	37	247	38
rect	246	49	247	50
rect	246	58	247	59
rect	246	67	247	68
rect	246	73	247	74
rect	246	76	247	77
rect	246	79	247	80
rect	246	82	247	83
rect	246	88	247	89
rect	246	91	247	92
rect	246	94	247	95
rect	246	97	247	98
rect	246	100	247	101
rect	246	109	247	110
rect	246	112	247	113
rect	246	115	247	116
rect	246	118	247	119
rect	246	121	247	122
rect	246	124	247	125
rect	246	133	247	134
rect	246	136	247	137
rect	246	139	247	140
rect	246	142	247	143
rect	246	145	247	146
rect	246	154	247	155
rect	246	160	247	161
rect	246	169	247	170
rect	246	172	247	173
rect	246	175	247	176
rect	246	181	247	182
rect	246	184	247	185
rect	246	187	247	188
rect	246	190	247	191
rect	246	193	247	194
rect	246	196	247	197
rect	246	199	247	200
rect	246	208	247	209
rect	246	217	247	218
rect	246	229	247	230
rect	246	232	247	233
rect	246	238	247	239
rect	246	241	247	242
rect	246	244	247	245
rect	246	247	247	248
rect	246	250	247	251
rect	246	262	247	263
rect	246	265	247	266
rect	246	268	247	269
rect	246	271	247	272
rect	246	277	247	278
rect	246	283	247	284
rect	246	286	247	287
rect	246	289	247	290
rect	246	292	247	293
rect	246	298	247	299
rect	246	304	247	305
rect	246	310	247	311
rect	246	319	247	320
rect	246	328	247	329
rect	246	337	247	338
rect	246	352	247	353
rect	246	355	247	356
rect	247	1	248	2
rect	247	10	248	11
rect	247	16	248	17
rect	247	19	248	20
rect	247	22	248	23
rect	247	28	248	29
rect	247	34	248	35
rect	247	37	248	38
rect	247	49	248	50
rect	247	58	248	59
rect	247	67	248	68
rect	247	73	248	74
rect	247	76	248	77
rect	247	79	248	80
rect	247	82	248	83
rect	247	88	248	89
rect	247	91	248	92
rect	247	94	248	95
rect	247	97	248	98
rect	247	109	248	110
rect	247	115	248	116
rect	247	118	248	119
rect	247	121	248	122
rect	247	133	248	134
rect	247	136	248	137
rect	247	139	248	140
rect	247	142	248	143
rect	247	145	248	146
rect	247	154	248	155
rect	247	169	248	170
rect	247	172	248	173
rect	247	175	248	176
rect	247	181	248	182
rect	247	184	248	185
rect	247	187	248	188
rect	247	190	248	191
rect	247	193	248	194
rect	247	199	248	200
rect	247	208	248	209
rect	247	217	248	218
rect	247	229	248	230
rect	247	232	248	233
rect	247	238	248	239
rect	247	244	248	245
rect	247	247	248	248
rect	247	250	248	251
rect	247	262	248	263
rect	247	265	248	266
rect	247	271	248	272
rect	247	277	248	278
rect	247	283	248	284
rect	247	286	248	287
rect	247	289	248	290
rect	247	298	248	299
rect	247	304	248	305
rect	247	310	248	311
rect	247	337	248	338
rect	247	352	248	353
rect	247	355	248	356
rect	248	1	249	2
rect	248	10	249	11
rect	248	13	249	14
rect	248	16	249	17
rect	248	19	249	20
rect	248	22	249	23
rect	248	28	249	29
rect	248	34	249	35
rect	248	37	249	38
rect	248	40	249	41
rect	248	49	249	50
rect	248	58	249	59
rect	248	61	249	62
rect	248	64	249	65
rect	248	67	249	68
rect	248	73	249	74
rect	248	76	249	77
rect	248	79	249	80
rect	248	82	249	83
rect	248	88	249	89
rect	248	91	249	92
rect	248	94	249	95
rect	248	97	249	98
rect	248	103	249	104
rect	248	106	249	107
rect	248	109	249	110
rect	248	115	249	116
rect	248	118	249	119
rect	248	121	249	122
rect	248	133	249	134
rect	248	136	249	137
rect	248	139	249	140
rect	248	142	249	143
rect	248	145	249	146
rect	248	151	249	152
rect	248	154	249	155
rect	248	157	249	158
rect	248	169	249	170
rect	248	172	249	173
rect	248	175	249	176
rect	248	181	249	182
rect	248	184	249	185
rect	248	187	249	188
rect	248	190	249	191
rect	248	193	249	194
rect	248	199	249	200
rect	248	208	249	209
rect	248	217	249	218
rect	248	220	249	221
rect	248	229	249	230
rect	248	232	249	233
rect	248	238	249	239
rect	248	244	249	245
rect	248	247	249	248
rect	248	250	249	251
rect	248	256	249	257
rect	248	262	249	263
rect	248	265	249	266
rect	248	271	249	272
rect	248	274	249	275
rect	248	277	249	278
rect	248	280	249	281
rect	248	283	249	284
rect	248	286	249	287
rect	248	289	249	290
rect	248	298	249	299
rect	248	304	249	305
rect	248	310	249	311
rect	248	325	249	326
rect	248	337	249	338
rect	248	352	249	353
rect	248	355	249	356
rect	248	364	249	365
rect	249	13	250	14
rect	249	16	250	17
rect	249	19	250	20
rect	249	22	250	23
rect	249	28	250	29
rect	249	34	250	35
rect	249	37	250	38
rect	249	40	250	41
rect	249	49	250	50
rect	249	58	250	59
rect	249	61	250	62
rect	249	64	250	65
rect	249	67	250	68
rect	249	73	250	74
rect	249	76	250	77
rect	249	79	250	80
rect	249	82	250	83
rect	249	88	250	89
rect	249	91	250	92
rect	249	94	250	95
rect	249	97	250	98
rect	249	103	250	104
rect	249	106	250	107
rect	249	115	250	116
rect	249	118	250	119
rect	249	133	250	134
rect	249	136	250	137
rect	249	139	250	140
rect	249	142	250	143
rect	249	151	250	152
rect	249	154	250	155
rect	249	157	250	158
rect	249	169	250	170
rect	249	172	250	173
rect	249	175	250	176
rect	249	181	250	182
rect	249	190	250	191
rect	249	193	250	194
rect	249	208	250	209
rect	249	217	250	218
rect	249	220	250	221
rect	249	229	250	230
rect	249	232	250	233
rect	249	244	250	245
rect	249	247	250	248
rect	249	256	250	257
rect	249	262	250	263
rect	249	271	250	272
rect	249	274	250	275
rect	249	277	250	278
rect	249	280	250	281
rect	249	283	250	284
rect	249	286	250	287
rect	249	289	250	290
rect	249	298	250	299
rect	249	310	250	311
rect	249	325	250	326
rect	249	337	250	338
rect	249	352	250	353
rect	249	355	250	356
rect	249	364	250	365
rect	250	7	251	8
rect	250	13	251	14
rect	250	16	251	17
rect	250	19	251	20
rect	250	22	251	23
rect	250	28	251	29
rect	250	34	251	35
rect	250	37	251	38
rect	250	40	251	41
rect	250	49	251	50
rect	250	58	251	59
rect	250	61	251	62
rect	250	64	251	65
rect	250	67	251	68
rect	250	73	251	74
rect	250	76	251	77
rect	250	79	251	80
rect	250	82	251	83
rect	250	88	251	89
rect	250	91	251	92
rect	250	94	251	95
rect	250	97	251	98
rect	250	103	251	104
rect	250	106	251	107
rect	250	115	251	116
rect	250	118	251	119
rect	250	127	251	128
rect	250	133	251	134
rect	250	136	251	137
rect	250	139	251	140
rect	250	142	251	143
rect	250	151	251	152
rect	250	154	251	155
rect	250	157	251	158
rect	250	166	251	167
rect	250	169	251	170
rect	250	172	251	173
rect	250	175	251	176
rect	250	178	251	179
rect	250	181	251	182
rect	250	190	251	191
rect	250	193	251	194
rect	250	196	251	197
rect	250	205	251	206
rect	250	208	251	209
rect	250	217	251	218
rect	250	220	251	221
rect	250	223	251	224
rect	250	226	251	227
rect	250	229	251	230
rect	250	232	251	233
rect	250	241	251	242
rect	250	244	251	245
rect	250	247	251	248
rect	250	256	251	257
rect	250	259	251	260
rect	250	262	251	263
rect	250	271	251	272
rect	250	274	251	275
rect	250	277	251	278
rect	250	280	251	281
rect	250	283	251	284
rect	250	286	251	287
rect	250	289	251	290
rect	250	298	251	299
rect	250	301	251	302
rect	250	310	251	311
rect	250	319	251	320
rect	250	322	251	323
rect	250	325	251	326
rect	250	337	251	338
rect	250	349	251	350
rect	250	352	251	353
rect	250	355	251	356
rect	250	364	251	365
rect	251	7	252	8
rect	251	13	252	14
rect	251	16	252	17
rect	251	19	252	20
rect	251	22	252	23
rect	251	34	252	35
rect	251	37	252	38
rect	251	40	252	41
rect	251	61	252	62
rect	251	64	252	65
rect	251	67	252	68
rect	251	73	252	74
rect	251	76	252	77
rect	251	79	252	80
rect	251	82	252	83
rect	251	91	252	92
rect	251	94	252	95
rect	251	97	252	98
rect	251	103	252	104
rect	251	106	252	107
rect	251	115	252	116
rect	251	118	252	119
rect	251	127	252	128
rect	251	133	252	134
rect	251	136	252	137
rect	251	139	252	140
rect	251	142	252	143
rect	251	151	252	152
rect	251	154	252	155
rect	251	157	252	158
rect	251	166	252	167
rect	251	169	252	170
rect	251	172	252	173
rect	251	175	252	176
rect	251	178	252	179
rect	251	181	252	182
rect	251	190	252	191
rect	251	193	252	194
rect	251	196	252	197
rect	251	205	252	206
rect	251	208	252	209
rect	251	217	252	218
rect	251	220	252	221
rect	251	223	252	224
rect	251	226	252	227
rect	251	229	252	230
rect	251	232	252	233
rect	251	241	252	242
rect	251	244	252	245
rect	251	247	252	248
rect	251	256	252	257
rect	251	259	252	260
rect	251	262	252	263
rect	251	271	252	272
rect	251	274	252	275
rect	251	277	252	278
rect	251	280	252	281
rect	251	283	252	284
rect	251	286	252	287
rect	251	289	252	290
rect	251	298	252	299
rect	251	301	252	302
rect	251	310	252	311
rect	251	319	252	320
rect	251	322	252	323
rect	251	325	252	326
rect	251	337	252	338
rect	251	349	252	350
rect	251	352	252	353
rect	251	355	252	356
rect	251	364	252	365
rect	252	1	253	2
rect	252	7	253	8
rect	252	10	253	11
rect	252	13	253	14
rect	252	16	253	17
rect	252	19	253	20
rect	252	22	253	23
rect	252	31	253	32
rect	252	34	253	35
rect	252	37	253	38
rect	252	40	253	41
rect	252	55	253	56
rect	252	61	253	62
rect	252	64	253	65
rect	252	67	253	68
rect	252	70	253	71
rect	252	73	253	74
rect	252	76	253	77
rect	252	79	253	80
rect	252	82	253	83
rect	252	91	253	92
rect	252	94	253	95
rect	252	97	253	98
rect	252	100	253	101
rect	252	103	253	104
rect	252	106	253	107
rect	252	112	253	113
rect	252	115	253	116
rect	252	118	253	119
rect	252	127	253	128
rect	252	133	253	134
rect	252	136	253	137
rect	252	139	253	140
rect	252	142	253	143
rect	252	151	253	152
rect	252	154	253	155
rect	252	157	253	158
rect	252	166	253	167
rect	252	169	253	170
rect	252	172	253	173
rect	252	175	253	176
rect	252	178	253	179
rect	252	181	253	182
rect	252	190	253	191
rect	252	193	253	194
rect	252	196	253	197
rect	252	205	253	206
rect	252	208	253	209
rect	252	217	253	218
rect	252	220	253	221
rect	252	223	253	224
rect	252	226	253	227
rect	252	229	253	230
rect	252	232	253	233
rect	252	241	253	242
rect	252	244	253	245
rect	252	247	253	248
rect	252	256	253	257
rect	252	259	253	260
rect	252	262	253	263
rect	252	271	253	272
rect	252	274	253	275
rect	252	277	253	278
rect	252	280	253	281
rect	252	283	253	284
rect	252	286	253	287
rect	252	289	253	290
rect	252	298	253	299
rect	252	301	253	302
rect	252	310	253	311
rect	252	319	253	320
rect	252	322	253	323
rect	252	325	253	326
rect	252	334	253	335
rect	252	337	253	338
rect	252	349	253	350
rect	252	352	253	353
rect	252	355	253	356
rect	252	364	253	365
rect	259	7	260	8
rect	259	10	260	11
rect	259	13	260	14
rect	259	16	260	17
rect	259	19	260	20
rect	259	22	260	23
rect	259	28	260	29
rect	259	31	260	32
rect	259	34	260	35
rect	259	37	260	38
rect	259	40	260	41
rect	259	55	260	56
rect	259	64	260	65
rect	259	67	260	68
rect	259	70	260	71
rect	259	73	260	74
rect	259	76	260	77
rect	259	79	260	80
rect	259	82	260	83
rect	259	91	260	92
rect	259	94	260	95
rect	259	97	260	98
rect	259	100	260	101
rect	259	103	260	104
rect	259	106	260	107
rect	259	115	260	116
rect	259	118	260	119
rect	259	130	260	131
rect	259	133	260	134
rect	259	136	260	137
rect	259	139	260	140
rect	259	142	260	143
rect	259	148	260	149
rect	259	151	260	152
rect	259	154	260	155
rect	259	157	260	158
rect	259	166	260	167
rect	259	169	260	170
rect	259	172	260	173
rect	259	175	260	176
rect	259	178	260	179
rect	259	181	260	182
rect	259	190	260	191
rect	259	193	260	194
rect	259	196	260	197
rect	259	205	260	206
rect	259	208	260	209
rect	259	217	260	218
rect	259	226	260	227
rect	259	229	260	230
rect	259	232	260	233
rect	259	238	260	239
rect	259	241	260	242
rect	259	244	260	245
rect	259	247	260	248
rect	259	253	260	254
rect	259	256	260	257
rect	259	259	260	260
rect	259	262	260	263
rect	259	271	260	272
rect	259	274	260	275
rect	259	277	260	278
rect	259	280	260	281
rect	259	283	260	284
rect	259	286	260	287
rect	259	289	260	290
rect	259	298	260	299
rect	259	301	260	302
rect	259	307	260	308
rect	259	310	260	311
rect	259	316	260	317
rect	259	319	260	320
rect	259	322	260	323
rect	259	325	260	326
rect	259	328	260	329
rect	259	334	260	335
rect	259	337	260	338
rect	259	352	260	353
rect	259	355	260	356
rect	259	364	260	365
rect	260	7	261	8
rect	260	10	261	11
rect	260	13	261	14
rect	260	16	261	17
rect	260	19	261	20
rect	260	22	261	23
rect	260	28	261	29
rect	260	31	261	32
rect	260	34	261	35
rect	260	37	261	38
rect	260	40	261	41
rect	260	55	261	56
rect	260	64	261	65
rect	260	67	261	68
rect	260	70	261	71
rect	260	73	261	74
rect	260	76	261	77
rect	260	79	261	80
rect	260	82	261	83
rect	260	91	261	92
rect	260	94	261	95
rect	260	97	261	98
rect	260	100	261	101
rect	260	103	261	104
rect	260	106	261	107
rect	260	115	261	116
rect	260	118	261	119
rect	260	130	261	131
rect	260	133	261	134
rect	260	136	261	137
rect	260	139	261	140
rect	260	142	261	143
rect	260	148	261	149
rect	260	151	261	152
rect	260	154	261	155
rect	260	157	261	158
rect	260	166	261	167
rect	260	169	261	170
rect	260	172	261	173
rect	260	175	261	176
rect	260	178	261	179
rect	260	181	261	182
rect	260	190	261	191
rect	260	193	261	194
rect	260	196	261	197
rect	260	205	261	206
rect	260	208	261	209
rect	260	217	261	218
rect	260	226	261	227
rect	260	229	261	230
rect	260	232	261	233
rect	260	238	261	239
rect	260	241	261	242
rect	260	244	261	245
rect	260	247	261	248
rect	260	253	261	254
rect	260	256	261	257
rect	260	259	261	260
rect	260	262	261	263
rect	260	271	261	272
rect	260	274	261	275
rect	260	277	261	278
rect	260	280	261	281
rect	260	283	261	284
rect	260	286	261	287
rect	260	289	261	290
rect	260	301	261	302
rect	260	307	261	308
rect	260	310	261	311
rect	260	316	261	317
rect	260	319	261	320
rect	260	322	261	323
rect	260	325	261	326
rect	260	328	261	329
rect	260	334	261	335
rect	260	337	261	338
rect	260	352	261	353
rect	260	355	261	356
rect	260	364	261	365
rect	261	7	262	8
rect	261	10	262	11
rect	261	13	262	14
rect	261	16	262	17
rect	261	19	262	20
rect	261	22	262	23
rect	261	28	262	29
rect	261	31	262	32
rect	261	34	262	35
rect	261	37	262	38
rect	261	40	262	41
rect	261	55	262	56
rect	261	64	262	65
rect	261	67	262	68
rect	261	70	262	71
rect	261	73	262	74
rect	261	76	262	77
rect	261	79	262	80
rect	261	82	262	83
rect	261	91	262	92
rect	261	94	262	95
rect	261	97	262	98
rect	261	100	262	101
rect	261	103	262	104
rect	261	106	262	107
rect	261	115	262	116
rect	261	118	262	119
rect	261	130	262	131
rect	261	133	262	134
rect	261	136	262	137
rect	261	139	262	140
rect	261	142	262	143
rect	261	148	262	149
rect	261	151	262	152
rect	261	154	262	155
rect	261	157	262	158
rect	261	166	262	167
rect	261	169	262	170
rect	261	172	262	173
rect	261	175	262	176
rect	261	178	262	179
rect	261	181	262	182
rect	261	190	262	191
rect	261	193	262	194
rect	261	196	262	197
rect	261	205	262	206
rect	261	208	262	209
rect	261	217	262	218
rect	261	226	262	227
rect	261	229	262	230
rect	261	232	262	233
rect	261	238	262	239
rect	261	241	262	242
rect	261	244	262	245
rect	261	247	262	248
rect	261	253	262	254
rect	261	256	262	257
rect	261	259	262	260
rect	261	262	262	263
rect	261	271	262	272
rect	261	274	262	275
rect	261	277	262	278
rect	261	280	262	281
rect	261	283	262	284
rect	261	286	262	287
rect	261	289	262	290
rect	261	301	262	302
rect	261	304	262	305
rect	261	307	262	308
rect	261	310	262	311
rect	261	316	262	317
rect	261	319	262	320
rect	261	322	262	323
rect	261	325	262	326
rect	261	328	262	329
rect	261	334	262	335
rect	261	337	262	338
rect	261	352	262	353
rect	261	355	262	356
rect	261	364	262	365
rect	262	7	263	8
rect	262	10	263	11
rect	262	13	263	14
rect	262	16	263	17
rect	262	19	263	20
rect	262	22	263	23
rect	262	28	263	29
rect	262	31	263	32
rect	262	34	263	35
rect	262	37	263	38
rect	262	40	263	41
rect	262	55	263	56
rect	262	64	263	65
rect	262	67	263	68
rect	262	70	263	71
rect	262	73	263	74
rect	262	76	263	77
rect	262	79	263	80
rect	262	82	263	83
rect	262	91	263	92
rect	262	94	263	95
rect	262	97	263	98
rect	262	100	263	101
rect	262	103	263	104
rect	262	106	263	107
rect	262	115	263	116
rect	262	118	263	119
rect	262	130	263	131
rect	262	133	263	134
rect	262	136	263	137
rect	262	139	263	140
rect	262	142	263	143
rect	262	148	263	149
rect	262	151	263	152
rect	262	154	263	155
rect	262	157	263	158
rect	262	166	263	167
rect	262	169	263	170
rect	262	172	263	173
rect	262	175	263	176
rect	262	178	263	179
rect	262	181	263	182
rect	262	190	263	191
rect	262	193	263	194
rect	262	196	263	197
rect	262	205	263	206
rect	262	208	263	209
rect	262	217	263	218
rect	262	226	263	227
rect	262	229	263	230
rect	262	232	263	233
rect	262	238	263	239
rect	262	241	263	242
rect	262	244	263	245
rect	262	247	263	248
rect	262	253	263	254
rect	262	256	263	257
rect	262	259	263	260
rect	262	262	263	263
rect	262	271	263	272
rect	262	274	263	275
rect	262	277	263	278
rect	262	280	263	281
rect	262	283	263	284
rect	262	289	263	290
rect	262	301	263	302
rect	262	304	263	305
rect	262	307	263	308
rect	262	310	263	311
rect	262	316	263	317
rect	262	319	263	320
rect	262	322	263	323
rect	262	325	263	326
rect	262	328	263	329
rect	262	334	263	335
rect	262	337	263	338
rect	262	352	263	353
rect	262	355	263	356
rect	262	364	263	365
rect	263	7	264	8
rect	263	10	264	11
rect	263	13	264	14
rect	263	16	264	17
rect	263	19	264	20
rect	263	22	264	23
rect	263	28	264	29
rect	263	31	264	32
rect	263	34	264	35
rect	263	37	264	38
rect	263	40	264	41
rect	263	55	264	56
rect	263	64	264	65
rect	263	67	264	68
rect	263	70	264	71
rect	263	73	264	74
rect	263	76	264	77
rect	263	79	264	80
rect	263	82	264	83
rect	263	91	264	92
rect	263	94	264	95
rect	263	97	264	98
rect	263	100	264	101
rect	263	103	264	104
rect	263	106	264	107
rect	263	115	264	116
rect	263	118	264	119
rect	263	130	264	131
rect	263	133	264	134
rect	263	136	264	137
rect	263	139	264	140
rect	263	142	264	143
rect	263	148	264	149
rect	263	151	264	152
rect	263	154	264	155
rect	263	157	264	158
rect	263	166	264	167
rect	263	169	264	170
rect	263	172	264	173
rect	263	175	264	176
rect	263	178	264	179
rect	263	181	264	182
rect	263	190	264	191
rect	263	193	264	194
rect	263	196	264	197
rect	263	205	264	206
rect	263	208	264	209
rect	263	217	264	218
rect	263	226	264	227
rect	263	229	264	230
rect	263	232	264	233
rect	263	238	264	239
rect	263	241	264	242
rect	263	244	264	245
rect	263	247	264	248
rect	263	253	264	254
rect	263	256	264	257
rect	263	259	264	260
rect	263	262	264	263
rect	263	271	264	272
rect	263	274	264	275
rect	263	277	264	278
rect	263	280	264	281
rect	263	283	264	284
rect	263	289	264	290
rect	263	298	264	299
rect	263	301	264	302
rect	263	304	264	305
rect	263	307	264	308
rect	263	310	264	311
rect	263	316	264	317
rect	263	319	264	320
rect	263	322	264	323
rect	263	325	264	326
rect	263	328	264	329
rect	263	334	264	335
rect	263	337	264	338
rect	263	352	264	353
rect	263	355	264	356
rect	263	364	264	365
rect	264	7	265	8
rect	264	10	265	11
rect	264	13	265	14
rect	264	16	265	17
rect	264	19	265	20
rect	264	22	265	23
rect	264	28	265	29
rect	264	31	265	32
rect	264	34	265	35
rect	264	37	265	38
rect	264	40	265	41
rect	264	55	265	56
rect	264	64	265	65
rect	264	67	265	68
rect	264	70	265	71
rect	264	73	265	74
rect	264	76	265	77
rect	264	79	265	80
rect	264	82	265	83
rect	264	91	265	92
rect	264	94	265	95
rect	264	97	265	98
rect	264	100	265	101
rect	264	103	265	104
rect	264	106	265	107
rect	264	115	265	116
rect	264	118	265	119
rect	264	130	265	131
rect	264	133	265	134
rect	264	136	265	137
rect	264	139	265	140
rect	264	142	265	143
rect	264	148	265	149
rect	264	151	265	152
rect	264	154	265	155
rect	264	157	265	158
rect	264	166	265	167
rect	264	169	265	170
rect	264	172	265	173
rect	264	175	265	176
rect	264	178	265	179
rect	264	181	265	182
rect	264	190	265	191
rect	264	193	265	194
rect	264	196	265	197
rect	264	205	265	206
rect	264	208	265	209
rect	264	217	265	218
rect	264	226	265	227
rect	264	229	265	230
rect	264	232	265	233
rect	264	238	265	239
rect	264	241	265	242
rect	264	244	265	245
rect	264	247	265	248
rect	264	253	265	254
rect	264	256	265	257
rect	264	259	265	260
rect	264	262	265	263
rect	264	271	265	272
rect	264	274	265	275
rect	264	277	265	278
rect	264	283	265	284
rect	264	289	265	290
rect	264	298	265	299
rect	264	301	265	302
rect	264	304	265	305
rect	264	307	265	308
rect	264	310	265	311
rect	264	316	265	317
rect	264	319	265	320
rect	264	322	265	323
rect	264	325	265	326
rect	264	328	265	329
rect	264	334	265	335
rect	264	337	265	338
rect	264	352	265	353
rect	264	355	265	356
rect	264	364	265	365
rect	265	7	266	8
rect	265	10	266	11
rect	265	13	266	14
rect	265	16	266	17
rect	265	19	266	20
rect	265	22	266	23
rect	265	28	266	29
rect	265	31	266	32
rect	265	34	266	35
rect	265	37	266	38
rect	265	40	266	41
rect	265	55	266	56
rect	265	64	266	65
rect	265	67	266	68
rect	265	70	266	71
rect	265	73	266	74
rect	265	76	266	77
rect	265	79	266	80
rect	265	82	266	83
rect	265	91	266	92
rect	265	94	266	95
rect	265	97	266	98
rect	265	100	266	101
rect	265	103	266	104
rect	265	106	266	107
rect	265	115	266	116
rect	265	118	266	119
rect	265	130	266	131
rect	265	133	266	134
rect	265	136	266	137
rect	265	139	266	140
rect	265	142	266	143
rect	265	148	266	149
rect	265	151	266	152
rect	265	154	266	155
rect	265	157	266	158
rect	265	166	266	167
rect	265	169	266	170
rect	265	172	266	173
rect	265	175	266	176
rect	265	178	266	179
rect	265	181	266	182
rect	265	190	266	191
rect	265	193	266	194
rect	265	196	266	197
rect	265	205	266	206
rect	265	208	266	209
rect	265	217	266	218
rect	265	226	266	227
rect	265	229	266	230
rect	265	232	266	233
rect	265	238	266	239
rect	265	241	266	242
rect	265	244	266	245
rect	265	247	266	248
rect	265	253	266	254
rect	265	256	266	257
rect	265	259	266	260
rect	265	262	266	263
rect	265	271	266	272
rect	265	274	266	275
rect	265	277	266	278
rect	265	283	266	284
rect	265	286	266	287
rect	265	289	266	290
rect	265	298	266	299
rect	265	301	266	302
rect	265	304	266	305
rect	265	307	266	308
rect	265	310	266	311
rect	265	316	266	317
rect	265	319	266	320
rect	265	322	266	323
rect	265	325	266	326
rect	265	328	266	329
rect	265	334	266	335
rect	265	337	266	338
rect	265	352	266	353
rect	265	355	266	356
rect	265	364	266	365
rect	266	7	267	8
rect	266	10	267	11
rect	266	13	267	14
rect	266	16	267	17
rect	266	19	267	20
rect	266	22	267	23
rect	266	28	267	29
rect	266	31	267	32
rect	266	34	267	35
rect	266	37	267	38
rect	266	40	267	41
rect	266	55	267	56
rect	266	64	267	65
rect	266	67	267	68
rect	266	70	267	71
rect	266	73	267	74
rect	266	76	267	77
rect	266	79	267	80
rect	266	82	267	83
rect	266	91	267	92
rect	266	94	267	95
rect	266	97	267	98
rect	266	100	267	101
rect	266	103	267	104
rect	266	106	267	107
rect	266	115	267	116
rect	266	118	267	119
rect	266	130	267	131
rect	266	133	267	134
rect	266	136	267	137
rect	266	139	267	140
rect	266	142	267	143
rect	266	148	267	149
rect	266	151	267	152
rect	266	154	267	155
rect	266	157	267	158
rect	266	166	267	167
rect	266	169	267	170
rect	266	172	267	173
rect	266	175	267	176
rect	266	178	267	179
rect	266	181	267	182
rect	266	190	267	191
rect	266	193	267	194
rect	266	196	267	197
rect	266	205	267	206
rect	266	208	267	209
rect	266	217	267	218
rect	266	229	267	230
rect	266	232	267	233
rect	266	238	267	239
rect	266	241	267	242
rect	266	244	267	245
rect	266	247	267	248
rect	266	253	267	254
rect	266	256	267	257
rect	266	259	267	260
rect	266	262	267	263
rect	266	271	267	272
rect	266	274	267	275
rect	266	277	267	278
rect	266	283	267	284
rect	266	286	267	287
rect	266	289	267	290
rect	266	298	267	299
rect	266	301	267	302
rect	266	304	267	305
rect	266	307	267	308
rect	266	310	267	311
rect	266	316	267	317
rect	266	319	267	320
rect	266	322	267	323
rect	266	325	267	326
rect	266	328	267	329
rect	266	334	267	335
rect	266	337	267	338
rect	266	352	267	353
rect	266	355	267	356
rect	266	364	267	365
rect	267	7	268	8
rect	267	10	268	11
rect	267	13	268	14
rect	267	16	268	17
rect	267	19	268	20
rect	267	22	268	23
rect	267	28	268	29
rect	267	31	268	32
rect	267	34	268	35
rect	267	37	268	38
rect	267	40	268	41
rect	267	55	268	56
rect	267	64	268	65
rect	267	67	268	68
rect	267	70	268	71
rect	267	73	268	74
rect	267	76	268	77
rect	267	79	268	80
rect	267	82	268	83
rect	267	91	268	92
rect	267	94	268	95
rect	267	97	268	98
rect	267	100	268	101
rect	267	103	268	104
rect	267	106	268	107
rect	267	115	268	116
rect	267	118	268	119
rect	267	130	268	131
rect	267	133	268	134
rect	267	136	268	137
rect	267	139	268	140
rect	267	142	268	143
rect	267	148	268	149
rect	267	151	268	152
rect	267	154	268	155
rect	267	157	268	158
rect	267	166	268	167
rect	267	169	268	170
rect	267	172	268	173
rect	267	175	268	176
rect	267	178	268	179
rect	267	181	268	182
rect	267	190	268	191
rect	267	193	268	194
rect	267	196	268	197
rect	267	205	268	206
rect	267	208	268	209
rect	267	217	268	218
rect	267	229	268	230
rect	267	232	268	233
rect	267	238	268	239
rect	267	241	268	242
rect	267	244	268	245
rect	267	247	268	248
rect	267	253	268	254
rect	267	256	268	257
rect	267	259	268	260
rect	267	262	268	263
rect	267	271	268	272
rect	267	274	268	275
rect	267	277	268	278
rect	267	280	268	281
rect	267	283	268	284
rect	267	286	268	287
rect	267	289	268	290
rect	267	298	268	299
rect	267	301	268	302
rect	267	304	268	305
rect	267	307	268	308
rect	267	310	268	311
rect	267	316	268	317
rect	267	319	268	320
rect	267	322	268	323
rect	267	325	268	326
rect	267	328	268	329
rect	267	334	268	335
rect	267	337	268	338
rect	267	352	268	353
rect	267	355	268	356
rect	267	364	268	365
rect	268	7	269	8
rect	268	10	269	11
rect	268	13	269	14
rect	268	16	269	17
rect	268	19	269	20
rect	268	22	269	23
rect	268	28	269	29
rect	268	31	269	32
rect	268	34	269	35
rect	268	37	269	38
rect	268	40	269	41
rect	268	55	269	56
rect	268	64	269	65
rect	268	67	269	68
rect	268	70	269	71
rect	268	73	269	74
rect	268	76	269	77
rect	268	79	269	80
rect	268	82	269	83
rect	268	91	269	92
rect	268	94	269	95
rect	268	97	269	98
rect	268	100	269	101
rect	268	103	269	104
rect	268	106	269	107
rect	268	115	269	116
rect	268	118	269	119
rect	268	130	269	131
rect	268	133	269	134
rect	268	136	269	137
rect	268	139	269	140
rect	268	142	269	143
rect	268	148	269	149
rect	268	151	269	152
rect	268	154	269	155
rect	268	157	269	158
rect	268	166	269	167
rect	268	169	269	170
rect	268	172	269	173
rect	268	175	269	176
rect	268	178	269	179
rect	268	181	269	182
rect	268	190	269	191
rect	268	193	269	194
rect	268	196	269	197
rect	268	205	269	206
rect	268	208	269	209
rect	268	229	269	230
rect	268	232	269	233
rect	268	238	269	239
rect	268	241	269	242
rect	268	244	269	245
rect	268	247	269	248
rect	268	253	269	254
rect	268	256	269	257
rect	268	259	269	260
rect	268	262	269	263
rect	268	271	269	272
rect	268	274	269	275
rect	268	277	269	278
rect	268	280	269	281
rect	268	283	269	284
rect	268	286	269	287
rect	268	289	269	290
rect	268	298	269	299
rect	268	301	269	302
rect	268	304	269	305
rect	268	307	269	308
rect	268	310	269	311
rect	268	316	269	317
rect	268	319	269	320
rect	268	322	269	323
rect	268	325	269	326
rect	268	328	269	329
rect	268	334	269	335
rect	268	337	269	338
rect	268	352	269	353
rect	268	355	269	356
rect	268	364	269	365
rect	269	7	270	8
rect	269	10	270	11
rect	269	13	270	14
rect	269	16	270	17
rect	269	19	270	20
rect	269	22	270	23
rect	269	28	270	29
rect	269	31	270	32
rect	269	34	270	35
rect	269	37	270	38
rect	269	40	270	41
rect	269	55	270	56
rect	269	64	270	65
rect	269	67	270	68
rect	269	70	270	71
rect	269	73	270	74
rect	269	76	270	77
rect	269	79	270	80
rect	269	82	270	83
rect	269	91	270	92
rect	269	94	270	95
rect	269	97	270	98
rect	269	100	270	101
rect	269	103	270	104
rect	269	106	270	107
rect	269	115	270	116
rect	269	118	270	119
rect	269	130	270	131
rect	269	133	270	134
rect	269	136	270	137
rect	269	139	270	140
rect	269	142	270	143
rect	269	148	270	149
rect	269	151	270	152
rect	269	154	270	155
rect	269	157	270	158
rect	269	166	270	167
rect	269	169	270	170
rect	269	172	270	173
rect	269	175	270	176
rect	269	178	270	179
rect	269	181	270	182
rect	269	190	270	191
rect	269	193	270	194
rect	269	196	270	197
rect	269	205	270	206
rect	269	208	270	209
rect	269	226	270	227
rect	269	229	270	230
rect	269	232	270	233
rect	269	238	270	239
rect	269	241	270	242
rect	269	244	270	245
rect	269	247	270	248
rect	269	253	270	254
rect	269	256	270	257
rect	269	259	270	260
rect	269	262	270	263
rect	269	271	270	272
rect	269	274	270	275
rect	269	277	270	278
rect	269	280	270	281
rect	269	283	270	284
rect	269	286	270	287
rect	269	289	270	290
rect	269	298	270	299
rect	269	301	270	302
rect	269	304	270	305
rect	269	307	270	308
rect	269	310	270	311
rect	269	316	270	317
rect	269	319	270	320
rect	269	322	270	323
rect	269	325	270	326
rect	269	328	270	329
rect	269	334	270	335
rect	269	337	270	338
rect	269	352	270	353
rect	269	355	270	356
rect	269	364	270	365
rect	270	7	271	8
rect	270	10	271	11
rect	270	13	271	14
rect	270	16	271	17
rect	270	19	271	20
rect	270	22	271	23
rect	270	28	271	29
rect	270	31	271	32
rect	270	34	271	35
rect	270	37	271	38
rect	270	40	271	41
rect	270	55	271	56
rect	270	64	271	65
rect	270	67	271	68
rect	270	70	271	71
rect	270	73	271	74
rect	270	76	271	77
rect	270	79	271	80
rect	270	82	271	83
rect	270	91	271	92
rect	270	94	271	95
rect	270	97	271	98
rect	270	100	271	101
rect	270	103	271	104
rect	270	106	271	107
rect	270	115	271	116
rect	270	118	271	119
rect	270	130	271	131
rect	270	133	271	134
rect	270	136	271	137
rect	270	139	271	140
rect	270	142	271	143
rect	270	148	271	149
rect	270	151	271	152
rect	270	154	271	155
rect	270	157	271	158
rect	270	166	271	167
rect	270	169	271	170
rect	270	172	271	173
rect	270	175	271	176
rect	270	178	271	179
rect	270	181	271	182
rect	270	190	271	191
rect	270	196	271	197
rect	270	205	271	206
rect	270	208	271	209
rect	270	226	271	227
rect	270	229	271	230
rect	270	232	271	233
rect	270	238	271	239
rect	270	241	271	242
rect	270	244	271	245
rect	270	247	271	248
rect	270	253	271	254
rect	270	256	271	257
rect	270	259	271	260
rect	270	262	271	263
rect	270	271	271	272
rect	270	274	271	275
rect	270	277	271	278
rect	270	280	271	281
rect	270	283	271	284
rect	270	286	271	287
rect	270	289	271	290
rect	270	298	271	299
rect	270	301	271	302
rect	270	304	271	305
rect	270	307	271	308
rect	270	310	271	311
rect	270	316	271	317
rect	270	319	271	320
rect	270	322	271	323
rect	270	325	271	326
rect	270	328	271	329
rect	270	334	271	335
rect	270	337	271	338
rect	270	352	271	353
rect	270	355	271	356
rect	270	364	271	365
rect	271	7	272	8
rect	271	10	272	11
rect	271	13	272	14
rect	271	16	272	17
rect	271	19	272	20
rect	271	22	272	23
rect	271	28	272	29
rect	271	31	272	32
rect	271	34	272	35
rect	271	37	272	38
rect	271	40	272	41
rect	271	55	272	56
rect	271	64	272	65
rect	271	67	272	68
rect	271	70	272	71
rect	271	73	272	74
rect	271	76	272	77
rect	271	79	272	80
rect	271	82	272	83
rect	271	91	272	92
rect	271	94	272	95
rect	271	97	272	98
rect	271	100	272	101
rect	271	103	272	104
rect	271	106	272	107
rect	271	115	272	116
rect	271	118	272	119
rect	271	130	272	131
rect	271	133	272	134
rect	271	136	272	137
rect	271	139	272	140
rect	271	142	272	143
rect	271	148	272	149
rect	271	151	272	152
rect	271	154	272	155
rect	271	157	272	158
rect	271	166	272	167
rect	271	169	272	170
rect	271	172	272	173
rect	271	175	272	176
rect	271	178	272	179
rect	271	181	272	182
rect	271	190	272	191
rect	271	196	272	197
rect	271	205	272	206
rect	271	208	272	209
rect	271	217	272	218
rect	271	226	272	227
rect	271	229	272	230
rect	271	232	272	233
rect	271	238	272	239
rect	271	241	272	242
rect	271	244	272	245
rect	271	247	272	248
rect	271	253	272	254
rect	271	256	272	257
rect	271	259	272	260
rect	271	262	272	263
rect	271	271	272	272
rect	271	274	272	275
rect	271	277	272	278
rect	271	280	272	281
rect	271	283	272	284
rect	271	286	272	287
rect	271	289	272	290
rect	271	298	272	299
rect	271	301	272	302
rect	271	304	272	305
rect	271	307	272	308
rect	271	310	272	311
rect	271	316	272	317
rect	271	319	272	320
rect	271	322	272	323
rect	271	325	272	326
rect	271	328	272	329
rect	271	334	272	335
rect	271	337	272	338
rect	271	352	272	353
rect	271	355	272	356
rect	271	364	272	365
rect	272	7	273	8
rect	272	10	273	11
rect	272	13	273	14
rect	272	16	273	17
rect	272	19	273	20
rect	272	22	273	23
rect	272	28	273	29
rect	272	31	273	32
rect	272	34	273	35
rect	272	37	273	38
rect	272	40	273	41
rect	272	55	273	56
rect	272	64	273	65
rect	272	67	273	68
rect	272	70	273	71
rect	272	73	273	74
rect	272	76	273	77
rect	272	79	273	80
rect	272	82	273	83
rect	272	91	273	92
rect	272	94	273	95
rect	272	97	273	98
rect	272	100	273	101
rect	272	103	273	104
rect	272	106	273	107
rect	272	115	273	116
rect	272	118	273	119
rect	272	130	273	131
rect	272	133	273	134
rect	272	136	273	137
rect	272	139	273	140
rect	272	142	273	143
rect	272	148	273	149
rect	272	151	273	152
rect	272	154	273	155
rect	272	157	273	158
rect	272	166	273	167
rect	272	169	273	170
rect	272	172	273	173
rect	272	178	273	179
rect	272	181	273	182
rect	272	190	273	191
rect	272	196	273	197
rect	272	205	273	206
rect	272	208	273	209
rect	272	217	273	218
rect	272	226	273	227
rect	272	229	273	230
rect	272	232	273	233
rect	272	238	273	239
rect	272	241	273	242
rect	272	244	273	245
rect	272	247	273	248
rect	272	253	273	254
rect	272	256	273	257
rect	272	259	273	260
rect	272	262	273	263
rect	272	271	273	272
rect	272	274	273	275
rect	272	277	273	278
rect	272	280	273	281
rect	272	283	273	284
rect	272	286	273	287
rect	272	289	273	290
rect	272	298	273	299
rect	272	301	273	302
rect	272	304	273	305
rect	272	307	273	308
rect	272	310	273	311
rect	272	316	273	317
rect	272	319	273	320
rect	272	322	273	323
rect	272	325	273	326
rect	272	328	273	329
rect	272	334	273	335
rect	272	337	273	338
rect	272	352	273	353
rect	272	355	273	356
rect	272	364	273	365
rect	273	7	274	8
rect	273	10	274	11
rect	273	13	274	14
rect	273	16	274	17
rect	273	19	274	20
rect	273	22	274	23
rect	273	28	274	29
rect	273	31	274	32
rect	273	34	274	35
rect	273	37	274	38
rect	273	40	274	41
rect	273	55	274	56
rect	273	64	274	65
rect	273	67	274	68
rect	273	70	274	71
rect	273	73	274	74
rect	273	76	274	77
rect	273	79	274	80
rect	273	82	274	83
rect	273	91	274	92
rect	273	94	274	95
rect	273	97	274	98
rect	273	100	274	101
rect	273	103	274	104
rect	273	106	274	107
rect	273	115	274	116
rect	273	118	274	119
rect	273	130	274	131
rect	273	133	274	134
rect	273	136	274	137
rect	273	139	274	140
rect	273	142	274	143
rect	273	148	274	149
rect	273	151	274	152
rect	273	154	274	155
rect	273	157	274	158
rect	273	166	274	167
rect	273	169	274	170
rect	273	172	274	173
rect	273	178	274	179
rect	273	181	274	182
rect	273	190	274	191
rect	273	193	274	194
rect	273	196	274	197
rect	273	205	274	206
rect	273	208	274	209
rect	273	217	274	218
rect	273	226	274	227
rect	273	229	274	230
rect	273	232	274	233
rect	273	238	274	239
rect	273	241	274	242
rect	273	244	274	245
rect	273	247	274	248
rect	273	253	274	254
rect	273	256	274	257
rect	273	259	274	260
rect	273	262	274	263
rect	273	271	274	272
rect	273	274	274	275
rect	273	277	274	278
rect	273	280	274	281
rect	273	283	274	284
rect	273	286	274	287
rect	273	289	274	290
rect	273	298	274	299
rect	273	301	274	302
rect	273	304	274	305
rect	273	307	274	308
rect	273	310	274	311
rect	273	316	274	317
rect	273	319	274	320
rect	273	322	274	323
rect	273	325	274	326
rect	273	328	274	329
rect	273	334	274	335
rect	273	337	274	338
rect	273	352	274	353
rect	273	355	274	356
rect	273	364	274	365
rect	274	7	275	8
rect	274	10	275	11
rect	274	13	275	14
rect	274	16	275	17
rect	274	19	275	20
rect	274	22	275	23
rect	274	28	275	29
rect	274	31	275	32
rect	274	34	275	35
rect	274	37	275	38
rect	274	40	275	41
rect	274	55	275	56
rect	274	64	275	65
rect	274	67	275	68
rect	274	70	275	71
rect	274	73	275	74
rect	274	76	275	77
rect	274	79	275	80
rect	274	91	275	92
rect	274	94	275	95
rect	274	97	275	98
rect	274	100	275	101
rect	274	103	275	104
rect	274	106	275	107
rect	274	115	275	116
rect	274	118	275	119
rect	274	130	275	131
rect	274	133	275	134
rect	274	136	275	137
rect	274	139	275	140
rect	274	142	275	143
rect	274	148	275	149
rect	274	151	275	152
rect	274	154	275	155
rect	274	157	275	158
rect	274	166	275	167
rect	274	169	275	170
rect	274	178	275	179
rect	274	181	275	182
rect	274	190	275	191
rect	274	193	275	194
rect	274	196	275	197
rect	274	205	275	206
rect	274	208	275	209
rect	274	217	275	218
rect	274	226	275	227
rect	274	229	275	230
rect	274	232	275	233
rect	274	238	275	239
rect	274	241	275	242
rect	274	244	275	245
rect	274	247	275	248
rect	274	253	275	254
rect	274	256	275	257
rect	274	259	275	260
rect	274	262	275	263
rect	274	271	275	272
rect	274	274	275	275
rect	274	277	275	278
rect	274	280	275	281
rect	274	283	275	284
rect	274	286	275	287
rect	274	289	275	290
rect	274	298	275	299
rect	274	301	275	302
rect	274	304	275	305
rect	274	307	275	308
rect	274	310	275	311
rect	274	316	275	317
rect	274	319	275	320
rect	274	322	275	323
rect	274	325	275	326
rect	274	328	275	329
rect	274	334	275	335
rect	274	337	275	338
rect	274	352	275	353
rect	274	355	275	356
rect	274	364	275	365
rect	275	7	276	8
rect	275	10	276	11
rect	275	13	276	14
rect	275	16	276	17
rect	275	19	276	20
rect	275	22	276	23
rect	275	28	276	29
rect	275	31	276	32
rect	275	34	276	35
rect	275	37	276	38
rect	275	40	276	41
rect	275	55	276	56
rect	275	58	276	59
rect	275	64	276	65
rect	275	67	276	68
rect	275	70	276	71
rect	275	73	276	74
rect	275	76	276	77
rect	275	79	276	80
rect	275	91	276	92
rect	275	94	276	95
rect	275	97	276	98
rect	275	100	276	101
rect	275	103	276	104
rect	275	106	276	107
rect	275	115	276	116
rect	275	118	276	119
rect	275	130	276	131
rect	275	133	276	134
rect	275	136	276	137
rect	275	139	276	140
rect	275	142	276	143
rect	275	148	276	149
rect	275	151	276	152
rect	275	154	276	155
rect	275	157	276	158
rect	275	166	276	167
rect	275	169	276	170
rect	275	178	276	179
rect	275	181	276	182
rect	275	187	276	188
rect	275	190	276	191
rect	275	193	276	194
rect	275	196	276	197
rect	275	205	276	206
rect	275	208	276	209
rect	275	217	276	218
rect	275	226	276	227
rect	275	229	276	230
rect	275	232	276	233
rect	275	238	276	239
rect	275	241	276	242
rect	275	244	276	245
rect	275	247	276	248
rect	275	253	276	254
rect	275	256	276	257
rect	275	259	276	260
rect	275	262	276	263
rect	275	271	276	272
rect	275	274	276	275
rect	275	277	276	278
rect	275	280	276	281
rect	275	283	276	284
rect	275	286	276	287
rect	275	289	276	290
rect	275	298	276	299
rect	275	301	276	302
rect	275	304	276	305
rect	275	307	276	308
rect	275	310	276	311
rect	275	316	276	317
rect	275	319	276	320
rect	275	322	276	323
rect	275	325	276	326
rect	275	328	276	329
rect	275	334	276	335
rect	275	337	276	338
rect	275	352	276	353
rect	275	355	276	356
rect	275	364	276	365
rect	276	7	277	8
rect	276	10	277	11
rect	276	13	277	14
rect	276	16	277	17
rect	276	19	277	20
rect	276	22	277	23
rect	276	28	277	29
rect	276	31	277	32
rect	276	34	277	35
rect	276	37	277	38
rect	276	40	277	41
rect	276	55	277	56
rect	276	58	277	59
rect	276	64	277	65
rect	276	67	277	68
rect	276	70	277	71
rect	276	73	277	74
rect	276	76	277	77
rect	276	91	277	92
rect	276	94	277	95
rect	276	97	277	98
rect	276	100	277	101
rect	276	103	277	104
rect	276	106	277	107
rect	276	115	277	116
rect	276	118	277	119
rect	276	130	277	131
rect	276	133	277	134
rect	276	136	277	137
rect	276	139	277	140
rect	276	142	277	143
rect	276	148	277	149
rect	276	154	277	155
rect	276	157	277	158
rect	276	166	277	167
rect	276	169	277	170
rect	276	178	277	179
rect	276	181	277	182
rect	276	187	277	188
rect	276	190	277	191
rect	276	193	277	194
rect	276	196	277	197
rect	276	205	277	206
rect	276	208	277	209
rect	276	217	277	218
rect	276	226	277	227
rect	276	229	277	230
rect	276	232	277	233
rect	276	238	277	239
rect	276	241	277	242
rect	276	244	277	245
rect	276	247	277	248
rect	276	253	277	254
rect	276	256	277	257
rect	276	259	277	260
rect	276	262	277	263
rect	276	271	277	272
rect	276	274	277	275
rect	276	277	277	278
rect	276	280	277	281
rect	276	283	277	284
rect	276	286	277	287
rect	276	289	277	290
rect	276	298	277	299
rect	276	301	277	302
rect	276	304	277	305
rect	276	307	277	308
rect	276	310	277	311
rect	276	316	277	317
rect	276	319	277	320
rect	276	322	277	323
rect	276	325	277	326
rect	276	328	277	329
rect	276	334	277	335
rect	276	337	277	338
rect	276	352	277	353
rect	276	355	277	356
rect	276	364	277	365
rect	277	7	278	8
rect	277	10	278	11
rect	277	13	278	14
rect	277	16	278	17
rect	277	19	278	20
rect	277	22	278	23
rect	277	28	278	29
rect	277	31	278	32
rect	277	34	278	35
rect	277	37	278	38
rect	277	40	278	41
rect	277	55	278	56
rect	277	58	278	59
rect	277	64	278	65
rect	277	67	278	68
rect	277	70	278	71
rect	277	73	278	74
rect	277	76	278	77
rect	277	82	278	83
rect	277	91	278	92
rect	277	94	278	95
rect	277	97	278	98
rect	277	100	278	101
rect	277	103	278	104
rect	277	106	278	107
rect	277	115	278	116
rect	277	118	278	119
rect	277	130	278	131
rect	277	133	278	134
rect	277	136	278	137
rect	277	139	278	140
rect	277	142	278	143
rect	277	148	278	149
rect	277	154	278	155
rect	277	157	278	158
rect	277	166	278	167
rect	277	169	278	170
rect	277	178	278	179
rect	277	181	278	182
rect	277	184	278	185
rect	277	187	278	188
rect	277	190	278	191
rect	277	193	278	194
rect	277	196	278	197
rect	277	205	278	206
rect	277	208	278	209
rect	277	217	278	218
rect	277	226	278	227
rect	277	229	278	230
rect	277	232	278	233
rect	277	238	278	239
rect	277	241	278	242
rect	277	244	278	245
rect	277	247	278	248
rect	277	253	278	254
rect	277	256	278	257
rect	277	259	278	260
rect	277	262	278	263
rect	277	271	278	272
rect	277	274	278	275
rect	277	277	278	278
rect	277	280	278	281
rect	277	283	278	284
rect	277	286	278	287
rect	277	289	278	290
rect	277	298	278	299
rect	277	301	278	302
rect	277	304	278	305
rect	277	307	278	308
rect	277	310	278	311
rect	277	316	278	317
rect	277	319	278	320
rect	277	322	278	323
rect	277	325	278	326
rect	277	328	278	329
rect	277	334	278	335
rect	277	337	278	338
rect	277	352	278	353
rect	277	355	278	356
rect	277	364	278	365
rect	278	7	279	8
rect	278	10	279	11
rect	278	13	279	14
rect	278	16	279	17
rect	278	19	279	20
rect	278	22	279	23
rect	278	31	279	32
rect	278	34	279	35
rect	278	40	279	41
rect	278	55	279	56
rect	278	58	279	59
rect	278	64	279	65
rect	278	67	279	68
rect	278	70	279	71
rect	278	73	279	74
rect	278	82	279	83
rect	278	91	279	92
rect	278	94	279	95
rect	278	97	279	98
rect	278	100	279	101
rect	278	103	279	104
rect	278	106	279	107
rect	278	115	279	116
rect	278	118	279	119
rect	278	130	279	131
rect	278	133	279	134
rect	278	139	279	140
rect	278	142	279	143
rect	278	148	279	149
rect	278	154	279	155
rect	278	157	279	158
rect	278	166	279	167
rect	278	178	279	179
rect	278	181	279	182
rect	278	184	279	185
rect	278	187	279	188
rect	278	190	279	191
rect	278	193	279	194
rect	278	196	279	197
rect	278	205	279	206
rect	278	208	279	209
rect	278	217	279	218
rect	278	226	279	227
rect	278	229	279	230
rect	278	232	279	233
rect	278	238	279	239
rect	278	241	279	242
rect	278	244	279	245
rect	278	247	279	248
rect	278	253	279	254
rect	278	256	279	257
rect	278	259	279	260
rect	278	271	279	272
rect	278	274	279	275
rect	278	277	279	278
rect	278	280	279	281
rect	278	283	279	284
rect	278	286	279	287
rect	278	298	279	299
rect	278	301	279	302
rect	278	304	279	305
rect	278	307	279	308
rect	278	319	279	320
rect	278	322	279	323
rect	278	325	279	326
rect	278	328	279	329
rect	278	334	279	335
rect	278	337	279	338
rect	278	352	279	353
rect	278	355	279	356
rect	278	364	279	365
rect	279	7	280	8
rect	279	10	280	11
rect	279	13	280	14
rect	279	16	280	17
rect	279	19	280	20
rect	279	22	280	23
rect	279	31	280	32
rect	279	34	280	35
rect	279	40	280	41
rect	279	55	280	56
rect	279	58	280	59
rect	279	64	280	65
rect	279	67	280	68
rect	279	70	280	71
rect	279	73	280	74
rect	279	82	280	83
rect	279	85	280	86
rect	279	91	280	92
rect	279	94	280	95
rect	279	97	280	98
rect	279	100	280	101
rect	279	103	280	104
rect	279	106	280	107
rect	279	115	280	116
rect	279	118	280	119
rect	279	130	280	131
rect	279	133	280	134
rect	279	139	280	140
rect	279	142	280	143
rect	279	148	280	149
rect	279	151	280	152
rect	279	154	280	155
rect	279	157	280	158
rect	279	166	280	167
rect	279	178	280	179
rect	279	181	280	182
rect	279	184	280	185
rect	279	187	280	188
rect	279	190	280	191
rect	279	193	280	194
rect	279	196	280	197
rect	279	205	280	206
rect	279	208	280	209
rect	279	211	280	212
rect	279	217	280	218
rect	279	226	280	227
rect	279	229	280	230
rect	279	232	280	233
rect	279	238	280	239
rect	279	241	280	242
rect	279	244	280	245
rect	279	247	280	248
rect	279	253	280	254
rect	279	256	280	257
rect	279	259	280	260
rect	279	268	280	269
rect	279	271	280	272
rect	279	274	280	275
rect	279	277	280	278
rect	279	280	280	281
rect	279	283	280	284
rect	279	286	280	287
rect	279	292	280	293
rect	279	298	280	299
rect	279	301	280	302
rect	279	304	280	305
rect	279	307	280	308
rect	279	319	280	320
rect	279	322	280	323
rect	279	325	280	326
rect	279	328	280	329
rect	279	334	280	335
rect	279	337	280	338
rect	279	352	280	353
rect	279	355	280	356
rect	279	364	280	365
rect	280	7	281	8
rect	280	10	281	11
rect	280	13	281	14
rect	280	16	281	17
rect	280	19	281	20
rect	280	22	281	23
rect	280	31	281	32
rect	280	40	281	41
rect	280	55	281	56
rect	280	58	281	59
rect	280	64	281	65
rect	280	67	281	68
rect	280	73	281	74
rect	280	82	281	83
rect	280	85	281	86
rect	280	91	281	92
rect	280	94	281	95
rect	280	97	281	98
rect	280	100	281	101
rect	280	103	281	104
rect	280	106	281	107
rect	280	115	281	116
rect	280	130	281	131
rect	280	133	281	134
rect	280	142	281	143
rect	280	148	281	149
rect	280	151	281	152
rect	280	157	281	158
rect	280	166	281	167
rect	280	181	281	182
rect	280	184	281	185
rect	280	187	281	188
rect	280	190	281	191
rect	280	193	281	194
rect	280	196	281	197
rect	280	205	281	206
rect	280	211	281	212
rect	280	217	281	218
rect	280	226	281	227
rect	280	229	281	230
rect	280	232	281	233
rect	280	238	281	239
rect	280	241	281	242
rect	280	244	281	245
rect	280	247	281	248
rect	280	253	281	254
rect	280	256	281	257
rect	280	268	281	269
rect	280	271	281	272
rect	280	274	281	275
rect	280	277	281	278
rect	280	280	281	281
rect	280	286	281	287
rect	280	292	281	293
rect	280	298	281	299
rect	280	301	281	302
rect	280	304	281	305
rect	280	319	281	320
rect	280	322	281	323
rect	280	325	281	326
rect	280	328	281	329
rect	280	334	281	335
rect	280	337	281	338
rect	280	352	281	353
rect	280	355	281	356
rect	280	364	281	365
rect	281	7	282	8
rect	281	10	282	11
rect	281	13	282	14
rect	281	16	282	17
rect	281	19	282	20
rect	281	22	282	23
rect	281	28	282	29
rect	281	31	282	32
rect	281	40	282	41
rect	281	55	282	56
rect	281	58	282	59
rect	281	64	282	65
rect	281	67	282	68
rect	281	73	282	74
rect	281	79	282	80
rect	281	82	282	83
rect	281	85	282	86
rect	281	91	282	92
rect	281	94	282	95
rect	281	97	282	98
rect	281	100	282	101
rect	281	103	282	104
rect	281	106	282	107
rect	281	115	282	116
rect	281	124	282	125
rect	281	130	282	131
rect	281	133	282	134
rect	281	136	282	137
rect	281	142	282	143
rect	281	148	282	149
rect	281	151	282	152
rect	281	157	282	158
rect	281	166	282	167
rect	281	172	282	173
rect	281	175	282	176
rect	281	181	282	182
rect	281	184	282	185
rect	281	187	282	188
rect	281	190	282	191
rect	281	193	282	194
rect	281	196	282	197
rect	281	199	282	200
rect	281	205	282	206
rect	281	211	282	212
rect	281	217	282	218
rect	281	226	282	227
rect	281	229	282	230
rect	281	232	282	233
rect	281	238	282	239
rect	281	241	282	242
rect	281	244	282	245
rect	281	247	282	248
rect	281	253	282	254
rect	281	256	282	257
rect	281	265	282	266
rect	281	268	282	269
rect	281	271	282	272
rect	281	274	282	275
rect	281	277	282	278
rect	281	280	282	281
rect	281	286	282	287
rect	281	289	282	290
rect	281	292	282	293
rect	281	298	282	299
rect	281	301	282	302
rect	281	304	282	305
rect	281	313	282	314
rect	281	319	282	320
rect	281	322	282	323
rect	281	325	282	326
rect	281	328	282	329
rect	281	334	282	335
rect	281	337	282	338
rect	281	352	282	353
rect	281	355	282	356
rect	281	364	282	365
rect	282	7	283	8
rect	282	10	283	11
rect	282	13	283	14
rect	282	19	283	20
rect	282	22	283	23
rect	282	28	283	29
rect	282	31	283	32
rect	282	40	283	41
rect	282	55	283	56
rect	282	58	283	59
rect	282	64	283	65
rect	282	79	283	80
rect	282	82	283	83
rect	282	85	283	86
rect	282	91	283	92
rect	282	94	283	95
rect	282	97	283	98
rect	282	100	283	101
rect	282	103	283	104
rect	282	106	283	107
rect	282	124	283	125
rect	282	130	283	131
rect	282	133	283	134
rect	282	136	283	137
rect	282	142	283	143
rect	282	148	283	149
rect	282	151	283	152
rect	282	157	283	158
rect	282	166	283	167
rect	282	172	283	173
rect	282	175	283	176
rect	282	181	283	182
rect	282	184	283	185
rect	282	187	283	188
rect	282	190	283	191
rect	282	193	283	194
rect	282	196	283	197
rect	282	199	283	200
rect	282	205	283	206
rect	282	211	283	212
rect	282	217	283	218
rect	282	226	283	227
rect	282	229	283	230
rect	282	232	283	233
rect	282	238	283	239
rect	282	241	283	242
rect	282	244	283	245
rect	282	247	283	248
rect	282	253	283	254
rect	282	256	283	257
rect	282	265	283	266
rect	282	268	283	269
rect	282	271	283	272
rect	282	274	283	275
rect	282	277	283	278
rect	282	280	283	281
rect	282	286	283	287
rect	282	289	283	290
rect	282	292	283	293
rect	282	298	283	299
rect	282	301	283	302
rect	282	304	283	305
rect	282	313	283	314
rect	282	319	283	320
rect	282	322	283	323
rect	282	325	283	326
rect	282	334	283	335
rect	282	337	283	338
rect	282	355	283	356
rect	282	364	283	365
rect	283	7	284	8
rect	283	10	284	11
rect	283	13	284	14
rect	283	19	284	20
rect	283	22	284	23
rect	283	28	284	29
rect	283	31	284	32
rect	283	34	284	35
rect	283	40	284	41
rect	283	55	284	56
rect	283	58	284	59
rect	283	64	284	65
rect	283	70	284	71
rect	283	76	284	77
rect	283	79	284	80
rect	283	82	284	83
rect	283	85	284	86
rect	283	91	284	92
rect	283	94	284	95
rect	283	97	284	98
rect	283	100	284	101
rect	283	103	284	104
rect	283	106	284	107
rect	283	118	284	119
rect	283	124	284	125
rect	283	130	284	131
rect	283	133	284	134
rect	283	136	284	137
rect	283	139	284	140
rect	283	142	284	143
rect	283	148	284	149
rect	283	151	284	152
rect	283	157	284	158
rect	283	166	284	167
rect	283	172	284	173
rect	283	175	284	176
rect	283	181	284	182
rect	283	184	284	185
rect	283	187	284	188
rect	283	190	284	191
rect	283	193	284	194
rect	283	196	284	197
rect	283	199	284	200
rect	283	205	284	206
rect	283	211	284	212
rect	283	217	284	218
rect	283	226	284	227
rect	283	229	284	230
rect	283	232	284	233
rect	283	238	284	239
rect	283	241	284	242
rect	283	244	284	245
rect	283	247	284	248
rect	283	253	284	254
rect	283	256	284	257
rect	283	265	284	266
rect	283	268	284	269
rect	283	271	284	272
rect	283	274	284	275
rect	283	277	284	278
rect	283	280	284	281
rect	283	286	284	287
rect	283	289	284	290
rect	283	292	284	293
rect	283	298	284	299
rect	283	301	284	302
rect	283	304	284	305
rect	283	313	284	314
rect	283	319	284	320
rect	283	322	284	323
rect	283	325	284	326
rect	283	334	284	335
rect	283	337	284	338
rect	283	355	284	356
rect	283	361	284	362
rect	283	364	284	365
rect	284	7	285	8
rect	284	13	285	14
rect	284	19	285	20
rect	284	28	285	29
rect	284	31	285	32
rect	284	34	285	35
rect	284	40	285	41
rect	284	55	285	56
rect	284	58	285	59
rect	284	64	285	65
rect	284	70	285	71
rect	284	76	285	77
rect	284	79	285	80
rect	284	82	285	83
rect	284	85	285	86
rect	284	91	285	92
rect	284	97	285	98
rect	284	100	285	101
rect	284	103	285	104
rect	284	106	285	107
rect	284	118	285	119
rect	284	124	285	125
rect	284	130	285	131
rect	284	136	285	137
rect	284	139	285	140
rect	284	142	285	143
rect	284	151	285	152
rect	284	172	285	173
rect	284	175	285	176
rect	284	181	285	182
rect	284	184	285	185
rect	284	187	285	188
rect	284	190	285	191
rect	284	193	285	194
rect	284	196	285	197
rect	284	199	285	200
rect	284	205	285	206
rect	284	211	285	212
rect	284	217	285	218
rect	284	226	285	227
rect	284	229	285	230
rect	284	232	285	233
rect	284	238	285	239
rect	284	244	285	245
rect	284	256	285	257
rect	284	265	285	266
rect	284	268	285	269
rect	284	271	285	272
rect	284	274	285	275
rect	284	277	285	278
rect	284	280	285	281
rect	284	286	285	287
rect	284	289	285	290
rect	284	292	285	293
rect	284	298	285	299
rect	284	301	285	302
rect	284	304	285	305
rect	284	313	285	314
rect	284	319	285	320
rect	284	322	285	323
rect	284	337	285	338
rect	284	361	285	362
rect	284	364	285	365
rect	285	7	286	8
rect	285	13	286	14
rect	285	16	286	17
rect	285	19	286	20
rect	285	28	286	29
rect	285	31	286	32
rect	285	34	286	35
rect	285	37	286	38
rect	285	40	286	41
rect	285	55	286	56
rect	285	58	286	59
rect	285	64	286	65
rect	285	67	286	68
rect	285	70	286	71
rect	285	76	286	77
rect	285	79	286	80
rect	285	82	286	83
rect	285	85	286	86
rect	285	88	286	89
rect	285	91	286	92
rect	285	97	286	98
rect	285	100	286	101
rect	285	103	286	104
rect	285	106	286	107
rect	285	118	286	119
rect	285	121	286	122
rect	285	124	286	125
rect	285	130	286	131
rect	285	136	286	137
rect	285	139	286	140
rect	285	142	286	143
rect	285	151	286	152
rect	285	154	286	155
rect	285	172	286	173
rect	285	175	286	176
rect	285	181	286	182
rect	285	184	286	185
rect	285	187	286	188
rect	285	190	286	191
rect	285	193	286	194
rect	285	196	286	197
rect	285	199	286	200
rect	285	205	286	206
rect	285	208	286	209
rect	285	211	286	212
rect	285	217	286	218
rect	285	226	286	227
rect	285	229	286	230
rect	285	232	286	233
rect	285	235	286	236
rect	285	238	286	239
rect	285	244	286	245
rect	285	250	286	251
rect	285	256	286	257
rect	285	265	286	266
rect	285	268	286	269
rect	285	271	286	272
rect	285	274	286	275
rect	285	277	286	278
rect	285	280	286	281
rect	285	286	286	287
rect	285	289	286	290
rect	285	292	286	293
rect	285	298	286	299
rect	285	301	286	302
rect	285	304	286	305
rect	285	313	286	314
rect	285	316	286	317
rect	285	319	286	320
rect	285	322	286	323
rect	285	331	286	332
rect	285	337	286	338
rect	285	349	286	350
rect	285	352	286	353
rect	285	361	286	362
rect	285	364	286	365
rect	286	7	287	8
rect	286	13	287	14
rect	286	16	287	17
rect	286	19	287	20
rect	286	28	287	29
rect	286	34	287	35
rect	286	37	287	38
rect	286	40	287	41
rect	286	55	287	56
rect	286	58	287	59
rect	286	67	287	68
rect	286	70	287	71
rect	286	76	287	77
rect	286	79	287	80
rect	286	82	287	83
rect	286	85	287	86
rect	286	88	287	89
rect	286	91	287	92
rect	286	97	287	98
rect	286	100	287	101
rect	286	103	287	104
rect	286	106	287	107
rect	286	118	287	119
rect	286	121	287	122
rect	286	124	287	125
rect	286	136	287	137
rect	286	139	287	140
rect	286	142	287	143
rect	286	151	287	152
rect	286	154	287	155
rect	286	172	287	173
rect	286	175	287	176
rect	286	184	287	185
rect	286	187	287	188
rect	286	190	287	191
rect	286	193	287	194
rect	286	196	287	197
rect	286	199	287	200
rect	286	205	287	206
rect	286	208	287	209
rect	286	211	287	212
rect	286	217	287	218
rect	286	226	287	227
rect	286	229	287	230
rect	286	235	287	236
rect	286	238	287	239
rect	286	244	287	245
rect	286	250	287	251
rect	286	256	287	257
rect	286	265	287	266
rect	286	268	287	269
rect	286	271	287	272
rect	286	274	287	275
rect	286	277	287	278
rect	286	280	287	281
rect	286	286	287	287
rect	286	289	287	290
rect	286	292	287	293
rect	286	298	287	299
rect	286	301	287	302
rect	286	304	287	305
rect	286	313	287	314
rect	286	316	287	317
rect	286	319	287	320
rect	286	322	287	323
rect	286	331	287	332
rect	286	337	287	338
rect	286	349	287	350
rect	286	352	287	353
rect	286	361	287	362
rect	286	364	287	365
rect	287	7	288	8
rect	287	10	288	11
rect	287	13	288	14
rect	287	16	288	17
rect	287	19	288	20
rect	287	28	288	29
rect	287	34	288	35
rect	287	37	288	38
rect	287	40	288	41
rect	287	55	288	56
rect	287	58	288	59
rect	287	67	288	68
rect	287	70	288	71
rect	287	76	288	77
rect	287	79	288	80
rect	287	82	288	83
rect	287	85	288	86
rect	287	88	288	89
rect	287	91	288	92
rect	287	97	288	98
rect	287	100	288	101
rect	287	103	288	104
rect	287	106	288	107
rect	287	115	288	116
rect	287	118	288	119
rect	287	121	288	122
rect	287	124	288	125
rect	287	136	288	137
rect	287	139	288	140
rect	287	142	288	143
rect	287	151	288	152
rect	287	154	288	155
rect	287	169	288	170
rect	287	172	288	173
rect	287	175	288	176
rect	287	178	288	179
rect	287	184	288	185
rect	287	187	288	188
rect	287	190	288	191
rect	287	193	288	194
rect	287	196	288	197
rect	287	199	288	200
rect	287	205	288	206
rect	287	208	288	209
rect	287	211	288	212
rect	287	217	288	218
rect	287	226	288	227
rect	287	229	288	230
rect	287	235	288	236
rect	287	238	288	239
rect	287	244	288	245
rect	287	250	288	251
rect	287	256	288	257
rect	287	265	288	266
rect	287	268	288	269
rect	287	271	288	272
rect	287	274	288	275
rect	287	277	288	278
rect	287	280	288	281
rect	287	286	288	287
rect	287	289	288	290
rect	287	292	288	293
rect	287	298	288	299
rect	287	301	288	302
rect	287	304	288	305
rect	287	313	288	314
rect	287	316	288	317
rect	287	319	288	320
rect	287	322	288	323
rect	287	331	288	332
rect	287	337	288	338
rect	287	349	288	350
rect	287	352	288	353
rect	287	355	288	356
rect	287	361	288	362
rect	287	364	288	365
rect	288	7	289	8
rect	288	10	289	11
rect	288	13	289	14
rect	288	16	289	17
rect	288	28	289	29
rect	288	34	289	35
rect	288	37	289	38
rect	288	40	289	41
rect	288	55	289	56
rect	288	58	289	59
rect	288	67	289	68
rect	288	70	289	71
rect	288	76	289	77
rect	288	79	289	80
rect	288	82	289	83
rect	288	85	289	86
rect	288	88	289	89
rect	288	91	289	92
rect	288	97	289	98
rect	288	100	289	101
rect	288	103	289	104
rect	288	106	289	107
rect	288	115	289	116
rect	288	118	289	119
rect	288	121	289	122
rect	288	124	289	125
rect	288	136	289	137
rect	288	139	289	140
rect	288	142	289	143
rect	288	151	289	152
rect	288	154	289	155
rect	288	169	289	170
rect	288	172	289	173
rect	288	175	289	176
rect	288	178	289	179
rect	288	184	289	185
rect	288	187	289	188
rect	288	190	289	191
rect	288	193	289	194
rect	288	196	289	197
rect	288	199	289	200
rect	288	205	289	206
rect	288	208	289	209
rect	288	211	289	212
rect	288	217	289	218
rect	288	226	289	227
rect	288	229	289	230
rect	288	235	289	236
rect	288	244	289	245
rect	288	250	289	251
rect	288	265	289	266
rect	288	268	289	269
rect	288	274	289	275
rect	288	277	289	278
rect	288	280	289	281
rect	288	286	289	287
rect	288	289	289	290
rect	288	292	289	293
rect	288	298	289	299
rect	288	301	289	302
rect	288	304	289	305
rect	288	313	289	314
rect	288	316	289	317
rect	288	322	289	323
rect	288	331	289	332
rect	288	337	289	338
rect	288	349	289	350
rect	288	352	289	353
rect	288	355	289	356
rect	288	361	289	362
rect	288	364	289	365
rect	289	7	290	8
rect	289	10	290	11
rect	289	13	290	14
rect	289	16	290	17
rect	289	22	290	23
rect	289	28	290	29
rect	289	31	290	32
rect	289	34	290	35
rect	289	37	290	38
rect	289	40	290	41
rect	289	55	290	56
rect	289	58	290	59
rect	289	67	290	68
rect	289	70	290	71
rect	289	76	290	77
rect	289	79	290	80
rect	289	82	290	83
rect	289	85	290	86
rect	289	88	290	89
rect	289	91	290	92
rect	289	97	290	98
rect	289	100	290	101
rect	289	103	290	104
rect	289	106	290	107
rect	289	115	290	116
rect	289	118	290	119
rect	289	121	290	122
rect	289	124	290	125
rect	289	136	290	137
rect	289	139	290	140
rect	289	142	290	143
rect	289	151	290	152
rect	289	154	290	155
rect	289	169	290	170
rect	289	172	290	173
rect	289	175	290	176
rect	289	178	290	179
rect	289	184	290	185
rect	289	187	290	188
rect	289	190	290	191
rect	289	193	290	194
rect	289	196	290	197
rect	289	199	290	200
rect	289	205	290	206
rect	289	208	290	209
rect	289	211	290	212
rect	289	217	290	218
rect	289	226	290	227
rect	289	229	290	230
rect	289	235	290	236
rect	289	244	290	245
rect	289	247	290	248
rect	289	250	290	251
rect	289	253	290	254
rect	289	262	290	263
rect	289	265	290	266
rect	289	268	290	269
rect	289	274	290	275
rect	289	277	290	278
rect	289	280	290	281
rect	289	286	290	287
rect	289	289	290	290
rect	289	292	290	293
rect	289	298	290	299
rect	289	301	290	302
rect	289	304	290	305
rect	289	307	290	308
rect	289	313	290	314
rect	289	316	290	317
rect	289	322	290	323
rect	289	331	290	332
rect	289	337	290	338
rect	289	346	290	347
rect	289	349	290	350
rect	289	352	290	353
rect	289	355	290	356
rect	289	361	290	362
rect	289	364	290	365
rect	290	7	291	8
rect	290	10	291	11
rect	290	16	291	17
rect	290	22	291	23
rect	290	28	291	29
rect	290	31	291	32
rect	290	34	291	35
rect	290	37	291	38
rect	290	40	291	41
rect	290	58	291	59
rect	290	67	291	68
rect	290	70	291	71
rect	290	76	291	77
rect	290	79	291	80
rect	290	82	291	83
rect	290	85	291	86
rect	290	88	291	89
rect	290	97	291	98
rect	290	100	291	101
rect	290	103	291	104
rect	290	106	291	107
rect	290	115	291	116
rect	290	118	291	119
rect	290	121	291	122
rect	290	124	291	125
rect	290	136	291	137
rect	290	139	291	140
rect	290	142	291	143
rect	290	151	291	152
rect	290	154	291	155
rect	290	169	291	170
rect	290	172	291	173
rect	290	175	291	176
rect	290	178	291	179
rect	290	184	291	185
rect	290	187	291	188
rect	290	190	291	191
rect	290	193	291	194
rect	290	196	291	197
rect	290	199	291	200
rect	290	208	291	209
rect	290	211	291	212
rect	290	217	291	218
rect	290	226	291	227
rect	290	235	291	236
rect	290	247	291	248
rect	290	250	291	251
rect	290	253	291	254
rect	290	262	291	263
rect	290	265	291	266
rect	290	268	291	269
rect	290	280	291	281
rect	290	286	291	287
rect	290	289	291	290
rect	290	292	291	293
rect	290	298	291	299
rect	290	304	291	305
rect	290	307	291	308
rect	290	313	291	314
rect	290	316	291	317
rect	290	331	291	332
rect	290	337	291	338
rect	290	346	291	347
rect	290	349	291	350
rect	290	352	291	353
rect	290	355	291	356
rect	290	361	291	362
rect	290	364	291	365
rect	291	7	292	8
rect	291	10	292	11
rect	291	16	292	17
rect	291	19	292	20
rect	291	22	292	23
rect	291	28	292	29
rect	291	31	292	32
rect	291	34	292	35
rect	291	37	292	38
rect	291	40	292	41
rect	291	58	292	59
rect	291	67	292	68
rect	291	70	292	71
rect	291	73	292	74
rect	291	76	292	77
rect	291	79	292	80
rect	291	82	292	83
rect	291	85	292	86
rect	291	88	292	89
rect	291	94	292	95
rect	291	97	292	98
rect	291	100	292	101
rect	291	103	292	104
rect	291	106	292	107
rect	291	115	292	116
rect	291	118	292	119
rect	291	121	292	122
rect	291	124	292	125
rect	291	127	292	128
rect	291	136	292	137
rect	291	139	292	140
rect	291	142	292	143
rect	291	151	292	152
rect	291	154	292	155
rect	291	169	292	170
rect	291	172	292	173
rect	291	175	292	176
rect	291	178	292	179
rect	291	181	292	182
rect	291	184	292	185
rect	291	187	292	188
rect	291	190	292	191
rect	291	193	292	194
rect	291	196	292	197
rect	291	199	292	200
rect	291	208	292	209
rect	291	211	292	212
rect	291	214	292	215
rect	291	217	292	218
rect	291	226	292	227
rect	291	235	292	236
rect	291	238	292	239
rect	291	247	292	248
rect	291	250	292	251
rect	291	253	292	254
rect	291	259	292	260
rect	291	262	292	263
rect	291	265	292	266
rect	291	268	292	269
rect	291	271	292	272
rect	291	280	292	281
rect	291	283	292	284
rect	291	286	292	287
rect	291	289	292	290
rect	291	292	292	293
rect	291	298	292	299
rect	291	304	292	305
rect	291	307	292	308
rect	291	313	292	314
rect	291	316	292	317
rect	291	319	292	320
rect	291	331	292	332
rect	291	337	292	338
rect	291	340	292	341
rect	291	346	292	347
rect	291	349	292	350
rect	291	352	292	353
rect	291	355	292	356
rect	291	361	292	362
rect	291	364	292	365
rect	292	10	293	11
rect	292	16	293	17
rect	292	19	293	20
rect	292	22	293	23
rect	292	28	293	29
rect	292	31	293	32
rect	292	34	293	35
rect	292	37	293	38
rect	292	58	293	59
rect	292	67	293	68
rect	292	70	293	71
rect	292	73	293	74
rect	292	76	293	77
rect	292	79	293	80
rect	292	82	293	83
rect	292	85	293	86
rect	292	88	293	89
rect	292	94	293	95
rect	292	97	293	98
rect	292	100	293	101
rect	292	103	293	104
rect	292	106	293	107
rect	292	115	293	116
rect	292	118	293	119
rect	292	121	293	122
rect	292	124	293	125
rect	292	127	293	128
rect	292	136	293	137
rect	292	139	293	140
rect	292	142	293	143
rect	292	151	293	152
rect	292	154	293	155
rect	292	169	293	170
rect	292	172	293	173
rect	292	175	293	176
rect	292	178	293	179
rect	292	181	293	182
rect	292	184	293	185
rect	292	187	293	188
rect	292	190	293	191
rect	292	193	293	194
rect	292	196	293	197
rect	292	199	293	200
rect	292	208	293	209
rect	292	211	293	212
rect	292	214	293	215
rect	292	217	293	218
rect	292	226	293	227
rect	292	235	293	236
rect	292	238	293	239
rect	292	247	293	248
rect	292	250	293	251
rect	292	253	293	254
rect	292	259	293	260
rect	292	262	293	263
rect	292	265	293	266
rect	292	268	293	269
rect	292	271	293	272
rect	292	280	293	281
rect	292	283	293	284
rect	292	286	293	287
rect	292	289	293	290
rect	292	292	293	293
rect	292	298	293	299
rect	292	304	293	305
rect	292	307	293	308
rect	292	313	293	314
rect	292	316	293	317
rect	292	319	293	320
rect	292	331	293	332
rect	292	340	293	341
rect	292	346	293	347
rect	292	349	293	350
rect	292	352	293	353
rect	292	355	293	356
rect	292	361	293	362
rect	292	364	293	365
rect	293	10	294	11
rect	293	13	294	14
rect	293	16	294	17
rect	293	19	294	20
rect	293	22	294	23
rect	293	28	294	29
rect	293	31	294	32
rect	293	34	294	35
rect	293	37	294	38
rect	293	46	294	47
rect	293	49	294	50
rect	293	58	294	59
rect	293	67	294	68
rect	293	70	294	71
rect	293	73	294	74
rect	293	76	294	77
rect	293	79	294	80
rect	293	82	294	83
rect	293	85	294	86
rect	293	88	294	89
rect	293	94	294	95
rect	293	97	294	98
rect	293	100	294	101
rect	293	103	294	104
rect	293	106	294	107
rect	293	115	294	116
rect	293	118	294	119
rect	293	121	294	122
rect	293	124	294	125
rect	293	127	294	128
rect	293	136	294	137
rect	293	139	294	140
rect	293	142	294	143
rect	293	151	294	152
rect	293	154	294	155
rect	293	169	294	170
rect	293	172	294	173
rect	293	175	294	176
rect	293	178	294	179
rect	293	181	294	182
rect	293	184	294	185
rect	293	187	294	188
rect	293	190	294	191
rect	293	193	294	194
rect	293	196	294	197
rect	293	199	294	200
rect	293	208	294	209
rect	293	211	294	212
rect	293	214	294	215
rect	293	217	294	218
rect	293	226	294	227
rect	293	235	294	236
rect	293	238	294	239
rect	293	247	294	248
rect	293	250	294	251
rect	293	253	294	254
rect	293	259	294	260
rect	293	262	294	263
rect	293	265	294	266
rect	293	268	294	269
rect	293	271	294	272
rect	293	280	294	281
rect	293	283	294	284
rect	293	286	294	287
rect	293	289	294	290
rect	293	292	294	293
rect	293	295	294	296
rect	293	298	294	299
rect	293	301	294	302
rect	293	304	294	305
rect	293	307	294	308
rect	293	310	294	311
rect	293	313	294	314
rect	293	316	294	317
rect	293	319	294	320
rect	293	322	294	323
rect	293	331	294	332
rect	293	340	294	341
rect	293	346	294	347
rect	293	349	294	350
rect	293	352	294	353
rect	293	355	294	356
rect	293	361	294	362
rect	293	364	294	365
rect	300	13	301	14
rect	300	16	301	17
rect	300	19	301	20
rect	300	22	301	23
rect	300	28	301	29
rect	300	31	301	32
rect	300	34	301	35
rect	300	37	301	38
rect	300	46	301	47
rect	300	49	301	50
rect	300	58	301	59
rect	300	61	301	62
rect	300	67	301	68
rect	300	70	301	71
rect	300	73	301	74
rect	300	76	301	77
rect	300	79	301	80
rect	300	82	301	83
rect	300	85	301	86
rect	300	88	301	89
rect	300	94	301	95
rect	300	97	301	98
rect	300	100	301	101
rect	300	103	301	104
rect	300	106	301	107
rect	300	115	301	116
rect	300	118	301	119
rect	300	121	301	122
rect	300	124	301	125
rect	300	127	301	128
rect	300	133	301	134
rect	300	136	301	137
rect	300	139	301	140
rect	300	142	301	143
rect	300	148	301	149
rect	300	151	301	152
rect	300	154	301	155
rect	300	169	301	170
rect	300	172	301	173
rect	300	175	301	176
rect	300	178	301	179
rect	300	187	301	188
rect	300	190	301	191
rect	300	193	301	194
rect	300	196	301	197
rect	300	199	301	200
rect	300	208	301	209
rect	300	211	301	212
rect	300	214	301	215
rect	300	217	301	218
rect	300	223	301	224
rect	300	226	301	227
rect	300	232	301	233
rect	300	235	301	236
rect	300	238	301	239
rect	300	247	301	248
rect	300	250	301	251
rect	300	259	301	260
rect	300	262	301	263
rect	300	265	301	266
rect	300	268	301	269
rect	300	271	301	272
rect	300	274	301	275
rect	300	280	301	281
rect	300	283	301	284
rect	300	286	301	287
rect	300	289	301	290
rect	300	292	301	293
rect	300	301	301	302
rect	300	304	301	305
rect	300	307	301	308
rect	300	313	301	314
rect	300	316	301	317
rect	300	319	301	320
rect	300	322	301	323
rect	300	331	301	332
rect	300	340	301	341
rect	300	349	301	350
rect	300	352	301	353
rect	300	358	301	359
rect	300	361	301	362
rect	300	364	301	365
rect	301	13	302	14
rect	301	16	302	17
rect	301	19	302	20
rect	301	22	302	23
rect	301	28	302	29
rect	301	31	302	32
rect	301	34	302	35
rect	301	37	302	38
rect	301	46	302	47
rect	301	49	302	50
rect	301	58	302	59
rect	301	61	302	62
rect	301	67	302	68
rect	301	70	302	71
rect	301	73	302	74
rect	301	76	302	77
rect	301	79	302	80
rect	301	82	302	83
rect	301	85	302	86
rect	301	88	302	89
rect	301	94	302	95
rect	301	97	302	98
rect	301	100	302	101
rect	301	103	302	104
rect	301	106	302	107
rect	301	115	302	116
rect	301	118	302	119
rect	301	121	302	122
rect	301	124	302	125
rect	301	127	302	128
rect	301	133	302	134
rect	301	136	302	137
rect	301	139	302	140
rect	301	142	302	143
rect	301	148	302	149
rect	301	151	302	152
rect	301	154	302	155
rect	301	169	302	170
rect	301	172	302	173
rect	301	175	302	176
rect	301	178	302	179
rect	301	187	302	188
rect	301	190	302	191
rect	301	193	302	194
rect	301	196	302	197
rect	301	199	302	200
rect	301	208	302	209
rect	301	211	302	212
rect	301	214	302	215
rect	301	217	302	218
rect	301	223	302	224
rect	301	226	302	227
rect	301	232	302	233
rect	301	235	302	236
rect	301	247	302	248
rect	301	250	302	251
rect	301	259	302	260
rect	301	262	302	263
rect	301	265	302	266
rect	301	268	302	269
rect	301	271	302	272
rect	301	274	302	275
rect	301	280	302	281
rect	301	283	302	284
rect	301	286	302	287
rect	301	289	302	290
rect	301	292	302	293
rect	301	301	302	302
rect	301	304	302	305
rect	301	307	302	308
rect	301	313	302	314
rect	301	316	302	317
rect	301	319	302	320
rect	301	322	302	323
rect	301	331	302	332
rect	301	340	302	341
rect	301	349	302	350
rect	301	352	302	353
rect	301	358	302	359
rect	301	361	302	362
rect	301	364	302	365
rect	302	13	303	14
rect	302	16	303	17
rect	302	19	303	20
rect	302	22	303	23
rect	302	28	303	29
rect	302	31	303	32
rect	302	34	303	35
rect	302	37	303	38
rect	302	46	303	47
rect	302	49	303	50
rect	302	58	303	59
rect	302	61	303	62
rect	302	67	303	68
rect	302	70	303	71
rect	302	73	303	74
rect	302	76	303	77
rect	302	79	303	80
rect	302	82	303	83
rect	302	85	303	86
rect	302	88	303	89
rect	302	94	303	95
rect	302	97	303	98
rect	302	100	303	101
rect	302	103	303	104
rect	302	106	303	107
rect	302	115	303	116
rect	302	118	303	119
rect	302	121	303	122
rect	302	124	303	125
rect	302	127	303	128
rect	302	133	303	134
rect	302	136	303	137
rect	302	139	303	140
rect	302	142	303	143
rect	302	148	303	149
rect	302	151	303	152
rect	302	154	303	155
rect	302	169	303	170
rect	302	172	303	173
rect	302	175	303	176
rect	302	178	303	179
rect	302	187	303	188
rect	302	190	303	191
rect	302	193	303	194
rect	302	196	303	197
rect	302	199	303	200
rect	302	208	303	209
rect	302	211	303	212
rect	302	214	303	215
rect	302	217	303	218
rect	302	223	303	224
rect	302	226	303	227
rect	302	232	303	233
rect	302	235	303	236
rect	302	247	303	248
rect	302	250	303	251
rect	302	253	303	254
rect	302	259	303	260
rect	302	262	303	263
rect	302	265	303	266
rect	302	268	303	269
rect	302	271	303	272
rect	302	274	303	275
rect	302	280	303	281
rect	302	283	303	284
rect	302	286	303	287
rect	302	289	303	290
rect	302	292	303	293
rect	302	301	303	302
rect	302	304	303	305
rect	302	307	303	308
rect	302	313	303	314
rect	302	316	303	317
rect	302	319	303	320
rect	302	322	303	323
rect	302	331	303	332
rect	302	340	303	341
rect	302	349	303	350
rect	302	352	303	353
rect	302	358	303	359
rect	302	361	303	362
rect	302	364	303	365
rect	303	13	304	14
rect	303	16	304	17
rect	303	19	304	20
rect	303	22	304	23
rect	303	28	304	29
rect	303	31	304	32
rect	303	34	304	35
rect	303	37	304	38
rect	303	46	304	47
rect	303	49	304	50
rect	303	58	304	59
rect	303	61	304	62
rect	303	67	304	68
rect	303	70	304	71
rect	303	73	304	74
rect	303	76	304	77
rect	303	79	304	80
rect	303	82	304	83
rect	303	85	304	86
rect	303	88	304	89
rect	303	94	304	95
rect	303	97	304	98
rect	303	100	304	101
rect	303	103	304	104
rect	303	106	304	107
rect	303	115	304	116
rect	303	118	304	119
rect	303	121	304	122
rect	303	124	304	125
rect	303	127	304	128
rect	303	133	304	134
rect	303	136	304	137
rect	303	139	304	140
rect	303	142	304	143
rect	303	148	304	149
rect	303	151	304	152
rect	303	154	304	155
rect	303	169	304	170
rect	303	172	304	173
rect	303	175	304	176
rect	303	178	304	179
rect	303	187	304	188
rect	303	190	304	191
rect	303	193	304	194
rect	303	196	304	197
rect	303	199	304	200
rect	303	208	304	209
rect	303	211	304	212
rect	303	214	304	215
rect	303	217	304	218
rect	303	223	304	224
rect	303	232	304	233
rect	303	235	304	236
rect	303	247	304	248
rect	303	250	304	251
rect	303	253	304	254
rect	303	259	304	260
rect	303	262	304	263
rect	303	265	304	266
rect	303	268	304	269
rect	303	271	304	272
rect	303	274	304	275
rect	303	280	304	281
rect	303	283	304	284
rect	303	286	304	287
rect	303	289	304	290
rect	303	292	304	293
rect	303	301	304	302
rect	303	304	304	305
rect	303	307	304	308
rect	303	313	304	314
rect	303	316	304	317
rect	303	319	304	320
rect	303	322	304	323
rect	303	331	304	332
rect	303	340	304	341
rect	303	349	304	350
rect	303	352	304	353
rect	303	358	304	359
rect	303	361	304	362
rect	303	364	304	365
rect	304	13	305	14
rect	304	16	305	17
rect	304	19	305	20
rect	304	22	305	23
rect	304	28	305	29
rect	304	31	305	32
rect	304	34	305	35
rect	304	37	305	38
rect	304	46	305	47
rect	304	49	305	50
rect	304	58	305	59
rect	304	61	305	62
rect	304	67	305	68
rect	304	70	305	71
rect	304	73	305	74
rect	304	76	305	77
rect	304	79	305	80
rect	304	82	305	83
rect	304	85	305	86
rect	304	88	305	89
rect	304	94	305	95
rect	304	97	305	98
rect	304	100	305	101
rect	304	103	305	104
rect	304	106	305	107
rect	304	115	305	116
rect	304	118	305	119
rect	304	121	305	122
rect	304	124	305	125
rect	304	127	305	128
rect	304	133	305	134
rect	304	136	305	137
rect	304	139	305	140
rect	304	142	305	143
rect	304	148	305	149
rect	304	151	305	152
rect	304	154	305	155
rect	304	169	305	170
rect	304	172	305	173
rect	304	175	305	176
rect	304	178	305	179
rect	304	187	305	188
rect	304	190	305	191
rect	304	193	305	194
rect	304	196	305	197
rect	304	199	305	200
rect	304	208	305	209
rect	304	211	305	212
rect	304	214	305	215
rect	304	217	305	218
rect	304	223	305	224
rect	304	232	305	233
rect	304	235	305	236
rect	304	241	305	242
rect	304	247	305	248
rect	304	250	305	251
rect	304	253	305	254
rect	304	259	305	260
rect	304	262	305	263
rect	304	265	305	266
rect	304	268	305	269
rect	304	271	305	272
rect	304	274	305	275
rect	304	280	305	281
rect	304	283	305	284
rect	304	286	305	287
rect	304	289	305	290
rect	304	292	305	293
rect	304	301	305	302
rect	304	304	305	305
rect	304	307	305	308
rect	304	313	305	314
rect	304	316	305	317
rect	304	319	305	320
rect	304	322	305	323
rect	304	331	305	332
rect	304	340	305	341
rect	304	349	305	350
rect	304	352	305	353
rect	304	358	305	359
rect	304	361	305	362
rect	304	364	305	365
rect	305	13	306	14
rect	305	16	306	17
rect	305	19	306	20
rect	305	22	306	23
rect	305	28	306	29
rect	305	31	306	32
rect	305	34	306	35
rect	305	37	306	38
rect	305	46	306	47
rect	305	49	306	50
rect	305	58	306	59
rect	305	61	306	62
rect	305	67	306	68
rect	305	70	306	71
rect	305	73	306	74
rect	305	76	306	77
rect	305	79	306	80
rect	305	82	306	83
rect	305	85	306	86
rect	305	88	306	89
rect	305	94	306	95
rect	305	97	306	98
rect	305	100	306	101
rect	305	103	306	104
rect	305	106	306	107
rect	305	115	306	116
rect	305	118	306	119
rect	305	121	306	122
rect	305	124	306	125
rect	305	127	306	128
rect	305	133	306	134
rect	305	136	306	137
rect	305	139	306	140
rect	305	142	306	143
rect	305	148	306	149
rect	305	151	306	152
rect	305	154	306	155
rect	305	169	306	170
rect	305	172	306	173
rect	305	175	306	176
rect	305	178	306	179
rect	305	187	306	188
rect	305	190	306	191
rect	305	193	306	194
rect	305	196	306	197
rect	305	199	306	200
rect	305	211	306	212
rect	305	214	306	215
rect	305	217	306	218
rect	305	223	306	224
rect	305	232	306	233
rect	305	235	306	236
rect	305	241	306	242
rect	305	247	306	248
rect	305	250	306	251
rect	305	253	306	254
rect	305	259	306	260
rect	305	262	306	263
rect	305	265	306	266
rect	305	268	306	269
rect	305	271	306	272
rect	305	274	306	275
rect	305	280	306	281
rect	305	283	306	284
rect	305	286	306	287
rect	305	289	306	290
rect	305	292	306	293
rect	305	301	306	302
rect	305	304	306	305
rect	305	307	306	308
rect	305	313	306	314
rect	305	316	306	317
rect	305	319	306	320
rect	305	322	306	323
rect	305	331	306	332
rect	305	340	306	341
rect	305	349	306	350
rect	305	352	306	353
rect	305	358	306	359
rect	305	361	306	362
rect	305	364	306	365
rect	306	13	307	14
rect	306	16	307	17
rect	306	19	307	20
rect	306	22	307	23
rect	306	28	307	29
rect	306	31	307	32
rect	306	34	307	35
rect	306	37	307	38
rect	306	46	307	47
rect	306	49	307	50
rect	306	58	307	59
rect	306	61	307	62
rect	306	67	307	68
rect	306	70	307	71
rect	306	73	307	74
rect	306	76	307	77
rect	306	79	307	80
rect	306	82	307	83
rect	306	85	307	86
rect	306	88	307	89
rect	306	94	307	95
rect	306	97	307	98
rect	306	100	307	101
rect	306	103	307	104
rect	306	106	307	107
rect	306	115	307	116
rect	306	118	307	119
rect	306	121	307	122
rect	306	124	307	125
rect	306	127	307	128
rect	306	133	307	134
rect	306	136	307	137
rect	306	139	307	140
rect	306	142	307	143
rect	306	148	307	149
rect	306	151	307	152
rect	306	154	307	155
rect	306	169	307	170
rect	306	172	307	173
rect	306	175	307	176
rect	306	178	307	179
rect	306	187	307	188
rect	306	190	307	191
rect	306	193	307	194
rect	306	196	307	197
rect	306	199	307	200
rect	306	211	307	212
rect	306	214	307	215
rect	306	217	307	218
rect	306	223	307	224
rect	306	232	307	233
rect	306	235	307	236
rect	306	238	307	239
rect	306	241	307	242
rect	306	247	307	248
rect	306	250	307	251
rect	306	253	307	254
rect	306	259	307	260
rect	306	262	307	263
rect	306	265	307	266
rect	306	268	307	269
rect	306	271	307	272
rect	306	274	307	275
rect	306	280	307	281
rect	306	283	307	284
rect	306	286	307	287
rect	306	289	307	290
rect	306	292	307	293
rect	306	301	307	302
rect	306	304	307	305
rect	306	307	307	308
rect	306	313	307	314
rect	306	316	307	317
rect	306	319	307	320
rect	306	322	307	323
rect	306	331	307	332
rect	306	340	307	341
rect	306	349	307	350
rect	306	352	307	353
rect	306	358	307	359
rect	306	361	307	362
rect	306	364	307	365
rect	307	13	308	14
rect	307	16	308	17
rect	307	19	308	20
rect	307	22	308	23
rect	307	28	308	29
rect	307	31	308	32
rect	307	34	308	35
rect	307	37	308	38
rect	307	46	308	47
rect	307	49	308	50
rect	307	58	308	59
rect	307	61	308	62
rect	307	67	308	68
rect	307	70	308	71
rect	307	73	308	74
rect	307	76	308	77
rect	307	79	308	80
rect	307	82	308	83
rect	307	85	308	86
rect	307	88	308	89
rect	307	94	308	95
rect	307	97	308	98
rect	307	100	308	101
rect	307	103	308	104
rect	307	106	308	107
rect	307	115	308	116
rect	307	118	308	119
rect	307	121	308	122
rect	307	124	308	125
rect	307	127	308	128
rect	307	133	308	134
rect	307	136	308	137
rect	307	139	308	140
rect	307	142	308	143
rect	307	148	308	149
rect	307	151	308	152
rect	307	154	308	155
rect	307	169	308	170
rect	307	172	308	173
rect	307	175	308	176
rect	307	178	308	179
rect	307	187	308	188
rect	307	190	308	191
rect	307	193	308	194
rect	307	199	308	200
rect	307	214	308	215
rect	307	217	308	218
rect	307	223	308	224
rect	307	232	308	233
rect	307	235	308	236
rect	307	238	308	239
rect	307	241	308	242
rect	307	247	308	248
rect	307	250	308	251
rect	307	253	308	254
rect	307	259	308	260
rect	307	262	308	263
rect	307	265	308	266
rect	307	268	308	269
rect	307	271	308	272
rect	307	274	308	275
rect	307	280	308	281
rect	307	283	308	284
rect	307	286	308	287
rect	307	289	308	290
rect	307	292	308	293
rect	307	301	308	302
rect	307	304	308	305
rect	307	307	308	308
rect	307	313	308	314
rect	307	316	308	317
rect	307	319	308	320
rect	307	322	308	323
rect	307	331	308	332
rect	307	340	308	341
rect	307	349	308	350
rect	307	352	308	353
rect	307	358	308	359
rect	307	361	308	362
rect	307	364	308	365
rect	308	13	309	14
rect	308	16	309	17
rect	308	19	309	20
rect	308	22	309	23
rect	308	28	309	29
rect	308	31	309	32
rect	308	34	309	35
rect	308	37	309	38
rect	308	46	309	47
rect	308	49	309	50
rect	308	58	309	59
rect	308	61	309	62
rect	308	67	309	68
rect	308	70	309	71
rect	308	73	309	74
rect	308	76	309	77
rect	308	79	309	80
rect	308	82	309	83
rect	308	85	309	86
rect	308	88	309	89
rect	308	94	309	95
rect	308	97	309	98
rect	308	100	309	101
rect	308	103	309	104
rect	308	106	309	107
rect	308	115	309	116
rect	308	118	309	119
rect	308	121	309	122
rect	308	124	309	125
rect	308	127	309	128
rect	308	133	309	134
rect	308	136	309	137
rect	308	139	309	140
rect	308	142	309	143
rect	308	148	309	149
rect	308	151	309	152
rect	308	154	309	155
rect	308	169	309	170
rect	308	172	309	173
rect	308	175	309	176
rect	308	178	309	179
rect	308	187	309	188
rect	308	190	309	191
rect	308	193	309	194
rect	308	199	309	200
rect	308	208	309	209
rect	308	214	309	215
rect	308	217	309	218
rect	308	223	309	224
rect	308	226	309	227
rect	308	232	309	233
rect	308	235	309	236
rect	308	238	309	239
rect	308	241	309	242
rect	308	247	309	248
rect	308	250	309	251
rect	308	253	309	254
rect	308	259	309	260
rect	308	262	309	263
rect	308	265	309	266
rect	308	268	309	269
rect	308	271	309	272
rect	308	274	309	275
rect	308	280	309	281
rect	308	283	309	284
rect	308	286	309	287
rect	308	289	309	290
rect	308	292	309	293
rect	308	301	309	302
rect	308	304	309	305
rect	308	307	309	308
rect	308	313	309	314
rect	308	316	309	317
rect	308	319	309	320
rect	308	322	309	323
rect	308	331	309	332
rect	308	340	309	341
rect	308	349	309	350
rect	308	352	309	353
rect	308	358	309	359
rect	308	361	309	362
rect	308	364	309	365
rect	309	13	310	14
rect	309	16	310	17
rect	309	19	310	20
rect	309	22	310	23
rect	309	28	310	29
rect	309	31	310	32
rect	309	34	310	35
rect	309	37	310	38
rect	309	46	310	47
rect	309	49	310	50
rect	309	58	310	59
rect	309	61	310	62
rect	309	67	310	68
rect	309	70	310	71
rect	309	73	310	74
rect	309	76	310	77
rect	309	79	310	80
rect	309	82	310	83
rect	309	85	310	86
rect	309	88	310	89
rect	309	94	310	95
rect	309	97	310	98
rect	309	100	310	101
rect	309	103	310	104
rect	309	106	310	107
rect	309	115	310	116
rect	309	118	310	119
rect	309	121	310	122
rect	309	124	310	125
rect	309	127	310	128
rect	309	133	310	134
rect	309	136	310	137
rect	309	139	310	140
rect	309	142	310	143
rect	309	148	310	149
rect	309	151	310	152
rect	309	154	310	155
rect	309	169	310	170
rect	309	172	310	173
rect	309	175	310	176
rect	309	178	310	179
rect	309	187	310	188
rect	309	190	310	191
rect	309	199	310	200
rect	309	208	310	209
rect	309	214	310	215
rect	309	217	310	218
rect	309	223	310	224
rect	309	226	310	227
rect	309	232	310	233
rect	309	235	310	236
rect	309	238	310	239
rect	309	241	310	242
rect	309	247	310	248
rect	309	250	310	251
rect	309	253	310	254
rect	309	259	310	260
rect	309	262	310	263
rect	309	265	310	266
rect	309	268	310	269
rect	309	271	310	272
rect	309	274	310	275
rect	309	280	310	281
rect	309	283	310	284
rect	309	286	310	287
rect	309	289	310	290
rect	309	292	310	293
rect	309	301	310	302
rect	309	304	310	305
rect	309	307	310	308
rect	309	313	310	314
rect	309	316	310	317
rect	309	319	310	320
rect	309	322	310	323
rect	309	331	310	332
rect	309	340	310	341
rect	309	349	310	350
rect	309	352	310	353
rect	309	358	310	359
rect	309	361	310	362
rect	309	364	310	365
rect	310	13	311	14
rect	310	16	311	17
rect	310	19	311	20
rect	310	22	311	23
rect	310	28	311	29
rect	310	31	311	32
rect	310	34	311	35
rect	310	37	311	38
rect	310	46	311	47
rect	310	49	311	50
rect	310	58	311	59
rect	310	61	311	62
rect	310	67	311	68
rect	310	70	311	71
rect	310	73	311	74
rect	310	76	311	77
rect	310	79	311	80
rect	310	82	311	83
rect	310	85	311	86
rect	310	88	311	89
rect	310	94	311	95
rect	310	97	311	98
rect	310	100	311	101
rect	310	103	311	104
rect	310	106	311	107
rect	310	115	311	116
rect	310	118	311	119
rect	310	121	311	122
rect	310	124	311	125
rect	310	127	311	128
rect	310	133	311	134
rect	310	136	311	137
rect	310	139	311	140
rect	310	142	311	143
rect	310	148	311	149
rect	310	151	311	152
rect	310	154	311	155
rect	310	169	311	170
rect	310	172	311	173
rect	310	175	311	176
rect	310	178	311	179
rect	310	187	311	188
rect	310	190	311	191
rect	310	199	311	200
rect	310	208	311	209
rect	310	211	311	212
rect	310	214	311	215
rect	310	217	311	218
rect	310	223	311	224
rect	310	226	311	227
rect	310	232	311	233
rect	310	235	311	236
rect	310	238	311	239
rect	310	241	311	242
rect	310	247	311	248
rect	310	250	311	251
rect	310	253	311	254
rect	310	259	311	260
rect	310	262	311	263
rect	310	265	311	266
rect	310	268	311	269
rect	310	271	311	272
rect	310	274	311	275
rect	310	280	311	281
rect	310	283	311	284
rect	310	286	311	287
rect	310	289	311	290
rect	310	292	311	293
rect	310	301	311	302
rect	310	304	311	305
rect	310	307	311	308
rect	310	313	311	314
rect	310	316	311	317
rect	310	319	311	320
rect	310	322	311	323
rect	310	331	311	332
rect	310	340	311	341
rect	310	349	311	350
rect	310	352	311	353
rect	310	358	311	359
rect	310	361	311	362
rect	310	364	311	365
rect	311	13	312	14
rect	311	16	312	17
rect	311	19	312	20
rect	311	22	312	23
rect	311	28	312	29
rect	311	31	312	32
rect	311	34	312	35
rect	311	37	312	38
rect	311	46	312	47
rect	311	49	312	50
rect	311	58	312	59
rect	311	61	312	62
rect	311	67	312	68
rect	311	70	312	71
rect	311	73	312	74
rect	311	76	312	77
rect	311	79	312	80
rect	311	82	312	83
rect	311	85	312	86
rect	311	88	312	89
rect	311	94	312	95
rect	311	97	312	98
rect	311	100	312	101
rect	311	103	312	104
rect	311	106	312	107
rect	311	115	312	116
rect	311	118	312	119
rect	311	121	312	122
rect	311	124	312	125
rect	311	127	312	128
rect	311	133	312	134
rect	311	136	312	137
rect	311	139	312	140
rect	311	142	312	143
rect	311	148	312	149
rect	311	154	312	155
rect	311	169	312	170
rect	311	172	312	173
rect	311	178	312	179
rect	311	187	312	188
rect	311	190	312	191
rect	311	199	312	200
rect	311	208	312	209
rect	311	211	312	212
rect	311	214	312	215
rect	311	217	312	218
rect	311	223	312	224
rect	311	226	312	227
rect	311	232	312	233
rect	311	235	312	236
rect	311	238	312	239
rect	311	241	312	242
rect	311	247	312	248
rect	311	250	312	251
rect	311	253	312	254
rect	311	259	312	260
rect	311	262	312	263
rect	311	265	312	266
rect	311	268	312	269
rect	311	271	312	272
rect	311	274	312	275
rect	311	280	312	281
rect	311	283	312	284
rect	311	286	312	287
rect	311	289	312	290
rect	311	292	312	293
rect	311	301	312	302
rect	311	304	312	305
rect	311	307	312	308
rect	311	313	312	314
rect	311	316	312	317
rect	311	319	312	320
rect	311	322	312	323
rect	311	331	312	332
rect	311	340	312	341
rect	311	349	312	350
rect	311	352	312	353
rect	311	358	312	359
rect	311	361	312	362
rect	311	364	312	365
rect	312	13	313	14
rect	312	16	313	17
rect	312	19	313	20
rect	312	22	313	23
rect	312	28	313	29
rect	312	31	313	32
rect	312	34	313	35
rect	312	37	313	38
rect	312	46	313	47
rect	312	49	313	50
rect	312	58	313	59
rect	312	61	313	62
rect	312	67	313	68
rect	312	70	313	71
rect	312	73	313	74
rect	312	76	313	77
rect	312	79	313	80
rect	312	82	313	83
rect	312	85	313	86
rect	312	88	313	89
rect	312	94	313	95
rect	312	97	313	98
rect	312	100	313	101
rect	312	103	313	104
rect	312	106	313	107
rect	312	115	313	116
rect	312	118	313	119
rect	312	121	313	122
rect	312	124	313	125
rect	312	127	313	128
rect	312	133	313	134
rect	312	136	313	137
rect	312	139	313	140
rect	312	142	313	143
rect	312	148	313	149
rect	312	154	313	155
rect	312	166	313	167
rect	312	169	313	170
rect	312	172	313	173
rect	312	178	313	179
rect	312	187	313	188
rect	312	190	313	191
rect	312	196	313	197
rect	312	199	313	200
rect	312	208	313	209
rect	312	211	313	212
rect	312	214	313	215
rect	312	217	313	218
rect	312	223	313	224
rect	312	226	313	227
rect	312	232	313	233
rect	312	235	313	236
rect	312	238	313	239
rect	312	241	313	242
rect	312	247	313	248
rect	312	250	313	251
rect	312	253	313	254
rect	312	259	313	260
rect	312	262	313	263
rect	312	265	313	266
rect	312	268	313	269
rect	312	271	313	272
rect	312	274	313	275
rect	312	280	313	281
rect	312	283	313	284
rect	312	286	313	287
rect	312	289	313	290
rect	312	292	313	293
rect	312	301	313	302
rect	312	304	313	305
rect	312	307	313	308
rect	312	313	313	314
rect	312	316	313	317
rect	312	319	313	320
rect	312	322	313	323
rect	312	331	313	332
rect	312	340	313	341
rect	312	349	313	350
rect	312	352	313	353
rect	312	358	313	359
rect	312	361	313	362
rect	312	364	313	365
rect	313	13	314	14
rect	313	16	314	17
rect	313	19	314	20
rect	313	22	314	23
rect	313	28	314	29
rect	313	31	314	32
rect	313	34	314	35
rect	313	37	314	38
rect	313	46	314	47
rect	313	49	314	50
rect	313	58	314	59
rect	313	61	314	62
rect	313	67	314	68
rect	313	70	314	71
rect	313	73	314	74
rect	313	76	314	77
rect	313	79	314	80
rect	313	82	314	83
rect	313	85	314	86
rect	313	88	314	89
rect	313	94	314	95
rect	313	97	314	98
rect	313	100	314	101
rect	313	103	314	104
rect	313	106	314	107
rect	313	115	314	116
rect	313	118	314	119
rect	313	121	314	122
rect	313	127	314	128
rect	313	133	314	134
rect	313	136	314	137
rect	313	139	314	140
rect	313	142	314	143
rect	313	154	314	155
rect	313	166	314	167
rect	313	169	314	170
rect	313	172	314	173
rect	313	190	314	191
rect	313	196	314	197
rect	313	199	314	200
rect	313	208	314	209
rect	313	211	314	212
rect	313	214	314	215
rect	313	217	314	218
rect	313	223	314	224
rect	313	226	314	227
rect	313	232	314	233
rect	313	235	314	236
rect	313	238	314	239
rect	313	241	314	242
rect	313	247	314	248
rect	313	250	314	251
rect	313	253	314	254
rect	313	259	314	260
rect	313	262	314	263
rect	313	265	314	266
rect	313	268	314	269
rect	313	271	314	272
rect	313	274	314	275
rect	313	280	314	281
rect	313	283	314	284
rect	313	286	314	287
rect	313	289	314	290
rect	313	292	314	293
rect	313	301	314	302
rect	313	304	314	305
rect	313	307	314	308
rect	313	313	314	314
rect	313	316	314	317
rect	313	319	314	320
rect	313	322	314	323
rect	313	331	314	332
rect	313	340	314	341
rect	313	349	314	350
rect	313	352	314	353
rect	313	358	314	359
rect	313	361	314	362
rect	313	364	314	365
rect	314	13	315	14
rect	314	16	315	17
rect	314	19	315	20
rect	314	22	315	23
rect	314	28	315	29
rect	314	31	315	32
rect	314	34	315	35
rect	314	37	315	38
rect	314	46	315	47
rect	314	49	315	50
rect	314	58	315	59
rect	314	61	315	62
rect	314	67	315	68
rect	314	70	315	71
rect	314	73	315	74
rect	314	76	315	77
rect	314	79	315	80
rect	314	82	315	83
rect	314	85	315	86
rect	314	88	315	89
rect	314	94	315	95
rect	314	97	315	98
rect	314	100	315	101
rect	314	103	315	104
rect	314	106	315	107
rect	314	115	315	116
rect	314	118	315	119
rect	314	121	315	122
rect	314	127	315	128
rect	314	130	315	131
rect	314	133	315	134
rect	314	136	315	137
rect	314	139	315	140
rect	314	142	315	143
rect	314	154	315	155
rect	314	166	315	167
rect	314	169	315	170
rect	314	172	315	173
rect	314	175	315	176
rect	314	184	315	185
rect	314	190	315	191
rect	314	196	315	197
rect	314	199	315	200
rect	314	205	315	206
rect	314	208	315	209
rect	314	211	315	212
rect	314	214	315	215
rect	314	217	315	218
rect	314	223	315	224
rect	314	226	315	227
rect	314	232	315	233
rect	314	235	315	236
rect	314	238	315	239
rect	314	241	315	242
rect	314	247	315	248
rect	314	250	315	251
rect	314	253	315	254
rect	314	259	315	260
rect	314	262	315	263
rect	314	265	315	266
rect	314	268	315	269
rect	314	271	315	272
rect	314	274	315	275
rect	314	280	315	281
rect	314	283	315	284
rect	314	286	315	287
rect	314	289	315	290
rect	314	292	315	293
rect	314	301	315	302
rect	314	304	315	305
rect	314	307	315	308
rect	314	313	315	314
rect	314	316	315	317
rect	314	319	315	320
rect	314	322	315	323
rect	314	331	315	332
rect	314	340	315	341
rect	314	349	315	350
rect	314	352	315	353
rect	314	358	315	359
rect	314	361	315	362
rect	314	364	315	365
rect	315	13	316	14
rect	315	16	316	17
rect	315	19	316	20
rect	315	22	316	23
rect	315	28	316	29
rect	315	31	316	32
rect	315	34	316	35
rect	315	37	316	38
rect	315	46	316	47
rect	315	49	316	50
rect	315	58	316	59
rect	315	67	316	68
rect	315	70	316	71
rect	315	73	316	74
rect	315	76	316	77
rect	315	79	316	80
rect	315	82	316	83
rect	315	85	316	86
rect	315	88	316	89
rect	315	94	316	95
rect	315	97	316	98
rect	315	100	316	101
rect	315	103	316	104
rect	315	106	316	107
rect	315	115	316	116
rect	315	118	316	119
rect	315	121	316	122
rect	315	127	316	128
rect	315	130	316	131
rect	315	133	316	134
rect	315	136	316	137
rect	315	139	316	140
rect	315	142	316	143
rect	315	154	316	155
rect	315	166	316	167
rect	315	169	316	170
rect	315	172	316	173
rect	315	175	316	176
rect	315	184	316	185
rect	315	190	316	191
rect	315	196	316	197
rect	315	199	316	200
rect	315	205	316	206
rect	315	208	316	209
rect	315	211	316	212
rect	315	214	316	215
rect	315	217	316	218
rect	315	223	316	224
rect	315	226	316	227
rect	315	232	316	233
rect	315	235	316	236
rect	315	238	316	239
rect	315	241	316	242
rect	315	247	316	248
rect	315	250	316	251
rect	315	253	316	254
rect	315	259	316	260
rect	315	262	316	263
rect	315	265	316	266
rect	315	268	316	269
rect	315	271	316	272
rect	315	274	316	275
rect	315	280	316	281
rect	315	283	316	284
rect	315	289	316	290
rect	315	292	316	293
rect	315	301	316	302
rect	315	304	316	305
rect	315	307	316	308
rect	315	313	316	314
rect	315	316	316	317
rect	315	319	316	320
rect	315	322	316	323
rect	315	331	316	332
rect	315	340	316	341
rect	315	349	316	350
rect	315	352	316	353
rect	315	358	316	359
rect	315	361	316	362
rect	315	364	316	365
rect	316	13	317	14
rect	316	16	317	17
rect	316	19	317	20
rect	316	22	317	23
rect	316	28	317	29
rect	316	31	317	32
rect	316	34	317	35
rect	316	37	317	38
rect	316	46	317	47
rect	316	49	317	50
rect	316	58	317	59
rect	316	67	317	68
rect	316	70	317	71
rect	316	73	317	74
rect	316	76	317	77
rect	316	79	317	80
rect	316	82	317	83
rect	316	85	317	86
rect	316	88	317	89
rect	316	94	317	95
rect	316	97	317	98
rect	316	100	317	101
rect	316	103	317	104
rect	316	106	317	107
rect	316	115	317	116
rect	316	118	317	119
rect	316	121	317	122
rect	316	127	317	128
rect	316	130	317	131
rect	316	133	317	134
rect	316	136	317	137
rect	316	139	317	140
rect	316	142	317	143
rect	316	154	317	155
rect	316	166	317	167
rect	316	169	317	170
rect	316	172	317	173
rect	316	175	317	176
rect	316	184	317	185
rect	316	190	317	191
rect	316	196	317	197
rect	316	199	317	200
rect	316	205	317	206
rect	316	208	317	209
rect	316	211	317	212
rect	316	214	317	215
rect	316	217	317	218
rect	316	223	317	224
rect	316	226	317	227
rect	316	232	317	233
rect	316	235	317	236
rect	316	238	317	239
rect	316	241	317	242
rect	316	247	317	248
rect	316	250	317	251
rect	316	253	317	254
rect	316	259	317	260
rect	316	262	317	263
rect	316	265	317	266
rect	316	268	317	269
rect	316	271	317	272
rect	316	274	317	275
rect	316	280	317	281
rect	316	283	317	284
rect	316	289	317	290
rect	316	292	317	293
rect	316	301	317	302
rect	316	304	317	305
rect	316	307	317	308
rect	316	313	317	314
rect	316	316	317	317
rect	316	319	317	320
rect	316	322	317	323
rect	316	331	317	332
rect	316	340	317	341
rect	316	349	317	350
rect	316	352	317	353
rect	316	358	317	359
rect	316	361	317	362
rect	316	364	317	365
rect	317	13	318	14
rect	317	16	318	17
rect	317	19	318	20
rect	317	22	318	23
rect	317	28	318	29
rect	317	31	318	32
rect	317	34	318	35
rect	317	37	318	38
rect	317	46	318	47
rect	317	49	318	50
rect	317	58	318	59
rect	317	67	318	68
rect	317	70	318	71
rect	317	73	318	74
rect	317	76	318	77
rect	317	79	318	80
rect	317	82	318	83
rect	317	85	318	86
rect	317	88	318	89
rect	317	94	318	95
rect	317	97	318	98
rect	317	100	318	101
rect	317	103	318	104
rect	317	106	318	107
rect	317	115	318	116
rect	317	121	318	122
rect	317	127	318	128
rect	317	130	318	131
rect	317	133	318	134
rect	317	136	318	137
rect	317	139	318	140
rect	317	142	318	143
rect	317	154	318	155
rect	317	166	318	167
rect	317	169	318	170
rect	317	175	318	176
rect	317	184	318	185
rect	317	190	318	191
rect	317	196	318	197
rect	317	205	318	206
rect	317	208	318	209
rect	317	211	318	212
rect	317	214	318	215
rect	317	223	318	224
rect	317	226	318	227
rect	317	232	318	233
rect	317	235	318	236
rect	317	238	318	239
rect	317	241	318	242
rect	317	247	318	248
rect	317	250	318	251
rect	317	253	318	254
rect	317	259	318	260
rect	317	262	318	263
rect	317	265	318	266
rect	317	271	318	272
rect	317	274	318	275
rect	317	280	318	281
rect	317	283	318	284
rect	317	289	318	290
rect	317	292	318	293
rect	317	301	318	302
rect	317	304	318	305
rect	317	307	318	308
rect	317	313	318	314
rect	317	316	318	317
rect	317	319	318	320
rect	317	322	318	323
rect	317	340	318	341
rect	317	349	318	350
rect	317	352	318	353
rect	317	358	318	359
rect	317	361	318	362
rect	317	364	318	365
rect	318	13	319	14
rect	318	16	319	17
rect	318	19	319	20
rect	318	22	319	23
rect	318	28	319	29
rect	318	31	319	32
rect	318	34	319	35
rect	318	37	319	38
rect	318	46	319	47
rect	318	49	319	50
rect	318	58	319	59
rect	318	67	319	68
rect	318	70	319	71
rect	318	73	319	74
rect	318	76	319	77
rect	318	79	319	80
rect	318	82	319	83
rect	318	85	319	86
rect	318	88	319	89
rect	318	94	319	95
rect	318	97	319	98
rect	318	100	319	101
rect	318	103	319	104
rect	318	106	319	107
rect	318	115	319	116
rect	318	121	319	122
rect	318	127	319	128
rect	318	130	319	131
rect	318	133	319	134
rect	318	136	319	137
rect	318	139	319	140
rect	318	142	319	143
rect	318	154	319	155
rect	318	157	319	158
rect	318	166	319	167
rect	318	169	319	170
rect	318	175	319	176
rect	318	178	319	179
rect	318	181	319	182
rect	318	184	319	185
rect	318	190	319	191
rect	318	196	319	197
rect	318	205	319	206
rect	318	208	319	209
rect	318	211	319	212
rect	318	214	319	215
rect	318	223	319	224
rect	318	226	319	227
rect	318	229	319	230
rect	318	232	319	233
rect	318	235	319	236
rect	318	238	319	239
rect	318	241	319	242
rect	318	247	319	248
rect	318	250	319	251
rect	318	253	319	254
rect	318	259	319	260
rect	318	262	319	263
rect	318	265	319	266
rect	318	271	319	272
rect	318	274	319	275
rect	318	280	319	281
rect	318	283	319	284
rect	318	286	319	287
rect	318	289	319	290
rect	318	292	319	293
rect	318	301	319	302
rect	318	304	319	305
rect	318	307	319	308
rect	318	313	319	314
rect	318	316	319	317
rect	318	319	319	320
rect	318	322	319	323
rect	318	340	319	341
rect	318	343	319	344
rect	318	349	319	350
rect	318	352	319	353
rect	318	358	319	359
rect	318	361	319	362
rect	318	364	319	365
rect	319	13	320	14
rect	319	16	320	17
rect	319	19	320	20
rect	319	22	320	23
rect	319	28	320	29
rect	319	31	320	32
rect	319	34	320	35
rect	319	37	320	38
rect	319	46	320	47
rect	319	49	320	50
rect	319	58	320	59
rect	319	67	320	68
rect	319	70	320	71
rect	319	73	320	74
rect	319	76	320	77
rect	319	79	320	80
rect	319	82	320	83
rect	319	85	320	86
rect	319	88	320	89
rect	319	94	320	95
rect	319	97	320	98
rect	319	100	320	101
rect	319	103	320	104
rect	319	121	320	122
rect	319	127	320	128
rect	319	130	320	131
rect	319	133	320	134
rect	319	136	320	137
rect	319	139	320	140
rect	319	142	320	143
rect	319	154	320	155
rect	319	157	320	158
rect	319	166	320	167
rect	319	175	320	176
rect	319	178	320	179
rect	319	181	320	182
rect	319	184	320	185
rect	319	190	320	191
rect	319	196	320	197
rect	319	205	320	206
rect	319	208	320	209
rect	319	211	320	212
rect	319	214	320	215
rect	319	223	320	224
rect	319	226	320	227
rect	319	229	320	230
rect	319	232	320	233
rect	319	235	320	236
rect	319	238	320	239
rect	319	241	320	242
rect	319	247	320	248
rect	319	250	320	251
rect	319	253	320	254
rect	319	259	320	260
rect	319	262	320	263
rect	319	271	320	272
rect	319	274	320	275
rect	319	280	320	281
rect	319	283	320	284
rect	319	286	320	287
rect	319	289	320	290
rect	319	292	320	293
rect	319	301	320	302
rect	319	304	320	305
rect	319	307	320	308
rect	319	313	320	314
rect	319	319	320	320
rect	319	322	320	323
rect	319	340	320	341
rect	319	343	320	344
rect	319	349	320	350
rect	319	352	320	353
rect	319	358	320	359
rect	319	361	320	362
rect	319	364	320	365
rect	320	13	321	14
rect	320	16	321	17
rect	320	19	321	20
rect	320	22	321	23
rect	320	28	321	29
rect	320	31	321	32
rect	320	34	321	35
rect	320	37	321	38
rect	320	46	321	47
rect	320	49	321	50
rect	320	58	321	59
rect	320	67	321	68
rect	320	70	321	71
rect	320	73	321	74
rect	320	76	321	77
rect	320	79	321	80
rect	320	82	321	83
rect	320	85	321	86
rect	320	88	321	89
rect	320	94	321	95
rect	320	97	321	98
rect	320	100	321	101
rect	320	103	321	104
rect	320	109	321	110
rect	320	121	321	122
rect	320	127	321	128
rect	320	130	321	131
rect	320	133	321	134
rect	320	136	321	137
rect	320	139	321	140
rect	320	142	321	143
rect	320	154	321	155
rect	320	157	321	158
rect	320	160	321	161
rect	320	166	321	167
rect	320	175	321	176
rect	320	178	321	179
rect	320	181	321	182
rect	320	184	321	185
rect	320	190	321	191
rect	320	196	321	197
rect	320	205	321	206
rect	320	208	321	209
rect	320	211	321	212
rect	320	214	321	215
rect	320	220	321	221
rect	320	223	321	224
rect	320	226	321	227
rect	320	229	321	230
rect	320	232	321	233
rect	320	235	321	236
rect	320	238	321	239
rect	320	241	321	242
rect	320	247	321	248
rect	320	250	321	251
rect	320	253	321	254
rect	320	259	321	260
rect	320	262	321	263
rect	320	268	321	269
rect	320	271	321	272
rect	320	274	321	275
rect	320	280	321	281
rect	320	283	321	284
rect	320	286	321	287
rect	320	289	321	290
rect	320	292	321	293
rect	320	301	321	302
rect	320	304	321	305
rect	320	307	321	308
rect	320	313	321	314
rect	320	319	321	320
rect	320	322	321	323
rect	320	331	321	332
rect	320	340	321	341
rect	320	343	321	344
rect	320	349	321	350
rect	320	352	321	353
rect	320	358	321	359
rect	320	361	321	362
rect	320	364	321	365
rect	321	13	322	14
rect	321	16	322	17
rect	321	22	322	23
rect	321	28	322	29
rect	321	31	322	32
rect	321	34	322	35
rect	321	37	322	38
rect	321	46	322	47
rect	321	49	322	50
rect	321	58	322	59
rect	321	67	322	68
rect	321	70	322	71
rect	321	73	322	74
rect	321	76	322	77
rect	321	79	322	80
rect	321	82	322	83
rect	321	85	322	86
rect	321	88	322	89
rect	321	94	322	95
rect	321	97	322	98
rect	321	100	322	101
rect	321	103	322	104
rect	321	109	322	110
rect	321	121	322	122
rect	321	127	322	128
rect	321	130	322	131
rect	321	133	322	134
rect	321	139	322	140
rect	321	142	322	143
rect	321	154	322	155
rect	321	157	322	158
rect	321	160	322	161
rect	321	166	322	167
rect	321	175	322	176
rect	321	178	322	179
rect	321	181	322	182
rect	321	184	322	185
rect	321	190	322	191
rect	321	196	322	197
rect	321	205	322	206
rect	321	208	322	209
rect	321	211	322	212
rect	321	214	322	215
rect	321	220	322	221
rect	321	223	322	224
rect	321	226	322	227
rect	321	229	322	230
rect	321	232	322	233
rect	321	235	322	236
rect	321	238	322	239
rect	321	241	322	242
rect	321	247	322	248
rect	321	250	322	251
rect	321	253	322	254
rect	321	259	322	260
rect	321	262	322	263
rect	321	268	322	269
rect	321	271	322	272
rect	321	283	322	284
rect	321	286	322	287
rect	321	289	322	290
rect	321	292	322	293
rect	321	301	322	302
rect	321	304	322	305
rect	321	307	322	308
rect	321	313	322	314
rect	321	319	322	320
rect	321	322	322	323
rect	321	331	322	332
rect	321	340	322	341
rect	321	343	322	344
rect	321	349	322	350
rect	321	352	322	353
rect	321	358	322	359
rect	321	361	322	362
rect	321	364	322	365
rect	322	11	323	12
rect	322	13	323	14
rect	322	16	323	17
rect	322	22	323	23
rect	322	28	323	29
rect	322	31	323	32
rect	322	34	323	35
rect	322	37	323	38
rect	322	46	323	47
rect	322	49	323	50
rect	322	58	323	59
rect	322	67	323	68
rect	322	70	323	71
rect	322	73	323	74
rect	322	76	323	77
rect	322	79	323	80
rect	322	82	323	83
rect	322	85	323	86
rect	322	88	323	89
rect	322	94	323	95
rect	322	97	323	98
rect	322	100	323	101
rect	322	103	323	104
rect	322	106	323	107
rect	322	109	323	110
rect	322	121	323	122
rect	322	127	323	128
rect	322	130	323	131
rect	322	133	323	134
rect	322	139	323	140
rect	322	142	323	143
rect	322	145	323	146
rect	322	154	323	155
rect	322	157	323	158
rect	322	160	323	161
rect	322	166	323	167
rect	322	175	323	176
rect	322	178	323	179
rect	322	181	323	182
rect	322	184	323	185
rect	322	190	323	191
rect	322	196	323	197
rect	322	205	323	206
rect	322	208	323	209
rect	322	211	323	212
rect	322	214	323	215
rect	322	220	323	221
rect	322	223	323	224
rect	322	226	323	227
rect	322	229	323	230
rect	322	232	323	233
rect	322	235	323	236
rect	322	238	323	239
rect	322	241	323	242
rect	322	247	323	248
rect	322	250	323	251
rect	322	253	323	254
rect	322	259	323	260
rect	322	262	323	263
rect	322	268	323	269
rect	322	271	323	272
rect	322	283	323	284
rect	322	286	323	287
rect	322	289	323	290
rect	322	292	323	293
rect	322	301	323	302
rect	322	304	323	305
rect	322	307	323	308
rect	322	313	323	314
rect	322	316	323	317
rect	322	319	323	320
rect	322	322	323	323
rect	322	331	323	332
rect	322	340	323	341
rect	322	343	323	344
rect	322	349	323	350
rect	322	352	323	353
rect	322	358	323	359
rect	322	361	323	362
rect	322	364	323	365
rect	323	11	324	12
rect	323	13	324	14
rect	323	22	324	23
rect	323	28	324	29
rect	323	31	324	32
rect	323	34	324	35
rect	323	37	324	38
rect	323	46	324	47
rect	323	49	324	50
rect	323	58	324	59
rect	323	67	324	68
rect	323	70	324	71
rect	323	73	324	74
rect	323	76	324	77
rect	323	82	324	83
rect	323	85	324	86
rect	323	88	324	89
rect	323	94	324	95
rect	323	97	324	98
rect	323	100	324	101
rect	323	103	324	104
rect	323	106	324	107
rect	323	109	324	110
rect	323	121	324	122
rect	323	127	324	128
rect	323	130	324	131
rect	323	133	324	134
rect	323	139	324	140
rect	323	142	324	143
rect	323	145	324	146
rect	323	154	324	155
rect	323	157	324	158
rect	323	160	324	161
rect	323	166	324	167
rect	323	175	324	176
rect	323	178	324	179
rect	323	181	324	182
rect	323	184	324	185
rect	323	190	324	191
rect	323	196	324	197
rect	323	205	324	206
rect	323	208	324	209
rect	323	211	324	212
rect	323	214	324	215
rect	323	220	324	221
rect	323	223	324	224
rect	323	226	324	227
rect	323	229	324	230
rect	323	232	324	233
rect	323	235	324	236
rect	323	238	324	239
rect	323	241	324	242
rect	323	247	324	248
rect	323	250	324	251
rect	323	253	324	254
rect	323	259	324	260
rect	323	262	324	263
rect	323	268	324	269
rect	323	271	324	272
rect	323	283	324	284
rect	323	286	324	287
rect	323	289	324	290
rect	323	292	324	293
rect	323	304	324	305
rect	323	307	324	308
rect	323	313	324	314
rect	323	316	324	317
rect	323	319	324	320
rect	323	322	324	323
rect	323	331	324	332
rect	323	340	324	341
rect	323	343	324	344
rect	323	349	324	350
rect	323	352	324	353
rect	323	358	324	359
rect	323	361	324	362
rect	323	364	324	365
rect	324	11	325	12
rect	324	13	325	14
rect	324	22	325	23
rect	324	25	325	26
rect	324	28	325	29
rect	324	31	325	32
rect	324	34	325	35
rect	324	37	325	38
rect	324	46	325	47
rect	324	49	325	50
rect	324	58	325	59
rect	324	67	325	68
rect	324	70	325	71
rect	324	73	325	74
rect	324	76	325	77
rect	324	82	325	83
rect	324	85	325	86
rect	324	88	325	89
rect	324	94	325	95
rect	324	97	325	98
rect	324	100	325	101
rect	324	103	325	104
rect	324	106	325	107
rect	324	109	325	110
rect	324	121	325	122
rect	324	127	325	128
rect	324	130	325	131
rect	324	133	325	134
rect	324	139	325	140
rect	324	142	325	143
rect	324	145	325	146
rect	324	154	325	155
rect	324	157	325	158
rect	324	160	325	161
rect	324	166	325	167
rect	324	175	325	176
rect	324	178	325	179
rect	324	181	325	182
rect	324	184	325	185
rect	324	190	325	191
rect	324	196	325	197
rect	324	205	325	206
rect	324	208	325	209
rect	324	211	325	212
rect	324	214	325	215
rect	324	220	325	221
rect	324	223	325	224
rect	324	226	325	227
rect	324	229	325	230
rect	324	232	325	233
rect	324	235	325	236
rect	324	238	325	239
rect	324	241	325	242
rect	324	247	325	248
rect	324	250	325	251
rect	324	253	325	254
rect	324	259	325	260
rect	324	262	325	263
rect	324	268	325	269
rect	324	271	325	272
rect	324	280	325	281
rect	324	283	325	284
rect	324	286	325	287
rect	324	289	325	290
rect	324	292	325	293
rect	324	304	325	305
rect	324	307	325	308
rect	324	310	325	311
rect	324	313	325	314
rect	324	316	325	317
rect	324	319	325	320
rect	324	322	325	323
rect	324	331	325	332
rect	324	340	325	341
rect	324	343	325	344
rect	324	349	325	350
rect	324	352	325	353
rect	324	358	325	359
rect	324	361	325	362
rect	324	364	325	365
rect	325	11	326	12
rect	325	13	326	14
rect	325	22	326	23
rect	325	25	326	26
rect	325	28	326	29
rect	325	34	326	35
rect	325	37	326	38
rect	325	46	326	47
rect	325	49	326	50
rect	325	58	326	59
rect	325	67	326	68
rect	325	70	326	71
rect	325	73	326	74
rect	325	76	326	77
rect	325	85	326	86
rect	325	88	326	89
rect	325	94	326	95
rect	325	100	326	101
rect	325	103	326	104
rect	325	106	326	107
rect	325	109	326	110
rect	325	121	326	122
rect	325	127	326	128
rect	325	130	326	131
rect	325	133	326	134
rect	325	142	326	143
rect	325	145	326	146
rect	325	157	326	158
rect	325	160	326	161
rect	325	166	326	167
rect	325	175	326	176
rect	325	178	326	179
rect	325	181	326	182
rect	325	184	326	185
rect	325	190	326	191
rect	325	196	326	197
rect	325	205	326	206
rect	325	208	326	209
rect	325	211	326	212
rect	325	214	326	215
rect	325	220	326	221
rect	325	226	326	227
rect	325	229	326	230
rect	325	232	326	233
rect	325	238	326	239
rect	325	241	326	242
rect	325	250	326	251
rect	325	253	326	254
rect	325	259	326	260
rect	325	262	326	263
rect	325	268	326	269
rect	325	280	326	281
rect	325	283	326	284
rect	325	286	326	287
rect	325	289	326	290
rect	325	304	326	305
rect	325	310	326	311
rect	325	316	326	317
rect	325	319	326	320
rect	325	322	326	323
rect	325	331	326	332
rect	325	340	326	341
rect	325	343	326	344
rect	325	352	326	353
rect	325	358	326	359
rect	325	361	326	362
rect	325	364	326	365
rect	326	11	327	12
rect	326	13	327	14
rect	326	16	327	17
rect	326	22	327	23
rect	326	25	327	26
rect	326	28	327	29
rect	326	34	327	35
rect	326	37	327	38
rect	326	46	327	47
rect	326	49	327	50
rect	326	58	327	59
rect	326	61	327	62
rect	326	67	327	68
rect	326	70	327	71
rect	326	73	327	74
rect	326	76	327	77
rect	326	85	327	86
rect	326	88	327	89
rect	326	94	327	95
rect	326	100	327	101
rect	326	103	327	104
rect	326	106	327	107
rect	326	109	327	110
rect	326	121	327	122
rect	326	124	327	125
rect	326	127	327	128
rect	326	130	327	131
rect	326	133	327	134
rect	326	136	327	137
rect	326	142	327	143
rect	326	145	327	146
rect	326	148	327	149
rect	326	157	327	158
rect	326	160	327	161
rect	326	163	327	164
rect	326	166	327	167
rect	326	175	327	176
rect	326	178	327	179
rect	326	181	327	182
rect	326	184	327	185
rect	326	190	327	191
rect	326	196	327	197
rect	326	205	327	206
rect	326	208	327	209
rect	326	211	327	212
rect	326	214	327	215
rect	326	220	327	221
rect	326	226	327	227
rect	326	229	327	230
rect	326	232	327	233
rect	326	238	327	239
rect	326	241	327	242
rect	326	244	327	245
rect	326	250	327	251
rect	326	253	327	254
rect	326	259	327	260
rect	326	262	327	263
rect	326	265	327	266
rect	326	268	327	269
rect	326	274	327	275
rect	326	280	327	281
rect	326	283	327	284
rect	326	286	327	287
rect	326	289	327	290
rect	326	301	327	302
rect	326	304	327	305
rect	326	310	327	311
rect	326	316	327	317
rect	326	319	327	320
rect	326	322	327	323
rect	326	331	327	332
rect	326	340	327	341
rect	326	343	327	344
rect	326	352	327	353
rect	326	358	327	359
rect	326	361	327	362
rect	326	364	327	365
rect	326	373	327	374
rect	327	11	328	12
rect	327	16	328	17
rect	327	22	328	23
rect	327	25	328	26
rect	327	28	328	29
rect	327	34	328	35
rect	327	37	328	38
rect	327	46	328	47
rect	327	49	328	50
rect	327	61	328	62
rect	327	67	328	68
rect	327	70	328	71
rect	327	76	328	77
rect	327	85	328	86
rect	327	88	328	89
rect	327	100	328	101
rect	327	103	328	104
rect	327	106	328	107
rect	327	109	328	110
rect	327	121	328	122
rect	327	124	328	125
rect	327	127	328	128
rect	327	130	328	131
rect	327	136	328	137
rect	327	142	328	143
rect	327	145	328	146
rect	327	148	328	149
rect	327	157	328	158
rect	327	160	328	161
rect	327	163	328	164
rect	327	166	328	167
rect	327	175	328	176
rect	327	178	328	179
rect	327	181	328	182
rect	327	184	328	185
rect	327	196	328	197
rect	327	205	328	206
rect	327	208	328	209
rect	327	211	328	212
rect	327	220	328	221
rect	327	226	328	227
rect	327	229	328	230
rect	327	238	328	239
rect	327	241	328	242
rect	327	244	328	245
rect	327	250	328	251
rect	327	253	328	254
rect	327	259	328	260
rect	327	265	328	266
rect	327	268	328	269
rect	327	274	328	275
rect	327	280	328	281
rect	327	286	328	287
rect	327	289	328	290
rect	327	301	328	302
rect	327	304	328	305
rect	327	310	328	311
rect	327	316	328	317
rect	327	319	328	320
rect	327	322	328	323
rect	327	331	328	332
rect	327	343	328	344
rect	327	352	328	353
rect	327	358	328	359
rect	327	361	328	362
rect	327	364	328	365
rect	327	373	328	374
rect	328	11	329	12
rect	328	16	329	17
rect	328	19	329	20
rect	328	22	329	23
rect	328	25	329	26
rect	328	28	329	29
rect	328	34	329	35
rect	328	37	329	38
rect	328	46	329	47
rect	328	49	329	50
rect	328	61	329	62
rect	328	64	329	65
rect	328	67	329	68
rect	328	70	329	71
rect	328	76	329	77
rect	328	79	329	80
rect	328	85	329	86
rect	328	88	329	89
rect	328	91	329	92
rect	328	97	329	98
rect	328	100	329	101
rect	328	103	329	104
rect	328	106	329	107
rect	328	109	329	110
rect	328	121	329	122
rect	328	124	329	125
rect	328	127	329	128
rect	328	130	329	131
rect	328	136	329	137
rect	328	139	329	140
rect	328	142	329	143
rect	328	145	329	146
rect	328	148	329	149
rect	328	157	329	158
rect	328	160	329	161
rect	328	163	329	164
rect	328	166	329	167
rect	328	175	329	176
rect	328	178	329	179
rect	328	181	329	182
rect	328	184	329	185
rect	328	187	329	188
rect	328	193	329	194
rect	328	196	329	197
rect	328	205	329	206
rect	328	208	329	209
rect	328	211	329	212
rect	328	220	329	221
rect	328	223	329	224
rect	328	226	329	227
rect	328	229	329	230
rect	328	238	329	239
rect	328	241	329	242
rect	328	244	329	245
rect	328	250	329	251
rect	328	253	329	254
rect	328	256	329	257
rect	328	259	329	260
rect	328	265	329	266
rect	328	268	329	269
rect	328	271	329	272
rect	328	274	329	275
rect	328	280	329	281
rect	328	286	329	287
rect	328	289	329	290
rect	328	301	329	302
rect	328	304	329	305
rect	328	310	329	311
rect	328	313	329	314
rect	328	316	329	317
rect	328	319	329	320
rect	328	322	329	323
rect	328	331	329	332
rect	328	343	329	344
rect	328	349	329	350
rect	328	352	329	353
rect	328	358	329	359
rect	328	361	329	362
rect	328	364	329	365
rect	328	373	329	374
rect	329	11	330	12
rect	329	16	330	17
rect	329	19	330	20
rect	329	22	330	23
rect	329	25	330	26
rect	329	34	330	35
rect	329	37	330	38
rect	329	46	330	47
rect	329	61	330	62
rect	329	64	330	65
rect	329	67	330	68
rect	329	70	330	71
rect	329	79	330	80
rect	329	85	330	86
rect	329	91	330	92
rect	329	97	330	98
rect	329	100	330	101
rect	329	103	330	104
rect	329	106	330	107
rect	329	109	330	110
rect	329	121	330	122
rect	329	124	330	125
rect	329	127	330	128
rect	329	130	330	131
rect	329	136	330	137
rect	329	139	330	140
rect	329	142	330	143
rect	329	145	330	146
rect	329	148	330	149
rect	329	157	330	158
rect	329	160	330	161
rect	329	163	330	164
rect	329	166	330	167
rect	329	175	330	176
rect	329	178	330	179
rect	329	181	330	182
rect	329	184	330	185
rect	329	187	330	188
rect	329	193	330	194
rect	329	196	330	197
rect	329	205	330	206
rect	329	208	330	209
rect	329	211	330	212
rect	329	220	330	221
rect	329	223	330	224
rect	329	226	330	227
rect	329	229	330	230
rect	329	238	330	239
rect	329	241	330	242
rect	329	244	330	245
rect	329	250	330	251
rect	329	253	330	254
rect	329	256	330	257
rect	329	259	330	260
rect	329	265	330	266
rect	329	268	330	269
rect	329	271	330	272
rect	329	274	330	275
rect	329	280	330	281
rect	329	286	330	287
rect	329	289	330	290
rect	329	301	330	302
rect	329	304	330	305
rect	329	310	330	311
rect	329	313	330	314
rect	329	316	330	317
rect	329	319	330	320
rect	329	322	330	323
rect	329	331	330	332
rect	329	343	330	344
rect	329	349	330	350
rect	329	352	330	353
rect	329	358	330	359
rect	329	361	330	362
rect	329	364	330	365
rect	329	373	330	374
rect	330	11	331	12
rect	330	13	331	14
rect	330	16	331	17
rect	330	19	331	20
rect	330	22	331	23
rect	330	25	331	26
rect	330	34	331	35
rect	330	37	331	38
rect	330	44	331	45
rect	330	46	331	47
rect	330	58	331	59
rect	330	61	331	62
rect	330	64	331	65
rect	330	67	331	68
rect	330	70	331	71
rect	330	79	331	80
rect	330	85	331	86
rect	330	91	331	92
rect	330	94	331	95
rect	330	97	331	98
rect	330	100	331	101
rect	330	103	331	104
rect	330	106	331	107
rect	330	109	331	110
rect	330	115	331	116
rect	330	118	331	119
rect	330	121	331	122
rect	330	124	331	125
rect	330	127	331	128
rect	330	130	331	131
rect	330	133	331	134
rect	330	136	331	137
rect	330	139	331	140
rect	330	142	331	143
rect	330	145	331	146
rect	330	148	331	149
rect	330	157	331	158
rect	330	160	331	161
rect	330	163	331	164
rect	330	166	331	167
rect	330	175	331	176
rect	330	178	331	179
rect	330	181	331	182
rect	330	184	331	185
rect	330	187	331	188
rect	330	193	331	194
rect	330	196	331	197
rect	330	205	331	206
rect	330	208	331	209
rect	330	211	331	212
rect	330	220	331	221
rect	330	223	331	224
rect	330	226	331	227
rect	330	229	331	230
rect	330	238	331	239
rect	330	241	331	242
rect	330	244	331	245
rect	330	250	331	251
rect	330	253	331	254
rect	330	256	331	257
rect	330	259	331	260
rect	330	265	331	266
rect	330	268	331	269
rect	330	271	331	272
rect	330	274	331	275
rect	330	280	331	281
rect	330	286	331	287
rect	330	289	331	290
rect	330	301	331	302
rect	330	304	331	305
rect	330	310	331	311
rect	330	313	331	314
rect	330	316	331	317
rect	330	319	331	320
rect	330	322	331	323
rect	330	331	331	332
rect	330	343	331	344
rect	330	346	331	347
rect	330	349	331	350
rect	330	352	331	353
rect	330	358	331	359
rect	330	361	331	362
rect	330	364	331	365
rect	330	373	331	374
rect	331	13	332	14
rect	331	16	332	17
rect	331	19	332	20
rect	331	22	332	23
rect	331	25	332	26
rect	331	37	332	38
rect	331	44	332	45
rect	331	58	332	59
rect	331	61	332	62
rect	331	64	332	65
rect	331	67	332	68
rect	331	79	332	80
rect	331	91	332	92
rect	331	94	332	95
rect	331	97	332	98
rect	331	100	332	101
rect	331	103	332	104
rect	331	106	332	107
rect	331	109	332	110
rect	331	115	332	116
rect	331	118	332	119
rect	331	121	332	122
rect	331	124	332	125
rect	331	127	332	128
rect	331	130	332	131
rect	331	133	332	134
rect	331	136	332	137
rect	331	139	332	140
rect	331	142	332	143
rect	331	145	332	146
rect	331	148	332	149
rect	331	157	332	158
rect	331	160	332	161
rect	331	163	332	164
rect	331	166	332	167
rect	331	175	332	176
rect	331	178	332	179
rect	331	181	332	182
rect	331	184	332	185
rect	331	187	332	188
rect	331	193	332	194
rect	331	196	332	197
rect	331	205	332	206
rect	331	208	332	209
rect	331	211	332	212
rect	331	220	332	221
rect	331	223	332	224
rect	331	226	332	227
rect	331	229	332	230
rect	331	238	332	239
rect	331	241	332	242
rect	331	244	332	245
rect	331	250	332	251
rect	331	253	332	254
rect	331	256	332	257
rect	331	259	332	260
rect	331	265	332	266
rect	331	268	332	269
rect	331	271	332	272
rect	331	274	332	275
rect	331	280	332	281
rect	331	286	332	287
rect	331	289	332	290
rect	331	301	332	302
rect	331	304	332	305
rect	331	310	332	311
rect	331	313	332	314
rect	331	316	332	317
rect	331	322	332	323
rect	331	331	332	332
rect	331	343	332	344
rect	331	346	332	347
rect	331	349	332	350
rect	331	352	332	353
rect	331	358	332	359
rect	331	361	332	362
rect	331	373	332	374
rect	332	13	333	14
rect	332	16	333	17
rect	332	19	333	20
rect	332	22	333	23
rect	332	25	333	26
rect	332	28	333	29
rect	332	31	333	32
rect	332	37	333	38
rect	332	44	333	45
rect	332	49	333	50
rect	332	58	333	59
rect	332	61	333	62
rect	332	64	333	65
rect	332	67	333	68
rect	332	76	333	77
rect	332	79	333	80
rect	332	82	333	83
rect	332	88	333	89
rect	332	91	333	92
rect	332	94	333	95
rect	332	97	333	98
rect	332	100	333	101
rect	332	103	333	104
rect	332	106	333	107
rect	332	109	333	110
rect	332	115	333	116
rect	332	118	333	119
rect	332	121	333	122
rect	332	124	333	125
rect	332	127	333	128
rect	332	130	333	131
rect	332	133	333	134
rect	332	136	333	137
rect	332	139	333	140
rect	332	142	333	143
rect	332	145	333	146
rect	332	148	333	149
rect	332	157	333	158
rect	332	160	333	161
rect	332	163	333	164
rect	332	166	333	167
rect	332	175	333	176
rect	332	178	333	179
rect	332	181	333	182
rect	332	184	333	185
rect	332	187	333	188
rect	332	193	333	194
rect	332	196	333	197
rect	332	205	333	206
rect	332	208	333	209
rect	332	211	333	212
rect	332	220	333	221
rect	332	223	333	224
rect	332	226	333	227
rect	332	229	333	230
rect	332	238	333	239
rect	332	241	333	242
rect	332	244	333	245
rect	332	250	333	251
rect	332	253	333	254
rect	332	256	333	257
rect	332	259	333	260
rect	332	265	333	266
rect	332	268	333	269
rect	332	271	333	272
rect	332	274	333	275
rect	332	280	333	281
rect	332	286	333	287
rect	332	289	333	290
rect	332	295	333	296
rect	332	301	333	302
rect	332	304	333	305
rect	332	310	333	311
rect	332	313	333	314
rect	332	316	333	317
rect	332	322	333	323
rect	332	331	333	332
rect	332	340	333	341
rect	332	343	333	344
rect	332	346	333	347
rect	332	349	333	350
rect	332	352	333	353
rect	332	358	333	359
rect	332	361	333	362
rect	332	373	333	374
rect	332	376	333	377
rect	333	13	334	14
rect	333	16	334	17
rect	333	19	334	20
rect	333	25	334	26
rect	333	28	334	29
rect	333	31	334	32
rect	333	37	334	38
rect	333	49	334	50
rect	333	58	334	59
rect	333	61	334	62
rect	333	64	334	65
rect	333	76	334	77
rect	333	79	334	80
rect	333	82	334	83
rect	333	88	334	89
rect	333	91	334	92
rect	333	94	334	95
rect	333	97	334	98
rect	333	100	334	101
rect	333	103	334	104
rect	333	106	334	107
rect	333	109	334	110
rect	333	115	334	116
rect	333	118	334	119
rect	333	121	334	122
rect	333	124	334	125
rect	333	127	334	128
rect	333	130	334	131
rect	333	133	334	134
rect	333	136	334	137
rect	333	139	334	140
rect	333	142	334	143
rect	333	145	334	146
rect	333	148	334	149
rect	333	157	334	158
rect	333	160	334	161
rect	333	163	334	164
rect	333	166	334	167
rect	333	175	334	176
rect	333	178	334	179
rect	333	181	334	182
rect	333	184	334	185
rect	333	187	334	188
rect	333	193	334	194
rect	333	196	334	197
rect	333	205	334	206
rect	333	208	334	209
rect	333	211	334	212
rect	333	220	334	221
rect	333	223	334	224
rect	333	226	334	227
rect	333	229	334	230
rect	333	238	334	239
rect	333	241	334	242
rect	333	244	334	245
rect	333	253	334	254
rect	333	256	334	257
rect	333	265	334	266
rect	333	268	334	269
rect	333	271	334	272
rect	333	274	334	275
rect	333	280	334	281
rect	333	286	334	287
rect	333	295	334	296
rect	333	301	334	302
rect	333	310	334	311
rect	333	313	334	314
rect	333	316	334	317
rect	333	322	334	323
rect	333	331	334	332
rect	333	340	334	341
rect	333	343	334	344
rect	333	346	334	347
rect	333	349	334	350
rect	333	358	334	359
rect	333	361	334	362
rect	333	373	334	374
rect	333	376	334	377
rect	334	13	335	14
rect	334	16	335	17
rect	334	19	335	20
rect	334	25	335	26
rect	334	28	335	29
rect	334	31	335	32
rect	334	34	335	35
rect	334	37	335	38
rect	334	46	335	47
rect	334	49	335	50
rect	334	58	335	59
rect	334	61	335	62
rect	334	64	335	65
rect	334	73	335	74
rect	334	76	335	77
rect	334	79	335	80
rect	334	82	335	83
rect	334	85	335	86
rect	334	88	335	89
rect	334	91	335	92
rect	334	94	335	95
rect	334	97	335	98
rect	334	100	335	101
rect	334	103	335	104
rect	334	106	335	107
rect	334	109	335	110
rect	334	115	335	116
rect	334	118	335	119
rect	334	121	335	122
rect	334	124	335	125
rect	334	127	335	128
rect	334	130	335	131
rect	334	133	335	134
rect	334	136	335	137
rect	334	139	335	140
rect	334	142	335	143
rect	334	145	335	146
rect	334	148	335	149
rect	334	157	335	158
rect	334	160	335	161
rect	334	163	335	164
rect	334	166	335	167
rect	334	175	335	176
rect	334	178	335	179
rect	334	181	335	182
rect	334	184	335	185
rect	334	187	335	188
rect	334	193	335	194
rect	334	196	335	197
rect	334	205	335	206
rect	334	208	335	209
rect	334	211	335	212
rect	334	220	335	221
rect	334	223	335	224
rect	334	226	335	227
rect	334	229	335	230
rect	334	238	335	239
rect	334	241	335	242
rect	334	244	335	245
rect	334	253	335	254
rect	334	256	335	257
rect	334	265	335	266
rect	334	268	335	269
rect	334	271	335	272
rect	334	274	335	275
rect	334	280	335	281
rect	334	283	335	284
rect	334	286	335	287
rect	334	295	335	296
rect	334	298	335	299
rect	334	301	335	302
rect	334	310	335	311
rect	334	313	335	314
rect	334	316	335	317
rect	334	319	335	320
rect	334	322	335	323
rect	334	331	335	332
rect	334	340	335	341
rect	334	343	335	344
rect	334	346	335	347
rect	334	349	335	350
rect	334	358	335	359
rect	334	361	335	362
rect	334	364	335	365
rect	334	373	335	374
rect	334	376	335	377
rect	335	13	336	14
rect	335	16	336	17
rect	335	19	336	20
rect	335	25	336	26
rect	335	28	336	29
rect	335	31	336	32
rect	335	34	336	35
rect	335	37	336	38
rect	335	46	336	47
rect	335	49	336	50
rect	335	58	336	59
rect	335	61	336	62
rect	335	64	336	65
rect	335	73	336	74
rect	335	76	336	77
rect	335	79	336	80
rect	335	82	336	83
rect	335	85	336	86
rect	335	88	336	89
rect	335	91	336	92
rect	335	94	336	95
rect	335	97	336	98
rect	335	100	336	101
rect	335	103	336	104
rect	335	106	336	107
rect	335	109	336	110
rect	335	115	336	116
rect	335	118	336	119
rect	335	121	336	122
rect	335	124	336	125
rect	335	127	336	128
rect	335	130	336	131
rect	335	133	336	134
rect	335	136	336	137
rect	335	139	336	140
rect	335	142	336	143
rect	335	145	336	146
rect	335	148	336	149
rect	335	157	336	158
rect	335	160	336	161
rect	335	163	336	164
rect	335	166	336	167
rect	335	175	336	176
rect	335	178	336	179
rect	335	181	336	182
rect	335	184	336	185
rect	335	187	336	188
rect	335	193	336	194
rect	335	196	336	197
rect	335	205	336	206
rect	335	208	336	209
rect	335	211	336	212
rect	335	220	336	221
rect	335	223	336	224
rect	335	226	336	227
rect	335	229	336	230
rect	335	238	336	239
rect	335	241	336	242
rect	335	244	336	245
rect	335	253	336	254
rect	335	256	336	257
rect	335	265	336	266
rect	335	268	336	269
rect	335	271	336	272
rect	335	274	336	275
rect	335	280	336	281
rect	335	283	336	284
rect	335	286	336	287
rect	335	295	336	296
rect	335	298	336	299
rect	335	301	336	302
rect	335	310	336	311
rect	335	313	336	314
rect	335	316	336	317
rect	335	319	336	320
rect	335	322	336	323
rect	335	331	336	332
rect	335	340	336	341
rect	335	343	336	344
rect	335	346	336	347
rect	335	349	336	350
rect	335	364	336	365
rect	335	373	336	374
rect	335	376	336	377
rect	336	13	337	14
rect	336	16	337	17
rect	336	19	337	20
rect	336	22	337	23
rect	336	25	337	26
rect	336	28	337	29
rect	336	31	337	32
rect	336	34	337	35
rect	336	37	337	38
rect	336	46	337	47
rect	336	49	337	50
rect	336	58	337	59
rect	336	61	337	62
rect	336	64	337	65
rect	336	73	337	74
rect	336	76	337	77
rect	336	79	337	80
rect	336	82	337	83
rect	336	85	337	86
rect	336	88	337	89
rect	336	91	337	92
rect	336	94	337	95
rect	336	97	337	98
rect	336	100	337	101
rect	336	103	337	104
rect	336	106	337	107
rect	336	109	337	110
rect	336	115	337	116
rect	336	118	337	119
rect	336	121	337	122
rect	336	124	337	125
rect	336	127	337	128
rect	336	130	337	131
rect	336	133	337	134
rect	336	136	337	137
rect	336	139	337	140
rect	336	142	337	143
rect	336	145	337	146
rect	336	148	337	149
rect	336	157	337	158
rect	336	160	337	161
rect	336	163	337	164
rect	336	166	337	167
rect	336	175	337	176
rect	336	178	337	179
rect	336	181	337	182
rect	336	184	337	185
rect	336	187	337	188
rect	336	193	337	194
rect	336	196	337	197
rect	336	205	337	206
rect	336	208	337	209
rect	336	211	337	212
rect	336	220	337	221
rect	336	223	337	224
rect	336	226	337	227
rect	336	229	337	230
rect	336	238	337	239
rect	336	241	337	242
rect	336	244	337	245
rect	336	253	337	254
rect	336	256	337	257
rect	336	265	337	266
rect	336	268	337	269
rect	336	271	337	272
rect	336	274	337	275
rect	336	280	337	281
rect	336	283	337	284
rect	336	286	337	287
rect	336	295	337	296
rect	336	298	337	299
rect	336	301	337	302
rect	336	310	337	311
rect	336	313	337	314
rect	336	316	337	317
rect	336	319	337	320
rect	336	322	337	323
rect	336	331	337	332
rect	336	340	337	341
rect	336	343	337	344
rect	336	346	337	347
rect	336	349	337	350
rect	336	364	337	365
rect	336	373	337	374
rect	336	376	337	377
rect	336	385	337	386
rect	343	10	344	11
rect	343	13	344	14
rect	343	16	344	17
rect	343	19	344	20
rect	343	22	344	23
rect	343	25	344	26
rect	343	28	344	29
rect	343	31	344	32
rect	343	34	344	35
rect	343	37	344	38
rect	343	43	344	44
rect	343	46	344	47
rect	343	49	344	50
rect	343	58	344	59
rect	343	61	344	62
rect	343	64	344	65
rect	343	73	344	74
rect	343	76	344	77
rect	343	79	344	80
rect	343	82	344	83
rect	343	91	344	92
rect	343	94	344	95
rect	343	97	344	98
rect	343	100	344	101
rect	343	103	344	104
rect	343	106	344	107
rect	343	109	344	110
rect	343	118	344	119
rect	343	121	344	122
rect	343	124	344	125
rect	343	127	344	128
rect	343	130	344	131
rect	343	133	344	134
rect	343	136	344	137
rect	343	139	344	140
rect	343	142	344	143
rect	343	145	344	146
rect	343	148	344	149
rect	343	157	344	158
rect	343	160	344	161
rect	343	163	344	164
rect	343	166	344	167
rect	343	169	344	170
rect	343	175	344	176
rect	343	178	344	179
rect	343	181	344	182
rect	343	184	344	185
rect	343	190	344	191
rect	343	193	344	194
rect	343	196	344	197
rect	343	205	344	206
rect	343	208	344	209
rect	343	211	344	212
rect	343	220	344	221
rect	343	223	344	224
rect	343	226	344	227
rect	343	229	344	230
rect	343	238	344	239
rect	343	241	344	242
rect	343	244	344	245
rect	343	253	344	254
rect	343	256	344	257
rect	343	259	344	260
rect	343	265	344	266
rect	343	268	344	269
rect	343	271	344	272
rect	343	274	344	275
rect	343	280	344	281
rect	343	283	344	284
rect	343	286	344	287
rect	343	295	344	296
rect	343	298	344	299
rect	343	301	344	302
rect	343	310	344	311
rect	343	313	344	314
rect	343	316	344	317
rect	343	319	344	320
rect	343	322	344	323
rect	343	328	344	329
rect	343	331	344	332
rect	343	337	344	338
rect	343	340	344	341
rect	343	343	344	344
rect	343	349	344	350
rect	343	364	344	365
rect	343	370	344	371
rect	343	373	344	374
rect	343	376	344	377
rect	343	379	344	380
rect	343	385	344	386
rect	344	10	345	11
rect	344	13	345	14
rect	344	16	345	17
rect	344	19	345	20
rect	344	22	345	23
rect	344	25	345	26
rect	344	28	345	29
rect	344	31	345	32
rect	344	34	345	35
rect	344	37	345	38
rect	344	43	345	44
rect	344	46	345	47
rect	344	49	345	50
rect	344	58	345	59
rect	344	61	345	62
rect	344	64	345	65
rect	344	73	345	74
rect	344	76	345	77
rect	344	79	345	80
rect	344	82	345	83
rect	344	91	345	92
rect	344	94	345	95
rect	344	97	345	98
rect	344	100	345	101
rect	344	103	345	104
rect	344	106	345	107
rect	344	109	345	110
rect	344	118	345	119
rect	344	121	345	122
rect	344	124	345	125
rect	344	127	345	128
rect	344	130	345	131
rect	344	133	345	134
rect	344	136	345	137
rect	344	139	345	140
rect	344	142	345	143
rect	344	145	345	146
rect	344	148	345	149
rect	344	157	345	158
rect	344	160	345	161
rect	344	163	345	164
rect	344	166	345	167
rect	344	169	345	170
rect	344	175	345	176
rect	344	178	345	179
rect	344	181	345	182
rect	344	184	345	185
rect	344	190	345	191
rect	344	193	345	194
rect	344	196	345	197
rect	344	205	345	206
rect	344	208	345	209
rect	344	211	345	212
rect	344	220	345	221
rect	344	223	345	224
rect	344	226	345	227
rect	344	229	345	230
rect	344	238	345	239
rect	344	241	345	242
rect	344	244	345	245
rect	344	253	345	254
rect	344	256	345	257
rect	344	259	345	260
rect	344	265	345	266
rect	344	268	345	269
rect	344	271	345	272
rect	344	274	345	275
rect	344	280	345	281
rect	344	283	345	284
rect	344	286	345	287
rect	344	298	345	299
rect	344	301	345	302
rect	344	310	345	311
rect	344	313	345	314
rect	344	316	345	317
rect	344	319	345	320
rect	344	322	345	323
rect	344	328	345	329
rect	344	331	345	332
rect	344	337	345	338
rect	344	340	345	341
rect	344	343	345	344
rect	344	349	345	350
rect	344	364	345	365
rect	344	370	345	371
rect	344	373	345	374
rect	344	376	345	377
rect	344	379	345	380
rect	344	385	345	386
rect	345	10	346	11
rect	345	13	346	14
rect	345	16	346	17
rect	345	19	346	20
rect	345	22	346	23
rect	345	25	346	26
rect	345	28	346	29
rect	345	31	346	32
rect	345	34	346	35
rect	345	37	346	38
rect	345	43	346	44
rect	345	46	346	47
rect	345	49	346	50
rect	345	58	346	59
rect	345	61	346	62
rect	345	64	346	65
rect	345	73	346	74
rect	345	76	346	77
rect	345	79	346	80
rect	345	82	346	83
rect	345	91	346	92
rect	345	94	346	95
rect	345	97	346	98
rect	345	100	346	101
rect	345	103	346	104
rect	345	106	346	107
rect	345	109	346	110
rect	345	118	346	119
rect	345	121	346	122
rect	345	124	346	125
rect	345	127	346	128
rect	345	130	346	131
rect	345	133	346	134
rect	345	136	346	137
rect	345	139	346	140
rect	345	142	346	143
rect	345	145	346	146
rect	345	148	346	149
rect	345	157	346	158
rect	345	160	346	161
rect	345	163	346	164
rect	345	166	346	167
rect	345	169	346	170
rect	345	175	346	176
rect	345	178	346	179
rect	345	181	346	182
rect	345	184	346	185
rect	345	190	346	191
rect	345	193	346	194
rect	345	196	346	197
rect	345	205	346	206
rect	345	208	346	209
rect	345	211	346	212
rect	345	220	346	221
rect	345	223	346	224
rect	345	226	346	227
rect	345	229	346	230
rect	345	233	346	234
rect	345	238	346	239
rect	345	241	346	242
rect	345	244	346	245
rect	345	253	346	254
rect	345	256	346	257
rect	345	259	346	260
rect	345	265	346	266
rect	345	268	346	269
rect	345	271	346	272
rect	345	274	346	275
rect	345	280	346	281
rect	345	283	346	284
rect	345	286	346	287
rect	345	298	346	299
rect	345	301	346	302
rect	345	310	346	311
rect	345	313	346	314
rect	345	316	346	317
rect	345	319	346	320
rect	345	322	346	323
rect	345	328	346	329
rect	345	331	346	332
rect	345	337	346	338
rect	345	340	346	341
rect	345	343	346	344
rect	345	349	346	350
rect	345	364	346	365
rect	345	370	346	371
rect	345	373	346	374
rect	345	376	346	377
rect	345	379	346	380
rect	345	385	346	386
rect	346	10	347	11
rect	346	13	347	14
rect	346	16	347	17
rect	346	19	347	20
rect	346	22	347	23
rect	346	25	347	26
rect	346	28	347	29
rect	346	31	347	32
rect	346	34	347	35
rect	346	37	347	38
rect	346	43	347	44
rect	346	46	347	47
rect	346	49	347	50
rect	346	58	347	59
rect	346	61	347	62
rect	346	64	347	65
rect	346	73	347	74
rect	346	76	347	77
rect	346	79	347	80
rect	346	82	347	83
rect	346	91	347	92
rect	346	94	347	95
rect	346	97	347	98
rect	346	100	347	101
rect	346	103	347	104
rect	346	106	347	107
rect	346	109	347	110
rect	346	118	347	119
rect	346	121	347	122
rect	346	124	347	125
rect	346	127	347	128
rect	346	130	347	131
rect	346	133	347	134
rect	346	136	347	137
rect	346	139	347	140
rect	346	142	347	143
rect	346	145	347	146
rect	346	148	347	149
rect	346	157	347	158
rect	346	160	347	161
rect	346	163	347	164
rect	346	166	347	167
rect	346	169	347	170
rect	346	175	347	176
rect	346	178	347	179
rect	346	181	347	182
rect	346	184	347	185
rect	346	190	347	191
rect	346	193	347	194
rect	346	196	347	197
rect	346	205	347	206
rect	346	208	347	209
rect	346	211	347	212
rect	346	220	347	221
rect	346	223	347	224
rect	346	226	347	227
rect	346	229	347	230
rect	346	233	347	234
rect	346	238	347	239
rect	346	241	347	242
rect	346	244	347	245
rect	346	253	347	254
rect	346	256	347	257
rect	346	259	347	260
rect	346	265	347	266
rect	346	268	347	269
rect	346	271	347	272
rect	346	274	347	275
rect	346	280	347	281
rect	346	283	347	284
rect	346	286	347	287
rect	346	298	347	299
rect	346	301	347	302
rect	346	313	347	314
rect	346	316	347	317
rect	346	319	347	320
rect	346	322	347	323
rect	346	328	347	329
rect	346	331	347	332
rect	346	337	347	338
rect	346	340	347	341
rect	346	343	347	344
rect	346	349	347	350
rect	346	364	347	365
rect	346	370	347	371
rect	346	373	347	374
rect	346	376	347	377
rect	346	379	347	380
rect	346	385	347	386
rect	347	10	348	11
rect	347	13	348	14
rect	347	16	348	17
rect	347	19	348	20
rect	347	22	348	23
rect	347	25	348	26
rect	347	28	348	29
rect	347	31	348	32
rect	347	34	348	35
rect	347	37	348	38
rect	347	43	348	44
rect	347	46	348	47
rect	347	49	348	50
rect	347	58	348	59
rect	347	61	348	62
rect	347	64	348	65
rect	347	73	348	74
rect	347	76	348	77
rect	347	79	348	80
rect	347	82	348	83
rect	347	91	348	92
rect	347	94	348	95
rect	347	97	348	98
rect	347	100	348	101
rect	347	103	348	104
rect	347	106	348	107
rect	347	109	348	110
rect	347	118	348	119
rect	347	121	348	122
rect	347	124	348	125
rect	347	127	348	128
rect	347	130	348	131
rect	347	133	348	134
rect	347	136	348	137
rect	347	139	348	140
rect	347	142	348	143
rect	347	145	348	146
rect	347	148	348	149
rect	347	157	348	158
rect	347	160	348	161
rect	347	163	348	164
rect	347	166	348	167
rect	347	169	348	170
rect	347	175	348	176
rect	347	178	348	179
rect	347	181	348	182
rect	347	184	348	185
rect	347	190	348	191
rect	347	193	348	194
rect	347	196	348	197
rect	347	205	348	206
rect	347	208	348	209
rect	347	211	348	212
rect	347	220	348	221
rect	347	223	348	224
rect	347	226	348	227
rect	347	229	348	230
rect	347	233	348	234
rect	347	238	348	239
rect	347	241	348	242
rect	347	244	348	245
rect	347	253	348	254
rect	347	256	348	257
rect	347	259	348	260
rect	347	265	348	266
rect	347	268	348	269
rect	347	271	348	272
rect	347	274	348	275
rect	347	280	348	281
rect	347	283	348	284
rect	347	286	348	287
rect	347	295	348	296
rect	347	298	348	299
rect	347	301	348	302
rect	347	313	348	314
rect	347	316	348	317
rect	347	319	348	320
rect	347	322	348	323
rect	347	328	348	329
rect	347	331	348	332
rect	347	337	348	338
rect	347	340	348	341
rect	347	343	348	344
rect	347	349	348	350
rect	347	364	348	365
rect	347	370	348	371
rect	347	373	348	374
rect	347	376	348	377
rect	347	379	348	380
rect	347	385	348	386
rect	348	10	349	11
rect	348	13	349	14
rect	348	16	349	17
rect	348	19	349	20
rect	348	22	349	23
rect	348	25	349	26
rect	348	28	349	29
rect	348	31	349	32
rect	348	34	349	35
rect	348	37	349	38
rect	348	43	349	44
rect	348	46	349	47
rect	348	49	349	50
rect	348	58	349	59
rect	348	61	349	62
rect	348	64	349	65
rect	348	73	349	74
rect	348	76	349	77
rect	348	79	349	80
rect	348	82	349	83
rect	348	91	349	92
rect	348	94	349	95
rect	348	97	349	98
rect	348	100	349	101
rect	348	103	349	104
rect	348	106	349	107
rect	348	118	349	119
rect	348	121	349	122
rect	348	124	349	125
rect	348	127	349	128
rect	348	130	349	131
rect	348	136	349	137
rect	348	139	349	140
rect	348	142	349	143
rect	348	145	349	146
rect	348	148	349	149
rect	348	157	349	158
rect	348	160	349	161
rect	348	163	349	164
rect	348	166	349	167
rect	348	169	349	170
rect	348	175	349	176
rect	348	178	349	179
rect	348	181	349	182
rect	348	184	349	185
rect	348	190	349	191
rect	348	193	349	194
rect	348	196	349	197
rect	348	205	349	206
rect	348	208	349	209
rect	348	211	349	212
rect	348	220	349	221
rect	348	223	349	224
rect	348	226	349	227
rect	348	229	349	230
rect	348	238	349	239
rect	348	241	349	242
rect	348	244	349	245
rect	348	253	349	254
rect	348	256	349	257
rect	348	259	349	260
rect	348	265	349	266
rect	348	268	349	269
rect	348	271	349	272
rect	348	274	349	275
rect	348	280	349	281
rect	348	283	349	284
rect	348	286	349	287
rect	348	295	349	296
rect	348	298	349	299
rect	348	301	349	302
rect	348	313	349	314
rect	348	316	349	317
rect	348	319	349	320
rect	348	322	349	323
rect	348	328	349	329
rect	348	331	349	332
rect	348	337	349	338
rect	348	340	349	341
rect	348	343	349	344
rect	348	349	349	350
rect	348	364	349	365
rect	348	370	349	371
rect	348	373	349	374
rect	348	376	349	377
rect	348	379	349	380
rect	348	385	349	386
rect	349	10	350	11
rect	349	13	350	14
rect	349	16	350	17
rect	349	19	350	20
rect	349	22	350	23
rect	349	25	350	26
rect	349	28	350	29
rect	349	31	350	32
rect	349	34	350	35
rect	349	37	350	38
rect	349	43	350	44
rect	349	46	350	47
rect	349	49	350	50
rect	349	58	350	59
rect	349	61	350	62
rect	349	64	350	65
rect	349	73	350	74
rect	349	76	350	77
rect	349	79	350	80
rect	349	82	350	83
rect	349	86	350	87
rect	349	91	350	92
rect	349	94	350	95
rect	349	97	350	98
rect	349	100	350	101
rect	349	103	350	104
rect	349	106	350	107
rect	349	112	350	113
rect	349	118	350	119
rect	349	121	350	122
rect	349	124	350	125
rect	349	127	350	128
rect	349	130	350	131
rect	349	136	350	137
rect	349	139	350	140
rect	349	142	350	143
rect	349	145	350	146
rect	349	148	350	149
rect	349	157	350	158
rect	349	160	350	161
rect	349	163	350	164
rect	349	166	350	167
rect	349	169	350	170
rect	349	175	350	176
rect	349	178	350	179
rect	349	181	350	182
rect	349	184	350	185
rect	349	190	350	191
rect	349	193	350	194
rect	349	196	350	197
rect	349	205	350	206
rect	349	208	350	209
rect	349	211	350	212
rect	349	220	350	221
rect	349	223	350	224
rect	349	226	350	227
rect	349	229	350	230
rect	349	238	350	239
rect	349	241	350	242
rect	349	244	350	245
rect	349	253	350	254
rect	349	256	350	257
rect	349	259	350	260
rect	349	265	350	266
rect	349	268	350	269
rect	349	271	350	272
rect	349	274	350	275
rect	349	280	350	281
rect	349	283	350	284
rect	349	286	350	287
rect	349	295	350	296
rect	349	298	350	299
rect	349	301	350	302
rect	349	310	350	311
rect	349	313	350	314
rect	349	316	350	317
rect	349	319	350	320
rect	349	322	350	323
rect	349	328	350	329
rect	349	331	350	332
rect	349	337	350	338
rect	349	340	350	341
rect	349	343	350	344
rect	349	349	350	350
rect	349	364	350	365
rect	349	370	350	371
rect	349	373	350	374
rect	349	376	350	377
rect	349	379	350	380
rect	349	385	350	386
rect	350	13	351	14
rect	350	19	351	20
rect	350	22	351	23
rect	350	25	351	26
rect	350	28	351	29
rect	350	31	351	32
rect	350	34	351	35
rect	350	37	351	38
rect	350	43	351	44
rect	350	46	351	47
rect	350	49	351	50
rect	350	58	351	59
rect	350	61	351	62
rect	350	64	351	65
rect	350	73	351	74
rect	350	76	351	77
rect	350	79	351	80
rect	350	82	351	83
rect	350	86	351	87
rect	350	91	351	92
rect	350	94	351	95
rect	350	97	351	98
rect	350	100	351	101
rect	350	103	351	104
rect	350	106	351	107
rect	350	112	351	113
rect	350	118	351	119
rect	350	121	351	122
rect	350	124	351	125
rect	350	130	351	131
rect	350	136	351	137
rect	350	139	351	140
rect	350	142	351	143
rect	350	145	351	146
rect	350	148	351	149
rect	350	157	351	158
rect	350	160	351	161
rect	350	163	351	164
rect	350	166	351	167
rect	350	169	351	170
rect	350	175	351	176
rect	350	178	351	179
rect	350	181	351	182
rect	350	184	351	185
rect	350	190	351	191
rect	350	193	351	194
rect	350	196	351	197
rect	350	205	351	206
rect	350	208	351	209
rect	350	211	351	212
rect	350	220	351	221
rect	350	223	351	224
rect	350	226	351	227
rect	350	229	351	230
rect	350	238	351	239
rect	350	241	351	242
rect	350	253	351	254
rect	350	256	351	257
rect	350	259	351	260
rect	350	265	351	266
rect	350	268	351	269
rect	350	271	351	272
rect	350	274	351	275
rect	350	280	351	281
rect	350	283	351	284
rect	350	286	351	287
rect	350	295	351	296
rect	350	298	351	299
rect	350	301	351	302
rect	350	310	351	311
rect	350	313	351	314
rect	350	316	351	317
rect	350	319	351	320
rect	350	322	351	323
rect	350	328	351	329
rect	350	331	351	332
rect	350	337	351	338
rect	350	340	351	341
rect	350	343	351	344
rect	350	349	351	350
rect	350	364	351	365
rect	350	370	351	371
rect	350	373	351	374
rect	350	376	351	377
rect	350	379	351	380
rect	350	385	351	386
rect	351	13	352	14
rect	351	19	352	20
rect	351	22	352	23
rect	351	25	352	26
rect	351	28	352	29
rect	351	31	352	32
rect	351	34	352	35
rect	351	37	352	38
rect	351	43	352	44
rect	351	46	352	47
rect	351	49	352	50
rect	351	58	352	59
rect	351	61	352	62
rect	351	64	352	65
rect	351	73	352	74
rect	351	76	352	77
rect	351	79	352	80
rect	351	82	352	83
rect	351	86	352	87
rect	351	91	352	92
rect	351	94	352	95
rect	351	97	352	98
rect	351	100	352	101
rect	351	103	352	104
rect	351	106	352	107
rect	351	109	352	110
rect	351	112	352	113
rect	351	118	352	119
rect	351	121	352	122
rect	351	124	352	125
rect	351	130	352	131
rect	351	136	352	137
rect	351	139	352	140
rect	351	142	352	143
rect	351	145	352	146
rect	351	148	352	149
rect	351	157	352	158
rect	351	160	352	161
rect	351	163	352	164
rect	351	166	352	167
rect	351	169	352	170
rect	351	175	352	176
rect	351	178	352	179
rect	351	181	352	182
rect	351	184	352	185
rect	351	190	352	191
rect	351	193	352	194
rect	351	196	352	197
rect	351	205	352	206
rect	351	208	352	209
rect	351	211	352	212
rect	351	220	352	221
rect	351	223	352	224
rect	351	226	352	227
rect	351	229	352	230
rect	351	238	352	239
rect	351	241	352	242
rect	351	247	352	248
rect	351	253	352	254
rect	351	256	352	257
rect	351	259	352	260
rect	351	265	352	266
rect	351	268	352	269
rect	351	271	352	272
rect	351	274	352	275
rect	351	280	352	281
rect	351	283	352	284
rect	351	286	352	287
rect	351	295	352	296
rect	351	298	352	299
rect	351	301	352	302
rect	351	310	352	311
rect	351	313	352	314
rect	351	316	352	317
rect	351	319	352	320
rect	351	322	352	323
rect	351	328	352	329
rect	351	331	352	332
rect	351	337	352	338
rect	351	340	352	341
rect	351	343	352	344
rect	351	349	352	350
rect	351	364	352	365
rect	351	370	352	371
rect	351	373	352	374
rect	351	376	352	377
rect	351	379	352	380
rect	351	385	352	386
rect	352	13	353	14
rect	352	19	353	20
rect	352	25	353	26
rect	352	28	353	29
rect	352	31	353	32
rect	352	34	353	35
rect	352	37	353	38
rect	352	43	353	44
rect	352	46	353	47
rect	352	49	353	50
rect	352	58	353	59
rect	352	61	353	62
rect	352	64	353	65
rect	352	73	353	74
rect	352	76	353	77
rect	352	79	353	80
rect	352	82	353	83
rect	352	91	353	92
rect	352	94	353	95
rect	352	97	353	98
rect	352	100	353	101
rect	352	103	353	104
rect	352	106	353	107
rect	352	109	353	110
rect	352	112	353	113
rect	352	118	353	119
rect	352	121	353	122
rect	352	124	353	125
rect	352	130	353	131
rect	352	136	353	137
rect	352	139	353	140
rect	352	142	353	143
rect	352	148	353	149
rect	352	157	353	158
rect	352	160	353	161
rect	352	163	353	164
rect	352	166	353	167
rect	352	169	353	170
rect	352	175	353	176
rect	352	178	353	179
rect	352	181	353	182
rect	352	184	353	185
rect	352	190	353	191
rect	352	193	353	194
rect	352	196	353	197
rect	352	205	353	206
rect	352	208	353	209
rect	352	211	353	212
rect	352	220	353	221
rect	352	223	353	224
rect	352	226	353	227
rect	352	229	353	230
rect	352	241	353	242
rect	352	247	353	248
rect	352	253	353	254
rect	352	256	353	257
rect	352	259	353	260
rect	352	265	353	266
rect	352	268	353	269
rect	352	271	353	272
rect	352	274	353	275
rect	352	280	353	281
rect	352	283	353	284
rect	352	286	353	287
rect	352	295	353	296
rect	352	298	353	299
rect	352	301	353	302
rect	352	310	353	311
rect	352	313	353	314
rect	352	316	353	317
rect	352	319	353	320
rect	352	322	353	323
rect	352	328	353	329
rect	352	331	353	332
rect	352	337	353	338
rect	352	340	353	341
rect	352	343	353	344
rect	352	349	353	350
rect	352	364	353	365
rect	352	370	353	371
rect	352	373	353	374
rect	352	376	353	377
rect	352	379	353	380
rect	352	385	353	386
rect	353	13	354	14
rect	353	16	354	17
rect	353	19	354	20
rect	353	25	354	26
rect	353	28	354	29
rect	353	31	354	32
rect	353	34	354	35
rect	353	37	354	38
rect	353	43	354	44
rect	353	46	354	47
rect	353	49	354	50
rect	353	58	354	59
rect	353	61	354	62
rect	353	64	354	65
rect	353	73	354	74
rect	353	76	354	77
rect	353	79	354	80
rect	353	82	354	83
rect	353	91	354	92
rect	353	94	354	95
rect	353	97	354	98
rect	353	100	354	101
rect	353	103	354	104
rect	353	106	354	107
rect	353	109	354	110
rect	353	112	354	113
rect	353	118	354	119
rect	353	121	354	122
rect	353	124	354	125
rect	353	127	354	128
rect	353	130	354	131
rect	353	133	354	134
rect	353	136	354	137
rect	353	139	354	140
rect	353	142	354	143
rect	353	148	354	149
rect	353	157	354	158
rect	353	160	354	161
rect	353	163	354	164
rect	353	166	354	167
rect	353	169	354	170
rect	353	175	354	176
rect	353	178	354	179
rect	353	181	354	182
rect	353	184	354	185
rect	353	190	354	191
rect	353	193	354	194
rect	353	196	354	197
rect	353	205	354	206
rect	353	208	354	209
rect	353	211	354	212
rect	353	220	354	221
rect	353	223	354	224
rect	353	226	354	227
rect	353	229	354	230
rect	353	241	354	242
rect	353	244	354	245
rect	353	247	354	248
rect	353	253	354	254
rect	353	256	354	257
rect	353	259	354	260
rect	353	265	354	266
rect	353	268	354	269
rect	353	271	354	272
rect	353	274	354	275
rect	353	280	354	281
rect	353	283	354	284
rect	353	286	354	287
rect	353	295	354	296
rect	353	298	354	299
rect	353	301	354	302
rect	353	310	354	311
rect	353	313	354	314
rect	353	316	354	317
rect	353	319	354	320
rect	353	322	354	323
rect	353	328	354	329
rect	353	331	354	332
rect	353	337	354	338
rect	353	340	354	341
rect	353	343	354	344
rect	353	349	354	350
rect	353	364	354	365
rect	353	370	354	371
rect	353	373	354	374
rect	353	376	354	377
rect	353	379	354	380
rect	353	385	354	386
rect	354	13	355	14
rect	354	16	355	17
rect	354	25	355	26
rect	354	28	355	29
rect	354	31	355	32
rect	354	34	355	35
rect	354	37	355	38
rect	354	43	355	44
rect	354	46	355	47
rect	354	49	355	50
rect	354	58	355	59
rect	354	61	355	62
rect	354	64	355	65
rect	354	73	355	74
rect	354	76	355	77
rect	354	79	355	80
rect	354	82	355	83
rect	354	91	355	92
rect	354	94	355	95
rect	354	97	355	98
rect	354	100	355	101
rect	354	103	355	104
rect	354	106	355	107
rect	354	109	355	110
rect	354	112	355	113
rect	354	121	355	122
rect	354	124	355	125
rect	354	127	355	128
rect	354	130	355	131
rect	354	133	355	134
rect	354	136	355	137
rect	354	139	355	140
rect	354	142	355	143
rect	354	148	355	149
rect	354	157	355	158
rect	354	160	355	161
rect	354	163	355	164
rect	354	166	355	167
rect	354	169	355	170
rect	354	175	355	176
rect	354	178	355	179
rect	354	181	355	182
rect	354	184	355	185
rect	354	190	355	191
rect	354	193	355	194
rect	354	196	355	197
rect	354	205	355	206
rect	354	208	355	209
rect	354	211	355	212
rect	354	220	355	221
rect	354	223	355	224
rect	354	226	355	227
rect	354	229	355	230
rect	354	244	355	245
rect	354	247	355	248
rect	354	253	355	254
rect	354	256	355	257
rect	354	259	355	260
rect	354	265	355	266
rect	354	268	355	269
rect	354	271	355	272
rect	354	274	355	275
rect	354	280	355	281
rect	354	283	355	284
rect	354	286	355	287
rect	354	295	355	296
rect	354	298	355	299
rect	354	301	355	302
rect	354	310	355	311
rect	354	313	355	314
rect	354	316	355	317
rect	354	319	355	320
rect	354	322	355	323
rect	354	328	355	329
rect	354	331	355	332
rect	354	337	355	338
rect	354	340	355	341
rect	354	343	355	344
rect	354	349	355	350
rect	354	364	355	365
rect	354	370	355	371
rect	354	373	355	374
rect	354	376	355	377
rect	354	379	355	380
rect	354	385	355	386
rect	355	13	356	14
rect	355	16	356	17
rect	355	22	356	23
rect	355	25	356	26
rect	355	28	356	29
rect	355	31	356	32
rect	355	34	356	35
rect	355	37	356	38
rect	355	43	356	44
rect	355	46	356	47
rect	355	49	356	50
rect	355	58	356	59
rect	355	61	356	62
rect	355	64	356	65
rect	355	73	356	74
rect	355	76	356	77
rect	355	79	356	80
rect	355	82	356	83
rect	355	91	356	92
rect	355	94	356	95
rect	355	97	356	98
rect	355	100	356	101
rect	355	103	356	104
rect	355	106	356	107
rect	355	109	356	110
rect	355	112	356	113
rect	355	121	356	122
rect	355	124	356	125
rect	355	127	356	128
rect	355	130	356	131
rect	355	133	356	134
rect	355	136	356	137
rect	355	139	356	140
rect	355	142	356	143
rect	355	148	356	149
rect	355	151	356	152
rect	355	157	356	158
rect	355	160	356	161
rect	355	163	356	164
rect	355	166	356	167
rect	355	169	356	170
rect	355	175	356	176
rect	355	178	356	179
rect	355	181	356	182
rect	355	184	356	185
rect	355	190	356	191
rect	355	193	356	194
rect	355	196	356	197
rect	355	205	356	206
rect	355	208	356	209
rect	355	211	356	212
rect	355	220	356	221
rect	355	223	356	224
rect	355	226	356	227
rect	355	229	356	230
rect	355	238	356	239
rect	355	244	356	245
rect	355	247	356	248
rect	355	253	356	254
rect	355	256	356	257
rect	355	259	356	260
rect	355	265	356	266
rect	355	268	356	269
rect	355	271	356	272
rect	355	274	356	275
rect	355	280	356	281
rect	355	283	356	284
rect	355	286	356	287
rect	355	295	356	296
rect	355	298	356	299
rect	355	301	356	302
rect	355	310	356	311
rect	355	313	356	314
rect	355	316	356	317
rect	355	319	356	320
rect	355	322	356	323
rect	355	328	356	329
rect	355	331	356	332
rect	355	337	356	338
rect	355	340	356	341
rect	355	343	356	344
rect	355	349	356	350
rect	355	364	356	365
rect	355	370	356	371
rect	355	373	356	374
rect	355	376	356	377
rect	355	379	356	380
rect	355	385	356	386
rect	356	13	357	14
rect	356	16	357	17
rect	356	22	357	23
rect	356	25	357	26
rect	356	28	357	29
rect	356	31	357	32
rect	356	34	357	35
rect	356	37	357	38
rect	356	46	357	47
rect	356	49	357	50
rect	356	58	357	59
rect	356	61	357	62
rect	356	64	357	65
rect	356	73	357	74
rect	356	76	357	77
rect	356	79	357	80
rect	356	91	357	92
rect	356	94	357	95
rect	356	97	357	98
rect	356	100	357	101
rect	356	103	357	104
rect	356	106	357	107
rect	356	109	357	110
rect	356	112	357	113
rect	356	121	357	122
rect	356	124	357	125
rect	356	127	357	128
rect	356	130	357	131
rect	356	133	357	134
rect	356	136	357	137
rect	356	139	357	140
rect	356	142	357	143
rect	356	148	357	149
rect	356	151	357	152
rect	356	157	357	158
rect	356	160	357	161
rect	356	163	357	164
rect	356	166	357	167
rect	356	169	357	170
rect	356	175	357	176
rect	356	178	357	179
rect	356	181	357	182
rect	356	184	357	185
rect	356	190	357	191
rect	356	193	357	194
rect	356	196	357	197
rect	356	205	357	206
rect	356	208	357	209
rect	356	211	357	212
rect	356	220	357	221
rect	356	223	357	224
rect	356	226	357	227
rect	356	229	357	230
rect	356	238	357	239
rect	356	244	357	245
rect	356	247	357	248
rect	356	253	357	254
rect	356	256	357	257
rect	356	259	357	260
rect	356	265	357	266
rect	356	268	357	269
rect	356	271	357	272
rect	356	274	357	275
rect	356	283	357	284
rect	356	286	357	287
rect	356	295	357	296
rect	356	298	357	299
rect	356	301	357	302
rect	356	310	357	311
rect	356	313	357	314
rect	356	316	357	317
rect	356	319	357	320
rect	356	322	357	323
rect	356	328	357	329
rect	356	331	357	332
rect	356	337	357	338
rect	356	340	357	341
rect	356	343	357	344
rect	356	349	357	350
rect	356	364	357	365
rect	356	370	357	371
rect	356	373	357	374
rect	356	376	357	377
rect	356	379	357	380
rect	356	385	357	386
rect	357	13	358	14
rect	357	16	358	17
rect	357	19	358	20
rect	357	22	358	23
rect	357	25	358	26
rect	357	28	358	29
rect	357	31	358	32
rect	357	34	358	35
rect	357	37	358	38
rect	357	46	358	47
rect	357	49	358	50
rect	357	58	358	59
rect	357	61	358	62
rect	357	64	358	65
rect	357	73	358	74
rect	357	76	358	77
rect	357	79	358	80
rect	357	91	358	92
rect	357	94	358	95
rect	357	97	358	98
rect	357	100	358	101
rect	357	103	358	104
rect	357	106	358	107
rect	357	109	358	110
rect	357	112	358	113
rect	357	121	358	122
rect	357	124	358	125
rect	357	127	358	128
rect	357	130	358	131
rect	357	133	358	134
rect	357	136	358	137
rect	357	139	358	140
rect	357	142	358	143
rect	357	148	358	149
rect	357	151	358	152
rect	357	157	358	158
rect	357	160	358	161
rect	357	163	358	164
rect	357	166	358	167
rect	357	169	358	170
rect	357	175	358	176
rect	357	178	358	179
rect	357	181	358	182
rect	357	184	358	185
rect	357	190	358	191
rect	357	193	358	194
rect	357	196	358	197
rect	357	205	358	206
rect	357	208	358	209
rect	357	211	358	212
rect	357	220	358	221
rect	357	223	358	224
rect	357	226	358	227
rect	357	229	358	230
rect	357	238	358	239
rect	357	244	358	245
rect	357	247	358	248
rect	357	253	358	254
rect	357	256	358	257
rect	357	259	358	260
rect	357	265	358	266
rect	357	268	358	269
rect	357	271	358	272
rect	357	274	358	275
rect	357	283	358	284
rect	357	286	358	287
rect	357	295	358	296
rect	357	298	358	299
rect	357	301	358	302
rect	357	310	358	311
rect	357	313	358	314
rect	357	316	358	317
rect	357	319	358	320
rect	357	322	358	323
rect	357	328	358	329
rect	357	331	358	332
rect	357	337	358	338
rect	357	340	358	341
rect	357	343	358	344
rect	357	349	358	350
rect	357	364	358	365
rect	357	370	358	371
rect	357	373	358	374
rect	357	376	358	377
rect	357	379	358	380
rect	357	385	358	386
rect	358	13	359	14
rect	358	16	359	17
rect	358	19	359	20
rect	358	22	359	23
rect	358	25	359	26
rect	358	31	359	32
rect	358	34	359	35
rect	358	37	359	38
rect	358	46	359	47
rect	358	49	359	50
rect	358	58	359	59
rect	358	61	359	62
rect	358	64	359	65
rect	358	73	359	74
rect	358	76	359	77
rect	358	79	359	80
rect	358	91	359	92
rect	358	94	359	95
rect	358	97	359	98
rect	358	100	359	101
rect	358	103	359	104
rect	358	106	359	107
rect	358	109	359	110
rect	358	112	359	113
rect	358	121	359	122
rect	358	124	359	125
rect	358	127	359	128
rect	358	130	359	131
rect	358	133	359	134
rect	358	139	359	140
rect	358	142	359	143
rect	358	148	359	149
rect	358	151	359	152
rect	358	160	359	161
rect	358	163	359	164
rect	358	166	359	167
rect	358	169	359	170
rect	358	175	359	176
rect	358	178	359	179
rect	358	181	359	182
rect	358	184	359	185
rect	358	190	359	191
rect	358	193	359	194
rect	358	196	359	197
rect	358	205	359	206
rect	358	208	359	209
rect	358	211	359	212
rect	358	220	359	221
rect	358	223	359	224
rect	358	226	359	227
rect	358	229	359	230
rect	358	238	359	239
rect	358	244	359	245
rect	358	247	359	248
rect	358	253	359	254
rect	358	256	359	257
rect	358	259	359	260
rect	358	268	359	269
rect	358	271	359	272
rect	358	274	359	275
rect	358	283	359	284
rect	358	286	359	287
rect	358	295	359	296
rect	358	301	359	302
rect	358	310	359	311
rect	358	313	359	314
rect	358	316	359	317
rect	358	322	359	323
rect	358	328	359	329
rect	358	331	359	332
rect	358	337	359	338
rect	358	340	359	341
rect	358	343	359	344
rect	358	364	359	365
rect	358	370	359	371
rect	358	373	359	374
rect	358	376	359	377
rect	358	379	359	380
rect	358	385	359	386
rect	359	13	360	14
rect	359	16	360	17
rect	359	19	360	20
rect	359	22	360	23
rect	359	25	360	26
rect	359	31	360	32
rect	359	34	360	35
rect	359	37	360	38
rect	359	43	360	44
rect	359	46	360	47
rect	359	49	360	50
rect	359	58	360	59
rect	359	61	360	62
rect	359	64	360	65
rect	359	73	360	74
rect	359	76	360	77
rect	359	79	360	80
rect	359	91	360	92
rect	359	94	360	95
rect	359	97	360	98
rect	359	100	360	101
rect	359	103	360	104
rect	359	106	360	107
rect	359	109	360	110
rect	359	112	360	113
rect	359	115	360	116
rect	359	121	360	122
rect	359	124	360	125
rect	359	127	360	128
rect	359	130	360	131
rect	359	133	360	134
rect	359	139	360	140
rect	359	142	360	143
rect	359	145	360	146
rect	359	148	360	149
rect	359	151	360	152
rect	359	160	360	161
rect	359	163	360	164
rect	359	166	360	167
rect	359	169	360	170
rect	359	175	360	176
rect	359	178	360	179
rect	359	181	360	182
rect	359	184	360	185
rect	359	190	360	191
rect	359	193	360	194
rect	359	196	360	197
rect	359	205	360	206
rect	359	208	360	209
rect	359	211	360	212
rect	359	220	360	221
rect	359	223	360	224
rect	359	226	360	227
rect	359	229	360	230
rect	359	238	360	239
rect	359	241	360	242
rect	359	244	360	245
rect	359	247	360	248
rect	359	253	360	254
rect	359	256	360	257
rect	359	259	360	260
rect	359	268	360	269
rect	359	271	360	272
rect	359	274	360	275
rect	359	280	360	281
rect	359	283	360	284
rect	359	286	360	287
rect	359	295	360	296
rect	359	301	360	302
rect	359	310	360	311
rect	359	313	360	314
rect	359	316	360	317
rect	359	322	360	323
rect	359	328	360	329
rect	359	331	360	332
rect	359	337	360	338
rect	359	340	360	341
rect	359	343	360	344
rect	359	364	360	365
rect	359	370	360	371
rect	359	373	360	374
rect	359	376	360	377
rect	359	379	360	380
rect	359	385	360	386
rect	360	13	361	14
rect	360	16	361	17
rect	360	19	361	20
rect	360	22	361	23
rect	360	25	361	26
rect	360	31	361	32
rect	360	34	361	35
rect	360	43	361	44
rect	360	46	361	47
rect	360	49	361	50
rect	360	58	361	59
rect	360	61	361	62
rect	360	64	361	65
rect	360	73	361	74
rect	360	76	361	77
rect	360	79	361	80
rect	360	91	361	92
rect	360	94	361	95
rect	360	100	361	101
rect	360	103	361	104
rect	360	106	361	107
rect	360	109	361	110
rect	360	112	361	113
rect	360	115	361	116
rect	360	121	361	122
rect	360	124	361	125
rect	360	127	361	128
rect	360	133	361	134
rect	360	139	361	140
rect	360	142	361	143
rect	360	145	361	146
rect	360	151	361	152
rect	360	163	361	164
rect	360	166	361	167
rect	360	169	361	170
rect	360	175	361	176
rect	360	178	361	179
rect	360	181	361	182
rect	360	184	361	185
rect	360	190	361	191
rect	360	193	361	194
rect	360	196	361	197
rect	360	205	361	206
rect	360	208	361	209
rect	360	211	361	212
rect	360	220	361	221
rect	360	223	361	224
rect	360	226	361	227
rect	360	229	361	230
rect	360	238	361	239
rect	360	241	361	242
rect	360	244	361	245
rect	360	247	361	248
rect	360	253	361	254
rect	360	256	361	257
rect	360	259	361	260
rect	360	271	361	272
rect	360	274	361	275
rect	360	280	361	281
rect	360	283	361	284
rect	360	286	361	287
rect	360	295	361	296
rect	360	301	361	302
rect	360	310	361	311
rect	360	313	361	314
rect	360	316	361	317
rect	360	328	361	329
rect	360	331	361	332
rect	360	337	361	338
rect	360	340	361	341
rect	360	343	361	344
rect	360	370	361	371
rect	360	373	361	374
rect	360	376	361	377
rect	360	379	361	380
rect	361	13	362	14
rect	361	16	362	17
rect	361	19	362	20
rect	361	22	362	23
rect	361	25	362	26
rect	361	28	362	29
rect	361	31	362	32
rect	361	34	362	35
rect	361	43	362	44
rect	361	46	362	47
rect	361	49	362	50
rect	361	58	362	59
rect	361	61	362	62
rect	361	64	362	65
rect	361	73	362	74
rect	361	76	362	77
rect	361	79	362	80
rect	361	88	362	89
rect	361	91	362	92
rect	361	94	362	95
rect	361	100	362	101
rect	361	103	362	104
rect	361	106	362	107
rect	361	109	362	110
rect	361	112	362	113
rect	361	115	362	116
rect	361	118	362	119
rect	361	121	362	122
rect	361	124	362	125
rect	361	127	362	128
rect	361	133	362	134
rect	361	136	362	137
rect	361	139	362	140
rect	361	142	362	143
rect	361	145	362	146
rect	361	151	362	152
rect	361	157	362	158
rect	361	163	362	164
rect	361	166	362	167
rect	361	169	362	170
rect	361	175	362	176
rect	361	178	362	179
rect	361	181	362	182
rect	361	184	362	185
rect	361	190	362	191
rect	361	193	362	194
rect	361	196	362	197
rect	361	205	362	206
rect	361	208	362	209
rect	361	211	362	212
rect	361	220	362	221
rect	361	223	362	224
rect	361	226	362	227
rect	361	229	362	230
rect	361	238	362	239
rect	361	241	362	242
rect	361	244	362	245
rect	361	247	362	248
rect	361	253	362	254
rect	361	256	362	257
rect	361	259	362	260
rect	361	265	362	266
rect	361	271	362	272
rect	361	274	362	275
rect	361	280	362	281
rect	361	283	362	284
rect	361	286	362	287
rect	361	295	362	296
rect	361	298	362	299
rect	361	301	362	302
rect	361	310	362	311
rect	361	313	362	314
rect	361	316	362	317
rect	361	328	362	329
rect	361	331	362	332
rect	361	337	362	338
rect	361	340	362	341
rect	361	343	362	344
rect	361	355	362	356
rect	361	367	362	368
rect	361	370	362	371
rect	361	373	362	374
rect	361	376	362	377
rect	361	379	362	380
rect	362	13	363	14
rect	362	16	363	17
rect	362	19	363	20
rect	362	22	363	23
rect	362	25	363	26
rect	362	28	363	29
rect	362	31	363	32
rect	362	34	363	35
rect	362	43	363	44
rect	362	46	363	47
rect	362	49	363	50
rect	362	58	363	59
rect	362	61	363	62
rect	362	64	363	65
rect	362	76	363	77
rect	362	79	363	80
rect	362	88	363	89
rect	362	91	363	92
rect	362	94	363	95
rect	362	100	363	101
rect	362	103	363	104
rect	362	109	363	110
rect	362	112	363	113
rect	362	115	363	116
rect	362	118	363	119
rect	362	121	363	122
rect	362	124	363	125
rect	362	127	363	128
rect	362	133	363	134
rect	362	136	363	137
rect	362	139	363	140
rect	362	145	363	146
rect	362	151	363	152
rect	362	157	363	158
rect	362	166	363	167
rect	362	169	363	170
rect	362	178	363	179
rect	362	181	363	182
rect	362	184	363	185
rect	362	193	363	194
rect	362	196	363	197
rect	362	205	363	206
rect	362	208	363	209
rect	362	211	363	212
rect	362	220	363	221
rect	362	223	363	224
rect	362	226	363	227
rect	362	229	363	230
rect	362	238	363	239
rect	362	241	363	242
rect	362	244	363	245
rect	362	247	363	248
rect	362	253	363	254
rect	362	256	363	257
rect	362	259	363	260
rect	362	265	363	266
rect	362	271	363	272
rect	362	280	363	281
rect	362	283	363	284
rect	362	286	363	287
rect	362	295	363	296
rect	362	298	363	299
rect	362	301	363	302
rect	362	310	363	311
rect	362	328	363	329
rect	362	331	363	332
rect	362	337	363	338
rect	362	340	363	341
rect	362	343	363	344
rect	362	355	363	356
rect	362	367	363	368
rect	362	370	363	371
rect	362	373	363	374
rect	362	376	363	377
rect	363	4	364	5
rect	363	13	364	14
rect	363	16	364	17
rect	363	19	364	20
rect	363	22	364	23
rect	363	25	364	26
rect	363	28	364	29
rect	363	31	364	32
rect	363	34	364	35
rect	363	43	364	44
rect	363	46	364	47
rect	363	49	364	50
rect	363	58	364	59
rect	363	61	364	62
rect	363	64	364	65
rect	363	76	364	77
rect	363	79	364	80
rect	363	88	364	89
rect	363	91	364	92
rect	363	94	364	95
rect	363	97	364	98
rect	363	100	364	101
rect	363	103	364	104
rect	363	109	364	110
rect	363	112	364	113
rect	363	115	364	116
rect	363	118	364	119
rect	363	121	364	122
rect	363	124	364	125
rect	363	127	364	128
rect	363	130	364	131
rect	363	133	364	134
rect	363	136	364	137
rect	363	139	364	140
rect	363	145	364	146
rect	363	151	364	152
rect	363	154	364	155
rect	363	157	364	158
rect	363	166	364	167
rect	363	169	364	170
rect	363	178	364	179
rect	363	181	364	182
rect	363	184	364	185
rect	363	193	364	194
rect	363	196	364	197
rect	363	205	364	206
rect	363	208	364	209
rect	363	211	364	212
rect	363	220	364	221
rect	363	223	364	224
rect	363	226	364	227
rect	363	229	364	230
rect	363	238	364	239
rect	363	241	364	242
rect	363	244	364	245
rect	363	247	364	248
rect	363	253	364	254
rect	363	256	364	257
rect	363	259	364	260
rect	363	265	364	266
rect	363	268	364	269
rect	363	271	364	272
rect	363	280	364	281
rect	363	283	364	284
rect	363	286	364	287
rect	363	292	364	293
rect	363	295	364	296
rect	363	298	364	299
rect	363	301	364	302
rect	363	310	364	311
rect	363	322	364	323
rect	363	328	364	329
rect	363	331	364	332
rect	363	337	364	338
rect	363	340	364	341
rect	363	343	364	344
rect	363	355	364	356
rect	363	364	364	365
rect	363	367	364	368
rect	363	370	364	371
rect	363	373	364	374
rect	363	376	364	377
rect	364	4	365	5
rect	364	13	365	14
rect	364	16	365	17
rect	364	19	365	20
rect	364	22	365	23
rect	364	28	365	29
rect	364	31	365	32
rect	364	34	365	35
rect	364	43	365	44
rect	364	46	365	47
rect	364	49	365	50
rect	364	58	365	59
rect	364	61	365	62
rect	364	76	365	77
rect	364	79	365	80
rect	364	88	365	89
rect	364	94	365	95
rect	364	97	365	98
rect	364	100	365	101
rect	364	103	365	104
rect	364	109	365	110
rect	364	112	365	113
rect	364	115	365	116
rect	364	118	365	119
rect	364	127	365	128
rect	364	130	365	131
rect	364	133	365	134
rect	364	136	365	137
rect	364	139	365	140
rect	364	145	365	146
rect	364	151	365	152
rect	364	154	365	155
rect	364	157	365	158
rect	364	169	365	170
rect	364	181	365	182
rect	364	184	365	185
rect	364	193	365	194
rect	364	205	365	206
rect	364	208	365	209
rect	364	223	365	224
rect	364	226	365	227
rect	364	229	365	230
rect	364	238	365	239
rect	364	241	365	242
rect	364	244	365	245
rect	364	247	365	248
rect	364	253	365	254
rect	364	256	365	257
rect	364	259	365	260
rect	364	265	365	266
rect	364	268	365	269
rect	364	280	365	281
rect	364	283	365	284
rect	364	292	365	293
rect	364	295	365	296
rect	364	298	365	299
rect	364	301	365	302
rect	364	310	365	311
rect	364	322	365	323
rect	364	328	365	329
rect	364	331	365	332
rect	364	337	365	338
rect	364	340	365	341
rect	364	355	365	356
rect	364	364	365	365
rect	364	367	365	368
rect	364	370	365	371
rect	364	376	365	377
rect	365	4	366	5
rect	365	13	366	14
rect	365	16	366	17
rect	365	19	366	20
rect	365	22	366	23
rect	365	28	366	29
rect	365	31	366	32
rect	365	34	366	35
rect	365	40	366	41
rect	365	43	366	44
rect	365	46	366	47
rect	365	49	366	50
rect	365	58	366	59
rect	365	61	366	62
rect	365	67	366	68
rect	365	73	366	74
rect	365	76	366	77
rect	365	79	366	80
rect	365	88	366	89
rect	365	94	366	95
rect	365	97	366	98
rect	365	100	366	101
rect	365	103	366	104
rect	365	106	366	107
rect	365	109	366	110
rect	365	112	366	113
rect	365	115	366	116
rect	365	118	366	119
rect	365	127	366	128
rect	365	130	366	131
rect	365	133	366	134
rect	365	136	366	137
rect	365	139	366	140
rect	365	145	366	146
rect	365	151	366	152
rect	365	154	366	155
rect	365	157	366	158
rect	365	160	366	161
rect	365	163	366	164
rect	365	169	366	170
rect	365	172	366	173
rect	365	181	366	182
rect	365	184	366	185
rect	365	187	366	188
rect	365	193	366	194
rect	365	199	366	200
rect	365	205	366	206
rect	365	208	366	209
rect	365	218	366	219
rect	365	223	366	224
rect	365	226	366	227
rect	365	229	366	230
rect	365	238	366	239
rect	365	241	366	242
rect	365	244	366	245
rect	365	247	366	248
rect	365	250	366	251
rect	365	253	366	254
rect	365	256	366	257
rect	365	259	366	260
rect	365	265	366	266
rect	365	268	366	269
rect	365	277	366	278
rect	365	280	366	281
rect	365	283	366	284
rect	365	292	366	293
rect	365	295	366	296
rect	365	298	366	299
rect	365	301	366	302
rect	365	310	366	311
rect	365	313	366	314
rect	365	319	366	320
rect	365	322	366	323
rect	365	325	366	326
rect	365	328	366	329
rect	365	331	366	332
rect	365	337	366	338
rect	365	340	366	341
rect	365	355	366	356
rect	365	358	366	359
rect	365	364	366	365
rect	365	367	366	368
rect	365	370	366	371
rect	365	376	366	377
rect	366	4	367	5
rect	366	13	367	14
rect	366	16	367	17
rect	366	19	367	20
rect	366	22	367	23
rect	366	28	367	29
rect	366	34	367	35
rect	366	40	367	41
rect	366	43	367	44
rect	366	49	367	50
rect	366	61	367	62
rect	366	67	367	68
rect	366	73	367	74
rect	366	76	367	77
rect	366	79	367	80
rect	366	88	367	89
rect	366	97	367	98
rect	366	100	367	101
rect	366	103	367	104
rect	366	106	367	107
rect	366	109	367	110
rect	366	112	367	113
rect	366	115	367	116
rect	366	118	367	119
rect	366	127	367	128
rect	366	130	367	131
rect	366	133	367	134
rect	366	136	367	137
rect	366	145	367	146
rect	366	151	367	152
rect	366	154	367	155
rect	366	157	367	158
rect	366	160	367	161
rect	366	163	367	164
rect	366	172	367	173
rect	366	187	367	188
rect	366	193	367	194
rect	366	199	367	200
rect	366	205	367	206
rect	366	218	367	219
rect	366	229	367	230
rect	366	238	367	239
rect	366	241	367	242
rect	366	244	367	245
rect	366	247	367	248
rect	366	250	367	251
rect	366	253	367	254
rect	366	256	367	257
rect	366	259	367	260
rect	366	265	367	266
rect	366	268	367	269
rect	366	277	367	278
rect	366	280	367	281
rect	366	283	367	284
rect	366	292	367	293
rect	366	295	367	296
rect	366	298	367	299
rect	366	301	367	302
rect	366	310	367	311
rect	366	313	367	314
rect	366	319	367	320
rect	366	322	367	323
rect	366	325	367	326
rect	366	328	367	329
rect	366	331	367	332
rect	366	337	367	338
rect	366	340	367	341
rect	366	355	367	356
rect	366	358	367	359
rect	366	364	367	365
rect	366	367	367	368
rect	366	370	367	371
rect	367	4	368	5
rect	367	13	368	14
rect	367	16	368	17
rect	367	19	368	20
rect	367	22	368	23
rect	367	25	368	26
rect	367	28	368	29
rect	367	34	368	35
rect	367	37	368	38
rect	367	40	368	41
rect	367	43	368	44
rect	367	49	368	50
rect	367	61	368	62
rect	367	64	368	65
rect	367	67	368	68
rect	367	73	368	74
rect	367	76	368	77
rect	367	79	368	80
rect	367	88	368	89
rect	367	91	368	92
rect	367	97	368	98
rect	367	100	368	101
rect	367	103	368	104
rect	367	106	368	107
rect	367	109	368	110
rect	367	112	368	113
rect	367	115	368	116
rect	367	118	368	119
rect	367	121	368	122
rect	367	127	368	128
rect	367	130	368	131
rect	367	133	368	134
rect	367	136	368	137
rect	367	142	368	143
rect	367	145	368	146
rect	367	151	368	152
rect	367	154	368	155
rect	367	157	368	158
rect	367	160	368	161
rect	367	163	368	164
rect	367	172	368	173
rect	367	178	368	179
rect	367	187	368	188
rect	367	190	368	191
rect	367	193	368	194
rect	367	199	368	200
rect	367	205	368	206
rect	367	211	368	212
rect	367	218	368	219
rect	367	220	368	221
rect	367	229	368	230
rect	367	238	368	239
rect	367	241	368	242
rect	367	244	368	245
rect	367	247	368	248
rect	367	250	368	251
rect	367	253	368	254
rect	367	256	368	257
rect	367	259	368	260
rect	367	265	368	266
rect	367	268	368	269
rect	367	277	368	278
rect	367	280	368	281
rect	367	283	368	284
rect	367	292	368	293
rect	367	295	368	296
rect	367	298	368	299
rect	367	301	368	302
rect	367	310	368	311
rect	367	313	368	314
rect	367	319	368	320
rect	367	322	368	323
rect	367	325	368	326
rect	367	328	368	329
rect	367	331	368	332
rect	367	337	368	338
rect	367	340	368	341
rect	367	349	368	350
rect	367	352	368	353
rect	367	355	368	356
rect	367	358	368	359
rect	367	364	368	365
rect	367	367	368	368
rect	367	370	368	371
rect	368	4	369	5
rect	368	13	369	14
rect	368	16	369	17
rect	368	19	369	20
rect	368	22	369	23
rect	368	25	369	26
rect	368	28	369	29
rect	368	37	369	38
rect	368	40	369	41
rect	368	43	369	44
rect	368	64	369	65
rect	368	67	369	68
rect	368	73	369	74
rect	368	76	369	77
rect	368	79	369	80
rect	368	88	369	89
rect	368	91	369	92
rect	368	97	369	98
rect	368	106	369	107
rect	368	109	369	110
rect	368	112	369	113
rect	368	115	369	116
rect	368	118	369	119
rect	368	121	369	122
rect	368	127	369	128
rect	368	130	369	131
rect	368	133	369	134
rect	368	136	369	137
rect	368	142	369	143
rect	368	145	369	146
rect	368	151	369	152
rect	368	154	369	155
rect	368	157	369	158
rect	368	160	369	161
rect	368	163	369	164
rect	368	172	369	173
rect	368	178	369	179
rect	368	187	369	188
rect	368	190	369	191
rect	368	199	369	200
rect	368	211	369	212
rect	368	220	369	221
rect	368	238	369	239
rect	368	241	369	242
rect	368	244	369	245
rect	368	247	369	248
rect	368	250	369	251
rect	368	253	369	254
rect	368	256	369	257
rect	368	265	369	266
rect	368	268	369	269
rect	368	277	369	278
rect	368	280	369	281
rect	368	292	369	293
rect	368	295	369	296
rect	368	298	369	299
rect	368	301	369	302
rect	368	310	369	311
rect	368	313	369	314
rect	368	319	369	320
rect	368	322	369	323
rect	368	325	369	326
rect	368	349	369	350
rect	368	352	369	353
rect	368	355	369	356
rect	368	358	369	359
rect	368	364	369	365
rect	368	367	369	368
rect	369	4	370	5
rect	369	13	370	14
rect	369	16	370	17
rect	369	19	370	20
rect	369	22	370	23
rect	369	25	370	26
rect	369	28	370	29
rect	369	31	370	32
rect	369	37	370	38
rect	369	40	370	41
rect	369	43	370	44
rect	369	46	370	47
rect	369	55	370	56
rect	369	64	370	65
rect	369	67	370	68
rect	369	73	370	74
rect	369	76	370	77
rect	369	79	370	80
rect	369	88	370	89
rect	369	91	370	92
rect	369	94	370	95
rect	369	97	370	98
rect	369	106	370	107
rect	369	109	370	110
rect	369	112	370	113
rect	369	115	370	116
rect	369	118	370	119
rect	369	121	370	122
rect	369	124	370	125
rect	369	127	370	128
rect	369	130	370	131
rect	369	133	370	134
rect	369	136	370	137
rect	369	142	370	143
rect	369	145	370	146
rect	369	148	370	149
rect	369	151	370	152
rect	369	154	370	155
rect	369	157	370	158
rect	369	160	370	161
rect	369	163	370	164
rect	369	169	370	170
rect	369	172	370	173
rect	369	175	370	176
rect	369	178	370	179
rect	369	187	370	188
rect	369	190	370	191
rect	369	199	370	200
rect	369	208	370	209
rect	369	211	370	212
rect	369	220	370	221
rect	369	223	370	224
rect	369	226	370	227
rect	369	235	370	236
rect	369	238	370	239
rect	369	241	370	242
rect	369	244	370	245
rect	369	247	370	248
rect	369	250	370	251
rect	369	253	370	254
rect	369	256	370	257
rect	369	262	370	263
rect	369	265	370	266
rect	369	268	370	269
rect	369	277	370	278
rect	369	280	370	281
rect	369	289	370	290
rect	369	292	370	293
rect	369	295	370	296
rect	369	298	370	299
rect	369	301	370	302
rect	369	310	370	311
rect	369	313	370	314
rect	369	319	370	320
rect	369	322	370	323
rect	369	325	370	326
rect	369	349	370	350
rect	369	352	370	353
rect	369	355	370	356
rect	369	358	370	359
rect	369	364	370	365
rect	369	367	370	368
rect	376	4	377	5
rect	376	10	377	11
rect	376	13	377	14
rect	376	16	377	17
rect	376	19	377	20
rect	376	22	377	23
rect	376	25	377	26
rect	376	28	377	29
rect	376	37	377	38
rect	376	40	377	41
rect	376	43	377	44
rect	376	46	377	47
rect	376	55	377	56
rect	376	64	377	65
rect	376	67	377	68
rect	376	76	377	77
rect	376	79	377	80
rect	376	85	377	86
rect	376	88	377	89
rect	376	91	377	92
rect	376	94	377	95
rect	376	97	377	98
rect	376	106	377	107
rect	376	109	377	110
rect	376	112	377	113
rect	376	115	377	116
rect	376	118	377	119
rect	376	121	377	122
rect	376	124	377	125
rect	376	127	377	128
rect	376	130	377	131
rect	376	133	377	134
rect	376	136	377	137
rect	376	145	377	146
rect	376	148	377	149
rect	376	151	377	152
rect	376	154	377	155
rect	376	157	377	158
rect	376	160	377	161
rect	376	163	377	164
rect	376	172	377	173
rect	376	175	377	176
rect	376	178	377	179
rect	376	187	377	188
rect	376	190	377	191
rect	376	199	377	200
rect	376	208	377	209
rect	376	211	377	212
rect	376	220	377	221
rect	376	223	377	224
rect	376	226	377	227
rect	376	229	377	230
rect	376	235	377	236
rect	376	238	377	239
rect	376	241	377	242
rect	376	244	377	245
rect	376	247	377	248
rect	376	250	377	251
rect	376	253	377	254
rect	376	256	377	257
rect	376	265	377	266
rect	376	268	377	269
rect	376	271	377	272
rect	376	277	377	278
rect	376	280	377	281
rect	376	289	377	290
rect	376	292	377	293
rect	376	295	377	296
rect	376	298	377	299
rect	376	301	377	302
rect	376	310	377	311
rect	376	319	377	320
rect	376	322	377	323
rect	376	325	377	326
rect	376	331	377	332
rect	376	352	377	353
rect	376	355	377	356
rect	376	358	377	359
rect	376	364	377	365
rect	376	367	377	368
rect	377	4	378	5
rect	377	10	378	11
rect	377	13	378	14
rect	377	16	378	17
rect	377	19	378	20
rect	377	22	378	23
rect	377	25	378	26
rect	377	28	378	29
rect	377	37	378	38
rect	377	40	378	41
rect	377	43	378	44
rect	377	46	378	47
rect	377	55	378	56
rect	377	64	378	65
rect	377	67	378	68
rect	377	76	378	77
rect	377	79	378	80
rect	377	85	378	86
rect	377	88	378	89
rect	377	91	378	92
rect	377	94	378	95
rect	377	97	378	98
rect	377	106	378	107
rect	377	109	378	110
rect	377	112	378	113
rect	377	115	378	116
rect	377	118	378	119
rect	377	121	378	122
rect	377	124	378	125
rect	377	127	378	128
rect	377	130	378	131
rect	377	133	378	134
rect	377	136	378	137
rect	377	145	378	146
rect	377	148	378	149
rect	377	151	378	152
rect	377	154	378	155
rect	377	157	378	158
rect	377	160	378	161
rect	377	163	378	164
rect	377	175	378	176
rect	377	178	378	179
rect	377	187	378	188
rect	377	190	378	191
rect	377	199	378	200
rect	377	208	378	209
rect	377	211	378	212
rect	377	220	378	221
rect	377	223	378	224
rect	377	226	378	227
rect	377	229	378	230
rect	377	235	378	236
rect	377	238	378	239
rect	377	241	378	242
rect	377	244	378	245
rect	377	247	378	248
rect	377	250	378	251
rect	377	253	378	254
rect	377	256	378	257
rect	377	265	378	266
rect	377	268	378	269
rect	377	271	378	272
rect	377	277	378	278
rect	377	280	378	281
rect	377	289	378	290
rect	377	292	378	293
rect	377	295	378	296
rect	377	298	378	299
rect	377	301	378	302
rect	377	310	378	311
rect	377	319	378	320
rect	377	322	378	323
rect	377	325	378	326
rect	377	331	378	332
rect	377	352	378	353
rect	377	355	378	356
rect	377	358	378	359
rect	377	364	378	365
rect	377	367	378	368
rect	378	4	379	5
rect	378	10	379	11
rect	378	13	379	14
rect	378	16	379	17
rect	378	19	379	20
rect	378	22	379	23
rect	378	25	379	26
rect	378	28	379	29
rect	378	37	379	38
rect	378	40	379	41
rect	378	43	379	44
rect	378	46	379	47
rect	378	55	379	56
rect	378	64	379	65
rect	378	67	379	68
rect	378	76	379	77
rect	378	79	379	80
rect	378	85	379	86
rect	378	88	379	89
rect	378	91	379	92
rect	378	94	379	95
rect	378	97	379	98
rect	378	106	379	107
rect	378	109	379	110
rect	378	112	379	113
rect	378	115	379	116
rect	378	118	379	119
rect	378	121	379	122
rect	378	124	379	125
rect	378	127	379	128
rect	378	130	379	131
rect	378	133	379	134
rect	378	136	379	137
rect	378	145	379	146
rect	378	148	379	149
rect	378	151	379	152
rect	378	154	379	155
rect	378	157	379	158
rect	378	160	379	161
rect	378	163	379	164
rect	378	169	379	170
rect	378	175	379	176
rect	378	178	379	179
rect	378	187	379	188
rect	378	190	379	191
rect	378	199	379	200
rect	378	208	379	209
rect	378	211	379	212
rect	378	220	379	221
rect	378	223	379	224
rect	378	226	379	227
rect	378	229	379	230
rect	378	235	379	236
rect	378	238	379	239
rect	378	241	379	242
rect	378	244	379	245
rect	378	247	379	248
rect	378	250	379	251
rect	378	253	379	254
rect	378	256	379	257
rect	378	265	379	266
rect	378	268	379	269
rect	378	271	379	272
rect	378	277	379	278
rect	378	280	379	281
rect	378	289	379	290
rect	378	292	379	293
rect	378	295	379	296
rect	378	298	379	299
rect	378	301	379	302
rect	378	310	379	311
rect	378	319	379	320
rect	378	322	379	323
rect	378	325	379	326
rect	378	331	379	332
rect	378	352	379	353
rect	378	355	379	356
rect	378	358	379	359
rect	378	364	379	365
rect	378	367	379	368
rect	379	4	380	5
rect	379	10	380	11
rect	379	13	380	14
rect	379	16	380	17
rect	379	19	380	20
rect	379	22	380	23
rect	379	25	380	26
rect	379	28	380	29
rect	379	37	380	38
rect	379	40	380	41
rect	379	43	380	44
rect	379	46	380	47
rect	379	55	380	56
rect	379	64	380	65
rect	379	67	380	68
rect	379	76	380	77
rect	379	79	380	80
rect	379	85	380	86
rect	379	88	380	89
rect	379	91	380	92
rect	379	94	380	95
rect	379	97	380	98
rect	379	106	380	107
rect	379	109	380	110
rect	379	112	380	113
rect	379	115	380	116
rect	379	118	380	119
rect	379	121	380	122
rect	379	124	380	125
rect	379	127	380	128
rect	379	130	380	131
rect	379	133	380	134
rect	379	136	380	137
rect	379	145	380	146
rect	379	148	380	149
rect	379	151	380	152
rect	379	154	380	155
rect	379	157	380	158
rect	379	160	380	161
rect	379	163	380	164
rect	379	169	380	170
rect	379	175	380	176
rect	379	178	380	179
rect	379	190	380	191
rect	379	199	380	200
rect	379	208	380	209
rect	379	211	380	212
rect	379	220	380	221
rect	379	223	380	224
rect	379	226	380	227
rect	379	229	380	230
rect	379	235	380	236
rect	379	238	380	239
rect	379	241	380	242
rect	379	244	380	245
rect	379	247	380	248
rect	379	250	380	251
rect	379	253	380	254
rect	379	256	380	257
rect	379	265	380	266
rect	379	268	380	269
rect	379	271	380	272
rect	379	277	380	278
rect	379	280	380	281
rect	379	289	380	290
rect	379	292	380	293
rect	379	295	380	296
rect	379	298	380	299
rect	379	301	380	302
rect	379	310	380	311
rect	379	319	380	320
rect	379	322	380	323
rect	379	325	380	326
rect	379	331	380	332
rect	379	352	380	353
rect	379	355	380	356
rect	379	358	380	359
rect	379	364	380	365
rect	379	367	380	368
rect	380	4	381	5
rect	380	10	381	11
rect	380	13	381	14
rect	380	16	381	17
rect	380	19	381	20
rect	380	22	381	23
rect	380	25	381	26
rect	380	28	381	29
rect	380	37	381	38
rect	380	40	381	41
rect	380	43	381	44
rect	380	46	381	47
rect	380	55	381	56
rect	380	64	381	65
rect	380	67	381	68
rect	380	76	381	77
rect	380	79	381	80
rect	380	85	381	86
rect	380	88	381	89
rect	380	91	381	92
rect	380	94	381	95
rect	380	97	381	98
rect	380	106	381	107
rect	380	109	381	110
rect	380	112	381	113
rect	380	115	381	116
rect	380	118	381	119
rect	380	121	381	122
rect	380	124	381	125
rect	380	127	381	128
rect	380	130	381	131
rect	380	133	381	134
rect	380	136	381	137
rect	380	145	381	146
rect	380	148	381	149
rect	380	151	381	152
rect	380	154	381	155
rect	380	157	381	158
rect	380	160	381	161
rect	380	163	381	164
rect	380	169	381	170
rect	380	172	381	173
rect	380	175	381	176
rect	380	178	381	179
rect	380	190	381	191
rect	380	199	381	200
rect	380	208	381	209
rect	380	211	381	212
rect	380	220	381	221
rect	380	223	381	224
rect	380	226	381	227
rect	380	229	381	230
rect	380	235	381	236
rect	380	238	381	239
rect	380	241	381	242
rect	380	244	381	245
rect	380	247	381	248
rect	380	250	381	251
rect	380	253	381	254
rect	380	256	381	257
rect	380	265	381	266
rect	380	268	381	269
rect	380	271	381	272
rect	380	277	381	278
rect	380	280	381	281
rect	380	289	381	290
rect	380	292	381	293
rect	380	295	381	296
rect	380	298	381	299
rect	380	301	381	302
rect	380	310	381	311
rect	380	319	381	320
rect	380	322	381	323
rect	380	325	381	326
rect	380	331	381	332
rect	380	352	381	353
rect	380	355	381	356
rect	380	358	381	359
rect	380	364	381	365
rect	380	367	381	368
rect	381	4	382	5
rect	381	10	382	11
rect	381	13	382	14
rect	381	16	382	17
rect	381	19	382	20
rect	381	22	382	23
rect	381	25	382	26
rect	381	28	382	29
rect	381	37	382	38
rect	381	40	382	41
rect	381	43	382	44
rect	381	46	382	47
rect	381	55	382	56
rect	381	64	382	65
rect	381	67	382	68
rect	381	76	382	77
rect	381	79	382	80
rect	381	85	382	86
rect	381	88	382	89
rect	381	91	382	92
rect	381	94	382	95
rect	381	97	382	98
rect	381	106	382	107
rect	381	109	382	110
rect	381	112	382	113
rect	381	115	382	116
rect	381	118	382	119
rect	381	121	382	122
rect	381	124	382	125
rect	381	127	382	128
rect	381	130	382	131
rect	381	133	382	134
rect	381	136	382	137
rect	381	145	382	146
rect	381	151	382	152
rect	381	154	382	155
rect	381	157	382	158
rect	381	160	382	161
rect	381	163	382	164
rect	381	169	382	170
rect	381	172	382	173
rect	381	175	382	176
rect	381	178	382	179
rect	381	190	382	191
rect	381	199	382	200
rect	381	208	382	209
rect	381	211	382	212
rect	381	220	382	221
rect	381	223	382	224
rect	381	226	382	227
rect	381	229	382	230
rect	381	235	382	236
rect	381	238	382	239
rect	381	241	382	242
rect	381	244	382	245
rect	381	247	382	248
rect	381	250	382	251
rect	381	253	382	254
rect	381	256	382	257
rect	381	265	382	266
rect	381	268	382	269
rect	381	271	382	272
rect	381	277	382	278
rect	381	280	382	281
rect	381	289	382	290
rect	381	292	382	293
rect	381	295	382	296
rect	381	298	382	299
rect	381	301	382	302
rect	381	310	382	311
rect	381	319	382	320
rect	381	322	382	323
rect	381	325	382	326
rect	381	331	382	332
rect	381	352	382	353
rect	381	355	382	356
rect	381	358	382	359
rect	381	364	382	365
rect	381	367	382	368
rect	382	4	383	5
rect	382	10	383	11
rect	382	13	383	14
rect	382	16	383	17
rect	382	19	383	20
rect	382	22	383	23
rect	382	25	383	26
rect	382	28	383	29
rect	382	37	383	38
rect	382	40	383	41
rect	382	43	383	44
rect	382	46	383	47
rect	382	55	383	56
rect	382	64	383	65
rect	382	67	383	68
rect	382	76	383	77
rect	382	79	383	80
rect	382	85	383	86
rect	382	88	383	89
rect	382	91	383	92
rect	382	94	383	95
rect	382	97	383	98
rect	382	106	383	107
rect	382	109	383	110
rect	382	112	383	113
rect	382	115	383	116
rect	382	118	383	119
rect	382	121	383	122
rect	382	124	383	125
rect	382	127	383	128
rect	382	130	383	131
rect	382	133	383	134
rect	382	136	383	137
rect	382	145	383	146
rect	382	151	383	152
rect	382	154	383	155
rect	382	157	383	158
rect	382	160	383	161
rect	382	163	383	164
rect	382	169	383	170
rect	382	172	383	173
rect	382	175	383	176
rect	382	178	383	179
rect	382	187	383	188
rect	382	190	383	191
rect	382	199	383	200
rect	382	208	383	209
rect	382	211	383	212
rect	382	220	383	221
rect	382	223	383	224
rect	382	226	383	227
rect	382	229	383	230
rect	382	235	383	236
rect	382	238	383	239
rect	382	241	383	242
rect	382	244	383	245
rect	382	247	383	248
rect	382	250	383	251
rect	382	253	383	254
rect	382	256	383	257
rect	382	265	383	266
rect	382	268	383	269
rect	382	271	383	272
rect	382	277	383	278
rect	382	280	383	281
rect	382	289	383	290
rect	382	292	383	293
rect	382	295	383	296
rect	382	298	383	299
rect	382	301	383	302
rect	382	310	383	311
rect	382	319	383	320
rect	382	322	383	323
rect	382	325	383	326
rect	382	331	383	332
rect	382	352	383	353
rect	382	355	383	356
rect	382	358	383	359
rect	382	364	383	365
rect	382	367	383	368
rect	383	4	384	5
rect	383	10	384	11
rect	383	13	384	14
rect	383	16	384	17
rect	383	19	384	20
rect	383	22	384	23
rect	383	25	384	26
rect	383	28	384	29
rect	383	37	384	38
rect	383	40	384	41
rect	383	43	384	44
rect	383	46	384	47
rect	383	55	384	56
rect	383	64	384	65
rect	383	67	384	68
rect	383	76	384	77
rect	383	79	384	80
rect	383	85	384	86
rect	383	88	384	89
rect	383	91	384	92
rect	383	94	384	95
rect	383	97	384	98
rect	383	106	384	107
rect	383	109	384	110
rect	383	112	384	113
rect	383	115	384	116
rect	383	118	384	119
rect	383	121	384	122
rect	383	124	384	125
rect	383	127	384	128
rect	383	130	384	131
rect	383	133	384	134
rect	383	136	384	137
rect	383	145	384	146
rect	383	151	384	152
rect	383	154	384	155
rect	383	157	384	158
rect	383	160	384	161
rect	383	163	384	164
rect	383	169	384	170
rect	383	172	384	173
rect	383	178	384	179
rect	383	187	384	188
rect	383	190	384	191
rect	383	199	384	200
rect	383	208	384	209
rect	383	211	384	212
rect	383	220	384	221
rect	383	223	384	224
rect	383	226	384	227
rect	383	229	384	230
rect	383	235	384	236
rect	383	238	384	239
rect	383	241	384	242
rect	383	244	384	245
rect	383	247	384	248
rect	383	250	384	251
rect	383	253	384	254
rect	383	256	384	257
rect	383	265	384	266
rect	383	271	384	272
rect	383	277	384	278
rect	383	280	384	281
rect	383	289	384	290
rect	383	292	384	293
rect	383	295	384	296
rect	383	298	384	299
rect	383	301	384	302
rect	383	310	384	311
rect	383	319	384	320
rect	383	322	384	323
rect	383	325	384	326
rect	383	331	384	332
rect	383	352	384	353
rect	383	355	384	356
rect	383	358	384	359
rect	383	364	384	365
rect	383	367	384	368
rect	384	4	385	5
rect	384	10	385	11
rect	384	13	385	14
rect	384	16	385	17
rect	384	19	385	20
rect	384	22	385	23
rect	384	25	385	26
rect	384	28	385	29
rect	384	37	385	38
rect	384	40	385	41
rect	384	43	385	44
rect	384	46	385	47
rect	384	55	385	56
rect	384	64	385	65
rect	384	67	385	68
rect	384	76	385	77
rect	384	79	385	80
rect	384	85	385	86
rect	384	88	385	89
rect	384	91	385	92
rect	384	94	385	95
rect	384	97	385	98
rect	384	106	385	107
rect	384	109	385	110
rect	384	112	385	113
rect	384	115	385	116
rect	384	118	385	119
rect	384	121	385	122
rect	384	124	385	125
rect	384	127	385	128
rect	384	130	385	131
rect	384	133	385	134
rect	384	136	385	137
rect	384	145	385	146
rect	384	148	385	149
rect	384	151	385	152
rect	384	154	385	155
rect	384	157	385	158
rect	384	160	385	161
rect	384	163	385	164
rect	384	169	385	170
rect	384	172	385	173
rect	384	178	385	179
rect	384	187	385	188
rect	384	190	385	191
rect	384	199	385	200
rect	384	203	385	204
rect	384	208	385	209
rect	384	211	385	212
rect	384	220	385	221
rect	384	223	385	224
rect	384	226	385	227
rect	384	229	385	230
rect	384	235	385	236
rect	384	238	385	239
rect	384	241	385	242
rect	384	244	385	245
rect	384	247	385	248
rect	384	250	385	251
rect	384	253	385	254
rect	384	256	385	257
rect	384	265	385	266
rect	384	271	385	272
rect	384	277	385	278
rect	384	280	385	281
rect	384	289	385	290
rect	384	292	385	293
rect	384	295	385	296
rect	384	298	385	299
rect	384	301	385	302
rect	384	310	385	311
rect	384	319	385	320
rect	384	322	385	323
rect	384	325	385	326
rect	384	331	385	332
rect	384	352	385	353
rect	384	355	385	356
rect	384	358	385	359
rect	384	364	385	365
rect	384	367	385	368
rect	385	4	386	5
rect	385	10	386	11
rect	385	13	386	14
rect	385	16	386	17
rect	385	19	386	20
rect	385	22	386	23
rect	385	25	386	26
rect	385	28	386	29
rect	385	37	386	38
rect	385	40	386	41
rect	385	43	386	44
rect	385	46	386	47
rect	385	55	386	56
rect	385	64	386	65
rect	385	67	386	68
rect	385	76	386	77
rect	385	79	386	80
rect	385	85	386	86
rect	385	88	386	89
rect	385	91	386	92
rect	385	94	386	95
rect	385	97	386	98
rect	385	106	386	107
rect	385	109	386	110
rect	385	112	386	113
rect	385	115	386	116
rect	385	118	386	119
rect	385	121	386	122
rect	385	124	386	125
rect	385	127	386	128
rect	385	130	386	131
rect	385	133	386	134
rect	385	136	386	137
rect	385	145	386	146
rect	385	148	386	149
rect	385	151	386	152
rect	385	154	386	155
rect	385	157	386	158
rect	385	160	386	161
rect	385	169	386	170
rect	385	172	386	173
rect	385	178	386	179
rect	385	187	386	188
rect	385	190	386	191
rect	385	199	386	200
rect	385	203	386	204
rect	385	208	386	209
rect	385	211	386	212
rect	385	220	386	221
rect	385	223	386	224
rect	385	226	386	227
rect	385	229	386	230
rect	385	235	386	236
rect	385	238	386	239
rect	385	241	386	242
rect	385	244	386	245
rect	385	247	386	248
rect	385	250	386	251
rect	385	253	386	254
rect	385	256	386	257
rect	385	265	386	266
rect	385	271	386	272
rect	385	277	386	278
rect	385	289	386	290
rect	385	292	386	293
rect	385	295	386	296
rect	385	298	386	299
rect	385	301	386	302
rect	385	310	386	311
rect	385	319	386	320
rect	385	322	386	323
rect	385	325	386	326
rect	385	331	386	332
rect	385	352	386	353
rect	385	355	386	356
rect	385	358	386	359
rect	385	364	386	365
rect	385	367	386	368
rect	386	4	387	5
rect	386	10	387	11
rect	386	13	387	14
rect	386	16	387	17
rect	386	19	387	20
rect	386	22	387	23
rect	386	25	387	26
rect	386	28	387	29
rect	386	37	387	38
rect	386	40	387	41
rect	386	43	387	44
rect	386	46	387	47
rect	386	55	387	56
rect	386	64	387	65
rect	386	67	387	68
rect	386	76	387	77
rect	386	79	387	80
rect	386	85	387	86
rect	386	88	387	89
rect	386	91	387	92
rect	386	94	387	95
rect	386	97	387	98
rect	386	106	387	107
rect	386	109	387	110
rect	386	112	387	113
rect	386	115	387	116
rect	386	118	387	119
rect	386	121	387	122
rect	386	124	387	125
rect	386	127	387	128
rect	386	130	387	131
rect	386	133	387	134
rect	386	136	387	137
rect	386	145	387	146
rect	386	148	387	149
rect	386	151	387	152
rect	386	154	387	155
rect	386	157	387	158
rect	386	160	387	161
rect	386	169	387	170
rect	386	172	387	173
rect	386	175	387	176
rect	386	178	387	179
rect	386	187	387	188
rect	386	190	387	191
rect	386	199	387	200
rect	386	203	387	204
rect	386	208	387	209
rect	386	211	387	212
rect	386	220	387	221
rect	386	223	387	224
rect	386	226	387	227
rect	386	229	387	230
rect	386	235	387	236
rect	386	238	387	239
rect	386	241	387	242
rect	386	244	387	245
rect	386	247	387	248
rect	386	250	387	251
rect	386	253	387	254
rect	386	256	387	257
rect	386	265	387	266
rect	386	268	387	269
rect	386	271	387	272
rect	386	277	387	278
rect	386	289	387	290
rect	386	292	387	293
rect	386	295	387	296
rect	386	298	387	299
rect	386	301	387	302
rect	386	310	387	311
rect	386	319	387	320
rect	386	322	387	323
rect	386	325	387	326
rect	386	331	387	332
rect	386	352	387	353
rect	386	355	387	356
rect	386	358	387	359
rect	386	364	387	365
rect	386	367	387	368
rect	387	4	388	5
rect	387	10	388	11
rect	387	13	388	14
rect	387	16	388	17
rect	387	19	388	20
rect	387	22	388	23
rect	387	25	388	26
rect	387	28	388	29
rect	387	37	388	38
rect	387	40	388	41
rect	387	43	388	44
rect	387	46	388	47
rect	387	55	388	56
rect	387	64	388	65
rect	387	67	388	68
rect	387	76	388	77
rect	387	79	388	80
rect	387	85	388	86
rect	387	88	388	89
rect	387	91	388	92
rect	387	94	388	95
rect	387	97	388	98
rect	387	106	388	107
rect	387	109	388	110
rect	387	112	388	113
rect	387	115	388	116
rect	387	118	388	119
rect	387	121	388	122
rect	387	124	388	125
rect	387	127	388	128
rect	387	130	388	131
rect	387	133	388	134
rect	387	136	388	137
rect	387	145	388	146
rect	387	148	388	149
rect	387	151	388	152
rect	387	154	388	155
rect	387	160	388	161
rect	387	169	388	170
rect	387	172	388	173
rect	387	175	388	176
rect	387	178	388	179
rect	387	187	388	188
rect	387	190	388	191
rect	387	199	388	200
rect	387	203	388	204
rect	387	208	388	209
rect	387	211	388	212
rect	387	220	388	221
rect	387	223	388	224
rect	387	226	388	227
rect	387	229	388	230
rect	387	235	388	236
rect	387	238	388	239
rect	387	241	388	242
rect	387	244	388	245
rect	387	247	388	248
rect	387	250	388	251
rect	387	253	388	254
rect	387	256	388	257
rect	387	265	388	266
rect	387	268	388	269
rect	387	271	388	272
rect	387	289	388	290
rect	387	292	388	293
rect	387	295	388	296
rect	387	298	388	299
rect	387	301	388	302
rect	387	310	388	311
rect	387	319	388	320
rect	387	322	388	323
rect	387	325	388	326
rect	387	331	388	332
rect	387	352	388	353
rect	387	355	388	356
rect	387	358	388	359
rect	387	364	388	365
rect	387	367	388	368
rect	388	4	389	5
rect	388	10	389	11
rect	388	13	389	14
rect	388	16	389	17
rect	388	19	389	20
rect	388	22	389	23
rect	388	25	389	26
rect	388	28	389	29
rect	388	37	389	38
rect	388	40	389	41
rect	388	43	389	44
rect	388	46	389	47
rect	388	55	389	56
rect	388	64	389	65
rect	388	67	389	68
rect	388	76	389	77
rect	388	79	389	80
rect	388	85	389	86
rect	388	88	389	89
rect	388	91	389	92
rect	388	94	389	95
rect	388	97	389	98
rect	388	106	389	107
rect	388	109	389	110
rect	388	112	389	113
rect	388	115	389	116
rect	388	118	389	119
rect	388	121	389	122
rect	388	124	389	125
rect	388	127	389	128
rect	388	130	389	131
rect	388	133	389	134
rect	388	136	389	137
rect	388	145	389	146
rect	388	148	389	149
rect	388	151	389	152
rect	388	154	389	155
rect	388	160	389	161
rect	388	163	389	164
rect	388	169	389	170
rect	388	172	389	173
rect	388	175	389	176
rect	388	178	389	179
rect	388	187	389	188
rect	388	190	389	191
rect	388	199	389	200
rect	388	203	389	204
rect	388	208	389	209
rect	388	211	389	212
rect	388	220	389	221
rect	388	223	389	224
rect	388	226	389	227
rect	388	229	389	230
rect	388	235	389	236
rect	388	238	389	239
rect	388	241	389	242
rect	388	244	389	245
rect	388	247	389	248
rect	388	250	389	251
rect	388	253	389	254
rect	388	256	389	257
rect	388	265	389	266
rect	388	268	389	269
rect	388	271	389	272
rect	388	280	389	281
rect	388	289	389	290
rect	388	292	389	293
rect	388	295	389	296
rect	388	298	389	299
rect	388	301	389	302
rect	388	310	389	311
rect	388	319	389	320
rect	388	322	389	323
rect	388	325	389	326
rect	388	331	389	332
rect	388	352	389	353
rect	388	355	389	356
rect	388	358	389	359
rect	388	364	389	365
rect	388	367	389	368
rect	389	4	390	5
rect	389	10	390	11
rect	389	13	390	14
rect	389	16	390	17
rect	389	19	390	20
rect	389	22	390	23
rect	389	25	390	26
rect	389	28	390	29
rect	389	37	390	38
rect	389	40	390	41
rect	389	43	390	44
rect	389	46	390	47
rect	389	55	390	56
rect	389	64	390	65
rect	389	67	390	68
rect	389	76	390	77
rect	389	79	390	80
rect	389	85	390	86
rect	389	88	390	89
rect	389	91	390	92
rect	389	94	390	95
rect	389	97	390	98
rect	389	106	390	107
rect	389	109	390	110
rect	389	112	390	113
rect	389	115	390	116
rect	389	118	390	119
rect	389	121	390	122
rect	389	124	390	125
rect	389	127	390	128
rect	389	130	390	131
rect	389	133	390	134
rect	389	136	390	137
rect	389	145	390	146
rect	389	148	390	149
rect	389	151	390	152
rect	389	160	390	161
rect	389	163	390	164
rect	389	169	390	170
rect	389	172	390	173
rect	389	175	390	176
rect	389	178	390	179
rect	389	187	390	188
rect	389	190	390	191
rect	389	199	390	200
rect	389	203	390	204
rect	389	208	390	209
rect	389	211	390	212
rect	389	220	390	221
rect	389	223	390	224
rect	389	226	390	227
rect	389	229	390	230
rect	389	235	390	236
rect	389	238	390	239
rect	389	241	390	242
rect	389	244	390	245
rect	389	247	390	248
rect	389	250	390	251
rect	389	253	390	254
rect	389	256	390	257
rect	389	268	390	269
rect	389	271	390	272
rect	389	280	390	281
rect	389	289	390	290
rect	389	292	390	293
rect	389	295	390	296
rect	389	298	390	299
rect	389	301	390	302
rect	389	310	390	311
rect	389	319	390	320
rect	389	322	390	323
rect	389	325	390	326
rect	389	331	390	332
rect	389	352	390	353
rect	389	355	390	356
rect	389	358	390	359
rect	389	364	390	365
rect	389	367	390	368
rect	390	4	391	5
rect	390	10	391	11
rect	390	13	391	14
rect	390	16	391	17
rect	390	19	391	20
rect	390	22	391	23
rect	390	25	391	26
rect	390	28	391	29
rect	390	37	391	38
rect	390	40	391	41
rect	390	43	391	44
rect	390	46	391	47
rect	390	55	391	56
rect	390	64	391	65
rect	390	67	391	68
rect	390	76	391	77
rect	390	79	391	80
rect	390	85	391	86
rect	390	88	391	89
rect	390	91	391	92
rect	390	94	391	95
rect	390	97	391	98
rect	390	106	391	107
rect	390	109	391	110
rect	390	112	391	113
rect	390	115	391	116
rect	390	118	391	119
rect	390	121	391	122
rect	390	124	391	125
rect	390	127	391	128
rect	390	130	391	131
rect	390	133	391	134
rect	390	136	391	137
rect	390	145	391	146
rect	390	148	391	149
rect	390	151	391	152
rect	390	157	391	158
rect	390	160	391	161
rect	390	163	391	164
rect	390	169	391	170
rect	390	172	391	173
rect	390	175	391	176
rect	390	178	391	179
rect	390	187	391	188
rect	390	190	391	191
rect	390	199	391	200
rect	390	203	391	204
rect	390	208	391	209
rect	390	211	391	212
rect	390	220	391	221
rect	390	223	391	224
rect	390	226	391	227
rect	390	229	391	230
rect	390	235	391	236
rect	390	238	391	239
rect	390	241	391	242
rect	390	244	391	245
rect	390	247	391	248
rect	390	250	391	251
rect	390	253	391	254
rect	390	256	391	257
rect	390	268	391	269
rect	390	271	391	272
rect	390	277	391	278
rect	390	280	391	281
rect	390	289	391	290
rect	390	292	391	293
rect	390	295	391	296
rect	390	298	391	299
rect	390	301	391	302
rect	390	310	391	311
rect	390	319	391	320
rect	390	322	391	323
rect	390	325	391	326
rect	390	331	391	332
rect	390	352	391	353
rect	390	355	391	356
rect	390	358	391	359
rect	390	364	391	365
rect	390	367	391	368
rect	391	4	392	5
rect	391	10	392	11
rect	391	13	392	14
rect	391	16	392	17
rect	391	19	392	20
rect	391	22	392	23
rect	391	25	392	26
rect	391	28	392	29
rect	391	37	392	38
rect	391	40	392	41
rect	391	43	392	44
rect	391	46	392	47
rect	391	55	392	56
rect	391	64	392	65
rect	391	67	392	68
rect	391	76	392	77
rect	391	79	392	80
rect	391	85	392	86
rect	391	88	392	89
rect	391	91	392	92
rect	391	94	392	95
rect	391	97	392	98
rect	391	106	392	107
rect	391	109	392	110
rect	391	112	392	113
rect	391	115	392	116
rect	391	118	392	119
rect	391	121	392	122
rect	391	124	392	125
rect	391	127	392	128
rect	391	130	392	131
rect	391	133	392	134
rect	391	136	392	137
rect	391	148	392	149
rect	391	151	392	152
rect	391	157	392	158
rect	391	160	392	161
rect	391	163	392	164
rect	391	169	392	170
rect	391	172	392	173
rect	391	175	392	176
rect	391	178	392	179
rect	391	187	392	188
rect	391	190	392	191
rect	391	199	392	200
rect	391	208	392	209
rect	391	211	392	212
rect	391	220	392	221
rect	391	223	392	224
rect	391	226	392	227
rect	391	229	392	230
rect	391	235	392	236
rect	391	238	392	239
rect	391	241	392	242
rect	391	244	392	245
rect	391	247	392	248
rect	391	250	392	251
rect	391	253	392	254
rect	391	256	392	257
rect	391	268	392	269
rect	391	271	392	272
rect	391	277	392	278
rect	391	280	392	281
rect	391	289	392	290
rect	391	292	392	293
rect	391	295	392	296
rect	391	298	392	299
rect	391	301	392	302
rect	391	310	392	311
rect	391	319	392	320
rect	391	322	392	323
rect	391	325	392	326
rect	391	331	392	332
rect	391	352	392	353
rect	391	355	392	356
rect	391	358	392	359
rect	391	364	392	365
rect	391	367	392	368
rect	392	4	393	5
rect	392	10	393	11
rect	392	13	393	14
rect	392	16	393	17
rect	392	19	393	20
rect	392	22	393	23
rect	392	25	393	26
rect	392	28	393	29
rect	392	37	393	38
rect	392	40	393	41
rect	392	43	393	44
rect	392	46	393	47
rect	392	55	393	56
rect	392	64	393	65
rect	392	67	393	68
rect	392	76	393	77
rect	392	79	393	80
rect	392	85	393	86
rect	392	88	393	89
rect	392	91	393	92
rect	392	94	393	95
rect	392	97	393	98
rect	392	106	393	107
rect	392	109	393	110
rect	392	112	393	113
rect	392	115	393	116
rect	392	118	393	119
rect	392	121	393	122
rect	392	124	393	125
rect	392	127	393	128
rect	392	130	393	131
rect	392	133	393	134
rect	392	136	393	137
rect	392	148	393	149
rect	392	151	393	152
rect	392	154	393	155
rect	392	157	393	158
rect	392	160	393	161
rect	392	163	393	164
rect	392	169	393	170
rect	392	172	393	173
rect	392	175	393	176
rect	392	178	393	179
rect	392	187	393	188
rect	392	190	393	191
rect	392	199	393	200
rect	392	208	393	209
rect	392	211	393	212
rect	392	220	393	221
rect	392	223	393	224
rect	392	226	393	227
rect	392	229	393	230
rect	392	235	393	236
rect	392	238	393	239
rect	392	241	393	242
rect	392	244	393	245
rect	392	247	393	248
rect	392	250	393	251
rect	392	253	393	254
rect	392	256	393	257
rect	392	265	393	266
rect	392	268	393	269
rect	392	271	393	272
rect	392	277	393	278
rect	392	280	393	281
rect	392	289	393	290
rect	392	292	393	293
rect	392	295	393	296
rect	392	298	393	299
rect	392	301	393	302
rect	392	310	393	311
rect	392	319	393	320
rect	392	322	393	323
rect	392	325	393	326
rect	392	331	393	332
rect	392	352	393	353
rect	392	355	393	356
rect	392	358	393	359
rect	392	364	393	365
rect	392	367	393	368
rect	393	4	394	5
rect	393	10	394	11
rect	393	13	394	14
rect	393	16	394	17
rect	393	19	394	20
rect	393	22	394	23
rect	393	25	394	26
rect	393	28	394	29
rect	393	37	394	38
rect	393	40	394	41
rect	393	43	394	44
rect	393	46	394	47
rect	393	55	394	56
rect	393	64	394	65
rect	393	67	394	68
rect	393	76	394	77
rect	393	79	394	80
rect	393	85	394	86
rect	393	88	394	89
rect	393	91	394	92
rect	393	94	394	95
rect	393	97	394	98
rect	393	106	394	107
rect	393	109	394	110
rect	393	112	394	113
rect	393	115	394	116
rect	393	118	394	119
rect	393	121	394	122
rect	393	127	394	128
rect	393	130	394	131
rect	393	133	394	134
rect	393	136	394	137
rect	393	148	394	149
rect	393	151	394	152
rect	393	154	394	155
rect	393	157	394	158
rect	393	160	394	161
rect	393	163	394	164
rect	393	169	394	170
rect	393	172	394	173
rect	393	175	394	176
rect	393	178	394	179
rect	393	187	394	188
rect	393	190	394	191
rect	393	199	394	200
rect	393	208	394	209
rect	393	211	394	212
rect	393	220	394	221
rect	393	223	394	224
rect	393	226	394	227
rect	393	229	394	230
rect	393	235	394	236
rect	393	238	394	239
rect	393	241	394	242
rect	393	244	394	245
rect	393	247	394	248
rect	393	250	394	251
rect	393	253	394	254
rect	393	265	394	266
rect	393	268	394	269
rect	393	271	394	272
rect	393	277	394	278
rect	393	280	394	281
rect	393	289	394	290
rect	393	292	394	293
rect	393	295	394	296
rect	393	298	394	299
rect	393	301	394	302
rect	393	310	394	311
rect	393	319	394	320
rect	393	322	394	323
rect	393	325	394	326
rect	393	331	394	332
rect	393	352	394	353
rect	393	355	394	356
rect	393	358	394	359
rect	393	364	394	365
rect	393	367	394	368
rect	394	4	395	5
rect	394	10	395	11
rect	394	13	395	14
rect	394	16	395	17
rect	394	19	395	20
rect	394	22	395	23
rect	394	25	395	26
rect	394	28	395	29
rect	394	37	395	38
rect	394	40	395	41
rect	394	43	395	44
rect	394	46	395	47
rect	394	55	395	56
rect	394	64	395	65
rect	394	67	395	68
rect	394	76	395	77
rect	394	79	395	80
rect	394	85	395	86
rect	394	88	395	89
rect	394	91	395	92
rect	394	94	395	95
rect	394	97	395	98
rect	394	106	395	107
rect	394	109	395	110
rect	394	112	395	113
rect	394	115	395	116
rect	394	118	395	119
rect	394	121	395	122
rect	394	127	395	128
rect	394	130	395	131
rect	394	133	395	134
rect	394	136	395	137
rect	394	145	395	146
rect	394	148	395	149
rect	394	151	395	152
rect	394	154	395	155
rect	394	157	395	158
rect	394	160	395	161
rect	394	163	395	164
rect	394	169	395	170
rect	394	172	395	173
rect	394	175	395	176
rect	394	178	395	179
rect	394	187	395	188
rect	394	190	395	191
rect	394	199	395	200
rect	394	208	395	209
rect	394	211	395	212
rect	394	220	395	221
rect	394	223	395	224
rect	394	226	395	227
rect	394	229	395	230
rect	394	235	395	236
rect	394	238	395	239
rect	394	241	395	242
rect	394	244	395	245
rect	394	247	395	248
rect	394	250	395	251
rect	394	253	395	254
rect	394	262	395	263
rect	394	265	395	266
rect	394	268	395	269
rect	394	271	395	272
rect	394	277	395	278
rect	394	280	395	281
rect	394	289	395	290
rect	394	292	395	293
rect	394	295	395	296
rect	394	298	395	299
rect	394	301	395	302
rect	394	310	395	311
rect	394	319	395	320
rect	394	322	395	323
rect	394	325	395	326
rect	394	331	395	332
rect	394	352	395	353
rect	394	355	395	356
rect	394	358	395	359
rect	394	364	395	365
rect	394	367	395	368
rect	395	4	396	5
rect	395	10	396	11
rect	395	13	396	14
rect	395	16	396	17
rect	395	19	396	20
rect	395	22	396	23
rect	395	25	396	26
rect	395	28	396	29
rect	395	37	396	38
rect	395	40	396	41
rect	395	43	396	44
rect	395	46	396	47
rect	395	55	396	56
rect	395	64	396	65
rect	395	67	396	68
rect	395	76	396	77
rect	395	79	396	80
rect	395	85	396	86
rect	395	88	396	89
rect	395	91	396	92
rect	395	94	396	95
rect	395	97	396	98
rect	395	106	396	107
rect	395	109	396	110
rect	395	115	396	116
rect	395	118	396	119
rect	395	121	396	122
rect	395	127	396	128
rect	395	130	396	131
rect	395	133	396	134
rect	395	145	396	146
rect	395	148	396	149
rect	395	151	396	152
rect	395	154	396	155
rect	395	157	396	158
rect	395	160	396	161
rect	395	163	396	164
rect	395	169	396	170
rect	395	172	396	173
rect	395	175	396	176
rect	395	178	396	179
rect	395	187	396	188
rect	395	190	396	191
rect	395	199	396	200
rect	395	208	396	209
rect	395	211	396	212
rect	395	220	396	221
rect	395	223	396	224
rect	395	226	396	227
rect	395	229	396	230
rect	395	235	396	236
rect	395	238	396	239
rect	395	241	396	242
rect	395	244	396	245
rect	395	250	396	251
rect	395	253	396	254
rect	395	262	396	263
rect	395	265	396	266
rect	395	268	396	269
rect	395	271	396	272
rect	395	277	396	278
rect	395	280	396	281
rect	395	289	396	290
rect	395	292	396	293
rect	395	295	396	296
rect	395	298	396	299
rect	395	301	396	302
rect	395	310	396	311
rect	395	319	396	320
rect	395	322	396	323
rect	395	325	396	326
rect	395	331	396	332
rect	395	352	396	353
rect	395	355	396	356
rect	395	358	396	359
rect	395	364	396	365
rect	395	367	396	368
rect	396	4	397	5
rect	396	10	397	11
rect	396	13	397	14
rect	396	16	397	17
rect	396	19	397	20
rect	396	22	397	23
rect	396	25	397	26
rect	396	28	397	29
rect	396	37	397	38
rect	396	40	397	41
rect	396	43	397	44
rect	396	46	397	47
rect	396	55	397	56
rect	396	64	397	65
rect	396	67	397	68
rect	396	76	397	77
rect	396	79	397	80
rect	396	85	397	86
rect	396	88	397	89
rect	396	91	397	92
rect	396	94	397	95
rect	396	97	397	98
rect	396	100	397	101
rect	396	106	397	107
rect	396	109	397	110
rect	396	115	397	116
rect	396	118	397	119
rect	396	121	397	122
rect	396	124	397	125
rect	396	127	397	128
rect	396	130	397	131
rect	396	133	397	134
rect	396	145	397	146
rect	396	148	397	149
rect	396	151	397	152
rect	396	154	397	155
rect	396	157	397	158
rect	396	160	397	161
rect	396	163	397	164
rect	396	169	397	170
rect	396	172	397	173
rect	396	175	397	176
rect	396	178	397	179
rect	396	187	397	188
rect	396	190	397	191
rect	396	199	397	200
rect	396	208	397	209
rect	396	211	397	212
rect	396	220	397	221
rect	396	223	397	224
rect	396	226	397	227
rect	396	229	397	230
rect	396	235	397	236
rect	396	238	397	239
rect	396	241	397	242
rect	396	244	397	245
rect	396	250	397	251
rect	396	253	397	254
rect	396	256	397	257
rect	396	262	397	263
rect	396	265	397	266
rect	396	268	397	269
rect	396	271	397	272
rect	396	277	397	278
rect	396	280	397	281
rect	396	289	397	290
rect	396	292	397	293
rect	396	295	397	296
rect	396	298	397	299
rect	396	301	397	302
rect	396	310	397	311
rect	396	319	397	320
rect	396	322	397	323
rect	396	325	397	326
rect	396	331	397	332
rect	396	352	397	353
rect	396	355	397	356
rect	396	358	397	359
rect	396	364	397	365
rect	396	367	397	368
rect	397	4	398	5
rect	397	10	398	11
rect	397	13	398	14
rect	397	16	398	17
rect	397	19	398	20
rect	397	22	398	23
rect	397	25	398	26
rect	397	28	398	29
rect	397	37	398	38
rect	397	40	398	41
rect	397	43	398	44
rect	397	46	398	47
rect	397	55	398	56
rect	397	64	398	65
rect	397	67	398	68
rect	397	76	398	77
rect	397	79	398	80
rect	397	85	398	86
rect	397	88	398	89
rect	397	91	398	92
rect	397	94	398	95
rect	397	97	398	98
rect	397	100	398	101
rect	397	106	398	107
rect	397	109	398	110
rect	397	115	398	116
rect	397	118	398	119
rect	397	124	398	125
rect	397	130	398	131
rect	397	133	398	134
rect	397	145	398	146
rect	397	148	398	149
rect	397	151	398	152
rect	397	154	398	155
rect	397	157	398	158
rect	397	160	398	161
rect	397	163	398	164
rect	397	169	398	170
rect	397	172	398	173
rect	397	175	398	176
rect	397	178	398	179
rect	397	187	398	188
rect	397	190	398	191
rect	397	199	398	200
rect	397	208	398	209
rect	397	211	398	212
rect	397	220	398	221
rect	397	223	398	224
rect	397	226	398	227
rect	397	229	398	230
rect	397	235	398	236
rect	397	238	398	239
rect	397	244	398	245
rect	397	250	398	251
rect	397	253	398	254
rect	397	256	398	257
rect	397	262	398	263
rect	397	265	398	266
rect	397	268	398	269
rect	397	271	398	272
rect	397	277	398	278
rect	397	280	398	281
rect	397	289	398	290
rect	397	292	398	293
rect	397	295	398	296
rect	397	298	398	299
rect	397	301	398	302
rect	397	310	398	311
rect	397	319	398	320
rect	397	322	398	323
rect	397	325	398	326
rect	397	331	398	332
rect	397	352	398	353
rect	397	355	398	356
rect	397	358	398	359
rect	397	364	398	365
rect	397	367	398	368
rect	398	4	399	5
rect	398	10	399	11
rect	398	13	399	14
rect	398	16	399	17
rect	398	19	399	20
rect	398	22	399	23
rect	398	25	399	26
rect	398	28	399	29
rect	398	37	399	38
rect	398	40	399	41
rect	398	43	399	44
rect	398	46	399	47
rect	398	55	399	56
rect	398	64	399	65
rect	398	67	399	68
rect	398	76	399	77
rect	398	79	399	80
rect	398	85	399	86
rect	398	88	399	89
rect	398	91	399	92
rect	398	94	399	95
rect	398	97	399	98
rect	398	100	399	101
rect	398	106	399	107
rect	398	109	399	110
rect	398	112	399	113
rect	398	115	399	116
rect	398	118	399	119
rect	398	124	399	125
rect	398	130	399	131
rect	398	133	399	134
rect	398	136	399	137
rect	398	145	399	146
rect	398	148	399	149
rect	398	151	399	152
rect	398	154	399	155
rect	398	157	399	158
rect	398	160	399	161
rect	398	163	399	164
rect	398	169	399	170
rect	398	172	399	173
rect	398	175	399	176
rect	398	178	399	179
rect	398	187	399	188
rect	398	190	399	191
rect	398	199	399	200
rect	398	208	399	209
rect	398	211	399	212
rect	398	220	399	221
rect	398	223	399	224
rect	398	226	399	227
rect	398	229	399	230
rect	398	235	399	236
rect	398	238	399	239
rect	398	244	399	245
rect	398	247	399	248
rect	398	250	399	251
rect	398	253	399	254
rect	398	256	399	257
rect	398	262	399	263
rect	398	265	399	266
rect	398	268	399	269
rect	398	271	399	272
rect	398	277	399	278
rect	398	280	399	281
rect	398	289	399	290
rect	398	292	399	293
rect	398	295	399	296
rect	398	298	399	299
rect	398	301	399	302
rect	398	310	399	311
rect	398	319	399	320
rect	398	322	399	323
rect	398	325	399	326
rect	398	331	399	332
rect	398	352	399	353
rect	398	355	399	356
rect	398	358	399	359
rect	398	364	399	365
rect	398	367	399	368
rect	399	4	400	5
rect	399	10	400	11
rect	399	13	400	14
rect	399	16	400	17
rect	399	19	400	20
rect	399	22	400	23
rect	399	25	400	26
rect	399	28	400	29
rect	399	37	400	38
rect	399	40	400	41
rect	399	43	400	44
rect	399	46	400	47
rect	399	55	400	56
rect	399	64	400	65
rect	399	67	400	68
rect	399	76	400	77
rect	399	79	400	80
rect	399	85	400	86
rect	399	88	400	89
rect	399	91	400	92
rect	399	94	400	95
rect	399	100	400	101
rect	399	106	400	107
rect	399	109	400	110
rect	399	112	400	113
rect	399	115	400	116
rect	399	118	400	119
rect	399	124	400	125
rect	399	130	400	131
rect	399	133	400	134
rect	399	136	400	137
rect	399	145	400	146
rect	399	148	400	149
rect	399	151	400	152
rect	399	154	400	155
rect	399	157	400	158
rect	399	160	400	161
rect	399	163	400	164
rect	399	169	400	170
rect	399	172	400	173
rect	399	175	400	176
rect	399	178	400	179
rect	399	187	400	188
rect	399	190	400	191
rect	399	199	400	200
rect	399	208	400	209
rect	399	211	400	212
rect	399	220	400	221
rect	399	223	400	224
rect	399	226	400	227
rect	399	229	400	230
rect	399	235	400	236
rect	399	244	400	245
rect	399	247	400	248
rect	399	253	400	254
rect	399	256	400	257
rect	399	262	400	263
rect	399	265	400	266
rect	399	268	400	269
rect	399	271	400	272
rect	399	277	400	278
rect	399	280	400	281
rect	399	289	400	290
rect	399	292	400	293
rect	399	295	400	296
rect	399	298	400	299
rect	399	301	400	302
rect	399	310	400	311
rect	399	319	400	320
rect	399	322	400	323
rect	399	325	400	326
rect	399	331	400	332
rect	399	352	400	353
rect	399	355	400	356
rect	399	358	400	359
rect	399	364	400	365
rect	399	367	400	368
rect	400	4	401	5
rect	400	10	401	11
rect	400	13	401	14
rect	400	16	401	17
rect	400	19	401	20
rect	400	22	401	23
rect	400	25	401	26
rect	400	28	401	29
rect	400	37	401	38
rect	400	40	401	41
rect	400	43	401	44
rect	400	46	401	47
rect	400	55	401	56
rect	400	64	401	65
rect	400	67	401	68
rect	400	76	401	77
rect	400	79	401	80
rect	400	85	401	86
rect	400	88	401	89
rect	400	91	401	92
rect	400	94	401	95
rect	400	100	401	101
rect	400	106	401	107
rect	400	109	401	110
rect	400	112	401	113
rect	400	115	401	116
rect	400	118	401	119
rect	400	124	401	125
rect	400	127	401	128
rect	400	130	401	131
rect	400	133	401	134
rect	400	136	401	137
rect	400	145	401	146
rect	400	148	401	149
rect	400	151	401	152
rect	400	154	401	155
rect	400	157	401	158
rect	400	160	401	161
rect	400	163	401	164
rect	400	169	401	170
rect	400	172	401	173
rect	400	175	401	176
rect	400	178	401	179
rect	400	187	401	188
rect	400	190	401	191
rect	400	199	401	200
rect	400	208	401	209
rect	400	211	401	212
rect	400	220	401	221
rect	400	223	401	224
rect	400	226	401	227
rect	400	229	401	230
rect	400	235	401	236
rect	400	241	401	242
rect	400	244	401	245
rect	400	247	401	248
rect	400	253	401	254
rect	400	256	401	257
rect	400	259	401	260
rect	400	262	401	263
rect	400	265	401	266
rect	400	268	401	269
rect	400	271	401	272
rect	400	277	401	278
rect	400	280	401	281
rect	400	289	401	290
rect	400	292	401	293
rect	400	295	401	296
rect	400	298	401	299
rect	400	301	401	302
rect	400	310	401	311
rect	400	319	401	320
rect	400	322	401	323
rect	400	325	401	326
rect	400	331	401	332
rect	400	352	401	353
rect	400	355	401	356
rect	400	358	401	359
rect	400	364	401	365
rect	400	367	401	368
rect	401	4	402	5
rect	401	10	402	11
rect	401	13	402	14
rect	401	16	402	17
rect	401	19	402	20
rect	401	22	402	23
rect	401	25	402	26
rect	401	28	402	29
rect	401	37	402	38
rect	401	40	402	41
rect	401	43	402	44
rect	401	46	402	47
rect	401	55	402	56
rect	401	64	402	65
rect	401	67	402	68
rect	401	76	402	77
rect	401	79	402	80
rect	401	91	402	92
rect	401	94	402	95
rect	401	100	402	101
rect	401	106	402	107
rect	401	112	402	113
rect	401	115	402	116
rect	401	124	402	125
rect	401	127	402	128
rect	401	130	402	131
rect	401	133	402	134
rect	401	136	402	137
rect	401	145	402	146
rect	401	148	402	149
rect	401	151	402	152
rect	401	154	402	155
rect	401	157	402	158
rect	401	160	402	161
rect	401	163	402	164
rect	401	169	402	170
rect	401	172	402	173
rect	401	175	402	176
rect	401	178	402	179
rect	401	187	402	188
rect	401	190	402	191
rect	401	199	402	200
rect	401	208	402	209
rect	401	211	402	212
rect	401	220	402	221
rect	401	226	402	227
rect	401	229	402	230
rect	401	235	402	236
rect	401	241	402	242
rect	401	244	402	245
rect	401	247	402	248
rect	401	253	402	254
rect	401	256	402	257
rect	401	259	402	260
rect	401	262	402	263
rect	401	265	402	266
rect	401	268	402	269
rect	401	271	402	272
rect	401	277	402	278
rect	401	280	402	281
rect	401	289	402	290
rect	401	292	402	293
rect	401	295	402	296
rect	401	298	402	299
rect	401	301	402	302
rect	401	310	402	311
rect	401	319	402	320
rect	401	322	402	323
rect	401	325	402	326
rect	401	331	402	332
rect	401	352	402	353
rect	401	355	402	356
rect	401	358	402	359
rect	401	364	402	365
rect	401	367	402	368
rect	402	4	403	5
rect	402	10	403	11
rect	402	13	403	14
rect	402	16	403	17
rect	402	19	403	20
rect	402	22	403	23
rect	402	25	403	26
rect	402	28	403	29
rect	402	37	403	38
rect	402	40	403	41
rect	402	43	403	44
rect	402	46	403	47
rect	402	55	403	56
rect	402	64	403	65
rect	402	67	403	68
rect	402	76	403	77
rect	402	79	403	80
rect	402	91	403	92
rect	402	94	403	95
rect	402	97	403	98
rect	402	100	403	101
rect	402	106	403	107
rect	402	112	403	113
rect	402	115	403	116
rect	402	121	403	122
rect	402	124	403	125
rect	402	127	403	128
rect	402	130	403	131
rect	402	133	403	134
rect	402	136	403	137
rect	402	145	403	146
rect	402	148	403	149
rect	402	151	403	152
rect	402	154	403	155
rect	402	157	403	158
rect	402	160	403	161
rect	402	163	403	164
rect	402	169	403	170
rect	402	172	403	173
rect	402	175	403	176
rect	402	178	403	179
rect	402	187	403	188
rect	402	190	403	191
rect	402	199	403	200
rect	402	208	403	209
rect	402	211	403	212
rect	402	220	403	221
rect	402	226	403	227
rect	402	229	403	230
rect	402	235	403	236
rect	402	241	403	242
rect	402	244	403	245
rect	402	247	403	248
rect	402	250	403	251
rect	402	253	403	254
rect	402	256	403	257
rect	402	259	403	260
rect	402	262	403	263
rect	402	265	403	266
rect	402	268	403	269
rect	402	271	403	272
rect	402	277	403	278
rect	402	280	403	281
rect	402	289	403	290
rect	402	292	403	293
rect	402	295	403	296
rect	402	298	403	299
rect	402	301	403	302
rect	402	310	403	311
rect	402	319	403	320
rect	402	322	403	323
rect	402	325	403	326
rect	402	331	403	332
rect	402	352	403	353
rect	402	355	403	356
rect	402	358	403	359
rect	402	364	403	365
rect	402	367	403	368
rect	403	4	404	5
rect	403	10	404	11
rect	403	13	404	14
rect	403	16	404	17
rect	403	19	404	20
rect	403	22	404	23
rect	403	25	404	26
rect	403	28	404	29
rect	403	37	404	38
rect	403	40	404	41
rect	403	43	404	44
rect	403	46	404	47
rect	403	55	404	56
rect	403	64	404	65
rect	403	67	404	68
rect	403	76	404	77
rect	403	79	404	80
rect	403	94	404	95
rect	403	97	404	98
rect	403	100	404	101
rect	403	106	404	107
rect	403	112	404	113
rect	403	121	404	122
rect	403	124	404	125
rect	403	127	404	128
rect	403	130	404	131
rect	403	136	404	137
rect	403	145	404	146
rect	403	148	404	149
rect	403	151	404	152
rect	403	154	404	155
rect	403	157	404	158
rect	403	163	404	164
rect	403	169	404	170
rect	403	172	404	173
rect	403	175	404	176
rect	403	178	404	179
rect	403	187	404	188
rect	403	190	404	191
rect	403	199	404	200
rect	403	208	404	209
rect	403	211	404	212
rect	403	226	404	227
rect	403	229	404	230
rect	403	235	404	236
rect	403	241	404	242
rect	403	244	404	245
rect	403	247	404	248
rect	403	250	404	251
rect	403	253	404	254
rect	403	256	404	257
rect	403	259	404	260
rect	403	262	404	263
rect	403	265	404	266
rect	403	268	404	269
rect	403	271	404	272
rect	403	277	404	278
rect	403	280	404	281
rect	403	289	404	290
rect	403	292	404	293
rect	403	295	404	296
rect	403	298	404	299
rect	403	301	404	302
rect	403	310	404	311
rect	403	319	404	320
rect	403	322	404	323
rect	403	325	404	326
rect	403	331	404	332
rect	403	352	404	353
rect	403	355	404	356
rect	403	358	404	359
rect	403	364	404	365
rect	403	367	404	368
rect	404	4	405	5
rect	404	10	405	11
rect	404	13	405	14
rect	404	16	405	17
rect	404	19	405	20
rect	404	22	405	23
rect	404	25	405	26
rect	404	28	405	29
rect	404	37	405	38
rect	404	40	405	41
rect	404	43	405	44
rect	404	46	405	47
rect	404	55	405	56
rect	404	64	405	65
rect	404	67	405	68
rect	404	76	405	77
rect	404	79	405	80
rect	404	85	405	86
rect	404	94	405	95
rect	404	97	405	98
rect	404	100	405	101
rect	404	106	405	107
rect	404	109	405	110
rect	404	112	405	113
rect	404	118	405	119
rect	404	121	405	122
rect	404	124	405	125
rect	404	127	405	128
rect	404	130	405	131
rect	404	136	405	137
rect	404	145	405	146
rect	404	148	405	149
rect	404	151	405	152
rect	404	154	405	155
rect	404	157	405	158
rect	404	163	405	164
rect	404	166	405	167
rect	404	169	405	170
rect	404	172	405	173
rect	404	175	405	176
rect	404	178	405	179
rect	404	187	405	188
rect	404	190	405	191
rect	404	199	405	200
rect	404	208	405	209
rect	404	211	405	212
rect	404	226	405	227
rect	404	229	405	230
rect	404	235	405	236
rect	404	238	405	239
rect	404	241	405	242
rect	404	244	405	245
rect	404	247	405	248
rect	404	250	405	251
rect	404	253	405	254
rect	404	256	405	257
rect	404	259	405	260
rect	404	262	405	263
rect	404	265	405	266
rect	404	268	405	269
rect	404	271	405	272
rect	404	277	405	278
rect	404	280	405	281
rect	404	289	405	290
rect	404	292	405	293
rect	404	295	405	296
rect	404	298	405	299
rect	404	301	405	302
rect	404	310	405	311
rect	404	319	405	320
rect	404	322	405	323
rect	404	325	405	326
rect	404	331	405	332
rect	404	352	405	353
rect	404	355	405	356
rect	404	358	405	359
rect	404	364	405	365
rect	404	367	405	368
rect	405	4	406	5
rect	405	10	406	11
rect	405	13	406	14
rect	405	16	406	17
rect	405	19	406	20
rect	405	22	406	23
rect	405	28	406	29
rect	405	37	406	38
rect	405	40	406	41
rect	405	43	406	44
rect	405	46	406	47
rect	405	55	406	56
rect	405	64	406	65
rect	405	67	406	68
rect	405	76	406	77
rect	405	79	406	80
rect	405	85	406	86
rect	405	94	406	95
rect	405	97	406	98
rect	405	100	406	101
rect	405	106	406	107
rect	405	109	406	110
rect	405	112	406	113
rect	405	118	406	119
rect	405	121	406	122
rect	405	124	406	125
rect	405	127	406	128
rect	405	130	406	131
rect	405	136	406	137
rect	405	145	406	146
rect	405	148	406	149
rect	405	151	406	152
rect	405	154	406	155
rect	405	157	406	158
rect	405	163	406	164
rect	405	166	406	167
rect	405	169	406	170
rect	405	172	406	173
rect	405	175	406	176
rect	405	178	406	179
rect	405	187	406	188
rect	405	190	406	191
rect	405	199	406	200
rect	405	208	406	209
rect	405	211	406	212
rect	405	226	406	227
rect	405	229	406	230
rect	405	235	406	236
rect	405	238	406	239
rect	405	241	406	242
rect	405	244	406	245
rect	405	247	406	248
rect	405	250	406	251
rect	405	253	406	254
rect	405	256	406	257
rect	405	259	406	260
rect	405	262	406	263
rect	405	265	406	266
rect	405	268	406	269
rect	405	271	406	272
rect	405	277	406	278
rect	405	280	406	281
rect	405	289	406	290
rect	405	292	406	293
rect	405	295	406	296
rect	405	298	406	299
rect	405	301	406	302
rect	405	310	406	311
rect	405	319	406	320
rect	405	322	406	323
rect	405	325	406	326
rect	405	331	406	332
rect	405	352	406	353
rect	405	355	406	356
rect	405	358	406	359
rect	405	364	406	365
rect	405	367	406	368
rect	406	4	407	5
rect	406	10	407	11
rect	406	13	407	14
rect	406	16	407	17
rect	406	19	407	20
rect	406	22	407	23
rect	406	28	407	29
rect	406	31	407	32
rect	406	37	407	38
rect	406	40	407	41
rect	406	43	407	44
rect	406	46	407	47
rect	406	55	407	56
rect	406	64	407	65
rect	406	67	407	68
rect	406	76	407	77
rect	406	79	407	80
rect	406	85	407	86
rect	406	91	407	92
rect	406	94	407	95
rect	406	97	407	98
rect	406	100	407	101
rect	406	106	407	107
rect	406	109	407	110
rect	406	112	407	113
rect	406	118	407	119
rect	406	121	407	122
rect	406	124	407	125
rect	406	127	407	128
rect	406	130	407	131
rect	406	136	407	137
rect	406	145	407	146
rect	406	148	407	149
rect	406	151	407	152
rect	406	154	407	155
rect	406	157	407	158
rect	406	163	407	164
rect	406	166	407	167
rect	406	169	407	170
rect	406	172	407	173
rect	406	175	407	176
rect	406	178	407	179
rect	406	187	407	188
rect	406	190	407	191
rect	406	199	407	200
rect	406	208	407	209
rect	406	211	407	212
rect	406	226	407	227
rect	406	229	407	230
rect	406	235	407	236
rect	406	238	407	239
rect	406	241	407	242
rect	406	244	407	245
rect	406	247	407	248
rect	406	250	407	251
rect	406	253	407	254
rect	406	256	407	257
rect	406	259	407	260
rect	406	262	407	263
rect	406	265	407	266
rect	406	268	407	269
rect	406	271	407	272
rect	406	277	407	278
rect	406	280	407	281
rect	406	289	407	290
rect	406	292	407	293
rect	406	295	407	296
rect	406	298	407	299
rect	406	301	407	302
rect	406	307	407	308
rect	406	310	407	311
rect	406	319	407	320
rect	406	322	407	323
rect	406	325	407	326
rect	406	331	407	332
rect	406	352	407	353
rect	406	355	407	356
rect	406	358	407	359
rect	406	364	407	365
rect	406	367	407	368
rect	407	4	408	5
rect	407	10	408	11
rect	407	13	408	14
rect	407	16	408	17
rect	407	19	408	20
rect	407	22	408	23
rect	407	28	408	29
rect	407	31	408	32
rect	407	40	408	41
rect	407	46	408	47
rect	407	55	408	56
rect	407	64	408	65
rect	407	67	408	68
rect	407	76	408	77
rect	407	79	408	80
rect	407	85	408	86
rect	407	91	408	92
rect	407	94	408	95
rect	407	97	408	98
rect	407	100	408	101
rect	407	106	408	107
rect	407	109	408	110
rect	407	112	408	113
rect	407	118	408	119
rect	407	121	408	122
rect	407	124	408	125
rect	407	127	408	128
rect	407	130	408	131
rect	407	136	408	137
rect	407	145	408	146
rect	407	148	408	149
rect	407	151	408	152
rect	407	154	408	155
rect	407	157	408	158
rect	407	163	408	164
rect	407	166	408	167
rect	407	169	408	170
rect	407	172	408	173
rect	407	175	408	176
rect	407	178	408	179
rect	407	187	408	188
rect	407	190	408	191
rect	407	199	408	200
rect	407	208	408	209
rect	407	211	408	212
rect	407	226	408	227
rect	407	235	408	236
rect	407	238	408	239
rect	407	241	408	242
rect	407	244	408	245
rect	407	247	408	248
rect	407	250	408	251
rect	407	253	408	254
rect	407	256	408	257
rect	407	259	408	260
rect	407	262	408	263
rect	407	265	408	266
rect	407	268	408	269
rect	407	271	408	272
rect	407	277	408	278
rect	407	280	408	281
rect	407	289	408	290
rect	407	292	408	293
rect	407	295	408	296
rect	407	298	408	299
rect	407	301	408	302
rect	407	307	408	308
rect	407	310	408	311
rect	407	319	408	320
rect	407	322	408	323
rect	407	325	408	326
rect	407	331	408	332
rect	407	352	408	353
rect	407	355	408	356
rect	407	358	408	359
rect	407	364	408	365
rect	407	367	408	368
rect	408	4	409	5
rect	408	10	409	11
rect	408	13	409	14
rect	408	16	409	17
rect	408	19	409	20
rect	408	22	409	23
rect	408	25	409	26
rect	408	28	409	29
rect	408	31	409	32
rect	408	40	409	41
rect	408	46	409	47
rect	408	55	409	56
rect	408	64	409	65
rect	408	67	409	68
rect	408	76	409	77
rect	408	79	409	80
rect	408	85	409	86
rect	408	91	409	92
rect	408	94	409	95
rect	408	97	409	98
rect	408	100	409	101
rect	408	106	409	107
rect	408	109	409	110
rect	408	112	409	113
rect	408	118	409	119
rect	408	121	409	122
rect	408	124	409	125
rect	408	127	409	128
rect	408	130	409	131
rect	408	136	409	137
rect	408	145	409	146
rect	408	148	409	149
rect	408	151	409	152
rect	408	154	409	155
rect	408	157	409	158
rect	408	163	409	164
rect	408	166	409	167
rect	408	169	409	170
rect	408	172	409	173
rect	408	175	409	176
rect	408	178	409	179
rect	408	187	409	188
rect	408	190	409	191
rect	408	199	409	200
rect	408	208	409	209
rect	408	211	409	212
rect	408	226	409	227
rect	408	235	409	236
rect	408	238	409	239
rect	408	241	409	242
rect	408	244	409	245
rect	408	247	409	248
rect	408	250	409	251
rect	408	253	409	254
rect	408	256	409	257
rect	408	259	409	260
rect	408	262	409	263
rect	408	265	409	266
rect	408	268	409	269
rect	408	271	409	272
rect	408	277	409	278
rect	408	280	409	281
rect	408	289	409	290
rect	408	292	409	293
rect	408	295	409	296
rect	408	298	409	299
rect	408	301	409	302
rect	408	307	409	308
rect	408	310	409	311
rect	408	319	409	320
rect	408	322	409	323
rect	408	325	409	326
rect	408	331	409	332
rect	408	352	409	353
rect	408	355	409	356
rect	408	358	409	359
rect	408	364	409	365
rect	408	367	409	368
rect	409	4	410	5
rect	409	10	410	11
rect	409	13	410	14
rect	409	16	410	17
rect	409	19	410	20
rect	409	25	410	26
rect	409	28	410	29
rect	409	31	410	32
rect	409	40	410	41
rect	409	46	410	47
rect	409	67	410	68
rect	409	76	410	77
rect	409	85	410	86
rect	409	91	410	92
rect	409	94	410	95
rect	409	97	410	98
rect	409	100	410	101
rect	409	106	410	107
rect	409	109	410	110
rect	409	112	410	113
rect	409	118	410	119
rect	409	121	410	122
rect	409	124	410	125
rect	409	127	410	128
rect	409	136	410	137
rect	409	145	410	146
rect	409	148	410	149
rect	409	154	410	155
rect	409	157	410	158
rect	409	163	410	164
rect	409	166	410	167
rect	409	169	410	170
rect	409	172	410	173
rect	409	175	410	176
rect	409	178	410	179
rect	409	187	410	188
rect	409	190	410	191
rect	409	199	410	200
rect	409	208	410	209
rect	409	235	410	236
rect	409	238	410	239
rect	409	241	410	242
rect	409	244	410	245
rect	409	247	410	248
rect	409	250	410	251
rect	409	256	410	257
rect	409	259	410	260
rect	409	262	410	263
rect	409	265	410	266
rect	409	268	410	269
rect	409	271	410	272
rect	409	277	410	278
rect	409	280	410	281
rect	409	289	410	290
rect	409	292	410	293
rect	409	295	410	296
rect	409	298	410	299
rect	409	301	410	302
rect	409	307	410	308
rect	409	310	410	311
rect	409	319	410	320
rect	409	325	410	326
rect	409	331	410	332
rect	409	352	410	353
rect	409	355	410	356
rect	409	358	410	359
rect	409	364	410	365
rect	409	367	410	368
rect	410	4	411	5
rect	410	10	411	11
rect	410	13	411	14
rect	410	16	411	17
rect	410	19	411	20
rect	410	25	411	26
rect	410	28	411	29
rect	410	31	411	32
rect	410	37	411	38
rect	410	40	411	41
rect	410	46	411	47
rect	410	52	411	53
rect	410	67	411	68
rect	410	70	411	71
rect	410	76	411	77
rect	410	85	411	86
rect	410	91	411	92
rect	410	94	411	95
rect	410	97	411	98
rect	410	100	411	101
rect	410	103	411	104
rect	410	106	411	107
rect	410	109	411	110
rect	410	112	411	113
rect	410	115	411	116
rect	410	118	411	119
rect	410	121	411	122
rect	410	124	411	125
rect	410	127	411	128
rect	410	136	411	137
rect	410	145	411	146
rect	410	148	411	149
rect	410	154	411	155
rect	410	157	411	158
rect	410	160	411	161
rect	410	163	411	164
rect	410	166	411	167
rect	410	169	411	170
rect	410	172	411	173
rect	410	175	411	176
rect	410	178	411	179
rect	410	187	411	188
rect	410	190	411	191
rect	410	199	411	200
rect	410	208	411	209
rect	410	214	411	215
rect	410	217	411	218
rect	410	229	411	230
rect	410	235	411	236
rect	410	238	411	239
rect	410	241	411	242
rect	410	244	411	245
rect	410	247	411	248
rect	410	250	411	251
rect	410	256	411	257
rect	410	259	411	260
rect	410	262	411	263
rect	410	265	411	266
rect	410	268	411	269
rect	410	271	411	272
rect	410	277	411	278
rect	410	280	411	281
rect	410	289	411	290
rect	410	292	411	293
rect	410	295	411	296
rect	410	298	411	299
rect	410	301	411	302
rect	410	307	411	308
rect	410	310	411	311
rect	410	319	411	320
rect	410	325	411	326
rect	410	331	411	332
rect	410	352	411	353
rect	410	355	411	356
rect	410	358	411	359
rect	410	361	411	362
rect	410	364	411	365
rect	410	367	411	368
rect	411	4	412	5
rect	411	13	412	14
rect	411	16	412	17
rect	411	19	412	20
rect	411	25	412	26
rect	411	28	412	29
rect	411	31	412	32
rect	411	37	412	38
rect	411	40	412	41
rect	411	46	412	47
rect	411	52	412	53
rect	411	70	412	71
rect	411	76	412	77
rect	411	85	412	86
rect	411	91	412	92
rect	411	94	412	95
rect	411	97	412	98
rect	411	100	412	101
rect	411	103	412	104
rect	411	106	412	107
rect	411	109	412	110
rect	411	112	412	113
rect	411	115	412	116
rect	411	118	412	119
rect	411	121	412	122
rect	411	124	412	125
rect	411	127	412	128
rect	411	136	412	137
rect	411	145	412	146
rect	411	148	412	149
rect	411	154	412	155
rect	411	157	412	158
rect	411	160	412	161
rect	411	163	412	164
rect	411	166	412	167
rect	411	169	412	170
rect	411	172	412	173
rect	411	175	412	176
rect	411	178	412	179
rect	411	187	412	188
rect	411	190	412	191
rect	411	199	412	200
rect	411	208	412	209
rect	411	214	412	215
rect	411	217	412	218
rect	411	229	412	230
rect	411	235	412	236
rect	411	238	412	239
rect	411	241	412	242
rect	411	244	412	245
rect	411	247	412	248
rect	411	250	412	251
rect	411	256	412	257
rect	411	259	412	260
rect	411	262	412	263
rect	411	265	412	266
rect	411	268	412	269
rect	411	277	412	278
rect	411	280	412	281
rect	411	289	412	290
rect	411	295	412	296
rect	411	298	412	299
rect	411	301	412	302
rect	411	307	412	308
rect	411	310	412	311
rect	411	325	412	326
rect	411	331	412	332
rect	411	352	412	353
rect	411	355	412	356
rect	411	358	412	359
rect	411	361	412	362
rect	411	364	412	365
rect	411	367	412	368
rect	412	4	413	5
rect	412	13	413	14
rect	412	16	413	17
rect	412	19	413	20
rect	412	22	413	23
rect	412	25	413	26
rect	412	28	413	29
rect	412	31	413	32
rect	412	37	413	38
rect	412	40	413	41
rect	412	46	413	47
rect	412	52	413	53
rect	412	55	413	56
rect	412	70	413	71
rect	412	73	413	74
rect	412	76	413	77
rect	412	79	413	80
rect	412	85	413	86
rect	412	88	413	89
rect	412	91	413	92
rect	412	94	413	95
rect	412	97	413	98
rect	412	100	413	101
rect	412	103	413	104
rect	412	106	413	107
rect	412	109	413	110
rect	412	112	413	113
rect	412	115	413	116
rect	412	118	413	119
rect	412	121	413	122
rect	412	124	413	125
rect	412	127	413	128
rect	412	136	413	137
rect	412	145	413	146
rect	412	148	413	149
rect	412	154	413	155
rect	412	157	413	158
rect	412	160	413	161
rect	412	163	413	164
rect	412	166	413	167
rect	412	169	413	170
rect	412	172	413	173
rect	412	175	413	176
rect	412	178	413	179
rect	412	187	413	188
rect	412	190	413	191
rect	412	199	413	200
rect	412	208	413	209
rect	412	214	413	215
rect	412	217	413	218
rect	412	229	413	230
rect	412	235	413	236
rect	412	238	413	239
rect	412	241	413	242
rect	412	244	413	245
rect	412	247	413	248
rect	412	250	413	251
rect	412	256	413	257
rect	412	259	413	260
rect	412	262	413	263
rect	412	265	413	266
rect	412	268	413	269
rect	412	277	413	278
rect	412	280	413	281
rect	412	286	413	287
rect	412	289	413	290
rect	412	295	413	296
rect	412	298	413	299
rect	412	301	413	302
rect	412	307	413	308
rect	412	310	413	311
rect	412	322	413	323
rect	412	325	413	326
rect	412	331	413	332
rect	412	352	413	353
rect	412	355	413	356
rect	412	358	413	359
rect	412	361	413	362
rect	412	364	413	365
rect	412	367	413	368
rect	413	4	414	5
rect	413	13	414	14
rect	413	16	414	17
rect	413	22	414	23
rect	413	25	414	26
rect	413	31	414	32
rect	413	37	414	38
rect	413	40	414	41
rect	413	52	414	53
rect	413	55	414	56
rect	413	70	414	71
rect	413	73	414	74
rect	413	76	414	77
rect	413	79	414	80
rect	413	85	414	86
rect	413	88	414	89
rect	413	91	414	92
rect	413	94	414	95
rect	413	97	414	98
rect	413	100	414	101
rect	413	103	414	104
rect	413	106	414	107
rect	413	109	414	110
rect	413	112	414	113
rect	413	115	414	116
rect	413	118	414	119
rect	413	121	414	122
rect	413	124	414	125
rect	413	127	414	128
rect	413	136	414	137
rect	413	145	414	146
rect	413	148	414	149
rect	413	154	414	155
rect	413	157	414	158
rect	413	160	414	161
rect	413	163	414	164
rect	413	166	414	167
rect	413	169	414	170
rect	413	172	414	173
rect	413	175	414	176
rect	413	178	414	179
rect	413	187	414	188
rect	413	190	414	191
rect	413	199	414	200
rect	413	208	414	209
rect	413	214	414	215
rect	413	217	414	218
rect	413	229	414	230
rect	413	235	414	236
rect	413	238	414	239
rect	413	241	414	242
rect	413	244	414	245
rect	413	247	414	248
rect	413	250	414	251
rect	413	256	414	257
rect	413	259	414	260
rect	413	262	414	263
rect	413	265	414	266
rect	413	268	414	269
rect	413	277	414	278
rect	413	280	414	281
rect	413	286	414	287
rect	413	289	414	290
rect	413	295	414	296
rect	413	298	414	299
rect	413	301	414	302
rect	413	307	414	308
rect	413	310	414	311
rect	413	322	414	323
rect	413	325	414	326
rect	413	331	414	332
rect	413	352	414	353
rect	413	355	414	356
rect	413	361	414	362
rect	413	364	414	365
rect	413	367	414	368
rect	414	4	415	5
rect	414	10	415	11
rect	414	13	415	14
rect	414	16	415	17
rect	414	22	415	23
rect	414	25	415	26
rect	414	31	415	32
rect	414	37	415	38
rect	414	40	415	41
rect	414	43	415	44
rect	414	52	415	53
rect	414	55	415	56
rect	414	70	415	71
rect	414	73	415	74
rect	414	76	415	77
rect	414	79	415	80
rect	414	85	415	86
rect	414	88	415	89
rect	414	91	415	92
rect	414	94	415	95
rect	414	97	415	98
rect	414	100	415	101
rect	414	103	415	104
rect	414	106	415	107
rect	414	109	415	110
rect	414	112	415	113
rect	414	115	415	116
rect	414	118	415	119
rect	414	121	415	122
rect	414	124	415	125
rect	414	127	415	128
rect	414	136	415	137
rect	414	145	415	146
rect	414	148	415	149
rect	414	154	415	155
rect	414	157	415	158
rect	414	160	415	161
rect	414	163	415	164
rect	414	166	415	167
rect	414	169	415	170
rect	414	172	415	173
rect	414	175	415	176
rect	414	178	415	179
rect	414	187	415	188
rect	414	190	415	191
rect	414	199	415	200
rect	414	208	415	209
rect	414	214	415	215
rect	414	217	415	218
rect	414	229	415	230
rect	414	235	415	236
rect	414	238	415	239
rect	414	241	415	242
rect	414	244	415	245
rect	414	247	415	248
rect	414	250	415	251
rect	414	256	415	257
rect	414	259	415	260
rect	414	262	415	263
rect	414	265	415	266
rect	414	268	415	269
rect	414	277	415	278
rect	414	280	415	281
rect	414	286	415	287
rect	414	289	415	290
rect	414	295	415	296
rect	414	298	415	299
rect	414	301	415	302
rect	414	307	415	308
rect	414	310	415	311
rect	414	322	415	323
rect	414	325	415	326
rect	414	331	415	332
rect	414	352	415	353
rect	414	355	415	356
rect	414	361	415	362
rect	414	364	415	365
rect	414	367	415	368
rect	415	4	416	5
rect	415	10	416	11
rect	415	13	416	14
rect	415	22	416	23
rect	415	25	416	26
rect	415	31	416	32
rect	415	37	416	38
rect	415	40	416	41
rect	415	43	416	44
rect	415	52	416	53
rect	415	55	416	56
rect	415	70	416	71
rect	415	73	416	74
rect	415	76	416	77
rect	415	79	416	80
rect	415	85	416	86
rect	415	88	416	89
rect	415	91	416	92
rect	415	94	416	95
rect	415	97	416	98
rect	415	100	416	101
rect	415	103	416	104
rect	415	106	416	107
rect	415	109	416	110
rect	415	112	416	113
rect	415	115	416	116
rect	415	118	416	119
rect	415	121	416	122
rect	415	124	416	125
rect	415	127	416	128
rect	415	136	416	137
rect	415	145	416	146
rect	415	148	416	149
rect	415	154	416	155
rect	415	157	416	158
rect	415	160	416	161
rect	415	163	416	164
rect	415	166	416	167
rect	415	169	416	170
rect	415	172	416	173
rect	415	175	416	176
rect	415	178	416	179
rect	415	187	416	188
rect	415	190	416	191
rect	415	199	416	200
rect	415	208	416	209
rect	415	214	416	215
rect	415	217	416	218
rect	415	229	416	230
rect	415	235	416	236
rect	415	238	416	239
rect	415	241	416	242
rect	415	247	416	248
rect	415	250	416	251
rect	415	256	416	257
rect	415	259	416	260
rect	415	262	416	263
rect	415	265	416	266
rect	415	268	416	269
rect	415	277	416	278
rect	415	280	416	281
rect	415	286	416	287
rect	415	295	416	296
rect	415	298	416	299
rect	415	301	416	302
rect	415	307	416	308
rect	415	310	416	311
rect	415	322	416	323
rect	415	331	416	332
rect	415	352	416	353
rect	415	355	416	356
rect	415	361	416	362
rect	415	364	416	365
rect	415	367	416	368
rect	416	4	417	5
rect	416	7	417	8
rect	416	10	417	11
rect	416	13	417	14
rect	416	19	417	20
rect	416	22	417	23
rect	416	25	417	26
rect	416	28	417	29
rect	416	31	417	32
rect	416	34	417	35
rect	416	37	417	38
rect	416	40	417	41
rect	416	43	417	44
rect	416	52	417	53
rect	416	55	417	56
rect	416	70	417	71
rect	416	73	417	74
rect	416	76	417	77
rect	416	79	417	80
rect	416	85	417	86
rect	416	88	417	89
rect	416	91	417	92
rect	416	94	417	95
rect	416	97	417	98
rect	416	100	417	101
rect	416	103	417	104
rect	416	106	417	107
rect	416	109	417	110
rect	416	112	417	113
rect	416	115	417	116
rect	416	118	417	119
rect	416	121	417	122
rect	416	124	417	125
rect	416	127	417	128
rect	416	136	417	137
rect	416	145	417	146
rect	416	148	417	149
rect	416	154	417	155
rect	416	157	417	158
rect	416	160	417	161
rect	416	163	417	164
rect	416	166	417	167
rect	416	169	417	170
rect	416	172	417	173
rect	416	175	417	176
rect	416	178	417	179
rect	416	187	417	188
rect	416	190	417	191
rect	416	199	417	200
rect	416	208	417	209
rect	416	214	417	215
rect	416	217	417	218
rect	416	229	417	230
rect	416	232	417	233
rect	416	235	417	236
rect	416	238	417	239
rect	416	241	417	242
rect	416	247	417	248
rect	416	250	417	251
rect	416	253	417	254
rect	416	256	417	257
rect	416	259	417	260
rect	416	262	417	263
rect	416	265	417	266
rect	416	268	417	269
rect	416	277	417	278
rect	416	280	417	281
rect	416	286	417	287
rect	416	292	417	293
rect	416	295	417	296
rect	416	298	417	299
rect	416	301	417	302
rect	416	307	417	308
rect	416	310	417	311
rect	416	313	417	314
rect	416	322	417	323
rect	416	331	417	332
rect	416	352	417	353
rect	416	355	417	356
rect	416	361	417	362
rect	416	364	417	365
rect	416	367	417	368
rect	417	7	418	8
rect	417	10	418	11
rect	417	13	418	14
rect	417	19	418	20
rect	417	22	418	23
rect	417	25	418	26
rect	417	28	418	29
rect	417	31	418	32
rect	417	34	418	35
rect	417	37	418	38
rect	417	40	418	41
rect	417	43	418	44
rect	417	52	418	53
rect	417	55	418	56
rect	417	70	418	71
rect	417	73	418	74
rect	417	79	418	80
rect	417	85	418	86
rect	417	88	418	89
rect	417	91	418	92
rect	417	94	418	95
rect	417	97	418	98
rect	417	100	418	101
rect	417	103	418	104
rect	417	106	418	107
rect	417	109	418	110
rect	417	112	418	113
rect	417	115	418	116
rect	417	118	418	119
rect	417	121	418	122
rect	417	124	418	125
rect	417	127	418	128
rect	417	136	418	137
rect	417	145	418	146
rect	417	148	418	149
rect	417	154	418	155
rect	417	157	418	158
rect	417	160	418	161
rect	417	163	418	164
rect	417	166	418	167
rect	417	169	418	170
rect	417	172	418	173
rect	417	175	418	176
rect	417	178	418	179
rect	417	187	418	188
rect	417	190	418	191
rect	417	199	418	200
rect	417	214	418	215
rect	417	217	418	218
rect	417	229	418	230
rect	417	232	418	233
rect	417	238	418	239
rect	417	241	418	242
rect	417	247	418	248
rect	417	250	418	251
rect	417	253	418	254
rect	417	256	418	257
rect	417	259	418	260
rect	417	262	418	263
rect	417	265	418	266
rect	417	268	418	269
rect	417	277	418	278
rect	417	280	418	281
rect	417	286	418	287
rect	417	292	418	293
rect	417	295	418	296
rect	417	301	418	302
rect	417	307	418	308
rect	417	313	418	314
rect	417	322	418	323
rect	417	331	418	332
rect	417	352	418	353
rect	417	355	418	356
rect	417	361	418	362
rect	417	364	418	365
rect	417	367	418	368
rect	418	7	419	8
rect	418	10	419	11
rect	418	13	419	14
rect	418	19	419	20
rect	418	22	419	23
rect	418	25	419	26
rect	418	28	419	29
rect	418	31	419	32
rect	418	34	419	35
rect	418	37	419	38
rect	418	40	419	41
rect	418	43	419	44
rect	418	52	419	53
rect	418	55	419	56
rect	418	70	419	71
rect	418	73	419	74
rect	418	79	419	80
rect	418	82	419	83
rect	418	85	419	86
rect	418	88	419	89
rect	418	91	419	92
rect	418	94	419	95
rect	418	97	419	98
rect	418	100	419	101
rect	418	103	419	104
rect	418	106	419	107
rect	418	109	419	110
rect	418	112	419	113
rect	418	115	419	116
rect	418	118	419	119
rect	418	121	419	122
rect	418	124	419	125
rect	418	127	419	128
rect	418	136	419	137
rect	418	145	419	146
rect	418	148	419	149
rect	418	154	419	155
rect	418	157	419	158
rect	418	160	419	161
rect	418	163	419	164
rect	418	166	419	167
rect	418	169	419	170
rect	418	172	419	173
rect	418	175	419	176
rect	418	178	419	179
rect	418	187	419	188
rect	418	190	419	191
rect	418	199	419	200
rect	418	205	419	206
rect	418	214	419	215
rect	418	217	419	218
rect	418	226	419	227
rect	418	229	419	230
rect	418	232	419	233
rect	418	238	419	239
rect	418	241	419	242
rect	418	244	419	245
rect	418	247	419	248
rect	418	250	419	251
rect	418	253	419	254
rect	418	256	419	257
rect	418	259	419	260
rect	418	262	419	263
rect	418	265	419	266
rect	418	268	419	269
rect	418	277	419	278
rect	418	280	419	281
rect	418	283	419	284
rect	418	286	419	287
rect	418	292	419	293
rect	418	295	419	296
rect	418	301	419	302
rect	418	307	419	308
rect	418	313	419	314
rect	418	322	419	323
rect	418	325	419	326
rect	418	331	419	332
rect	418	352	419	353
rect	418	355	419	356
rect	418	361	419	362
rect	418	364	419	365
rect	418	367	419	368
rect	419	7	420	8
rect	419	10	420	11
rect	419	13	420	14
rect	419	19	420	20
rect	419	22	420	23
rect	419	25	420	26
rect	419	28	420	29
rect	419	31	420	32
rect	419	34	420	35
rect	419	37	420	38
rect	419	40	420	41
rect	419	43	420	44
rect	419	52	420	53
rect	419	55	420	56
rect	419	70	420	71
rect	419	73	420	74
rect	419	79	420	80
rect	419	82	420	83
rect	419	85	420	86
rect	419	88	420	89
rect	419	91	420	92
rect	419	94	420	95
rect	419	97	420	98
rect	419	100	420	101
rect	419	103	420	104
rect	419	106	420	107
rect	419	109	420	110
rect	419	112	420	113
rect	419	115	420	116
rect	419	118	420	119
rect	419	121	420	122
rect	419	124	420	125
rect	419	127	420	128
rect	419	136	420	137
rect	419	145	420	146
rect	419	148	420	149
rect	419	154	420	155
rect	419	157	420	158
rect	419	160	420	161
rect	419	163	420	164
rect	419	166	420	167
rect	419	169	420	170
rect	419	172	420	173
rect	419	175	420	176
rect	419	178	420	179
rect	419	187	420	188
rect	419	190	420	191
rect	419	199	420	200
rect	419	205	420	206
rect	419	214	420	215
rect	419	217	420	218
rect	419	226	420	227
rect	419	229	420	230
rect	419	232	420	233
rect	419	238	420	239
rect	419	241	420	242
rect	419	244	420	245
rect	419	247	420	248
rect	419	250	420	251
rect	419	253	420	254
rect	419	256	420	257
rect	419	259	420	260
rect	419	262	420	263
rect	419	265	420	266
rect	419	268	420	269
rect	419	277	420	278
rect	419	280	420	281
rect	419	283	420	284
rect	419	286	420	287
rect	419	292	420	293
rect	419	301	420	302
rect	419	307	420	308
rect	419	313	420	314
rect	419	322	420	323
rect	419	325	420	326
rect	419	355	420	356
rect	419	361	420	362
rect	419	364	420	365
rect	419	367	420	368
rect	420	1	421	2
rect	420	7	421	8
rect	420	10	421	11
rect	420	13	421	14
rect	420	19	421	20
rect	420	22	421	23
rect	420	25	421	26
rect	420	28	421	29
rect	420	31	421	32
rect	420	34	421	35
rect	420	37	421	38
rect	420	40	421	41
rect	420	43	421	44
rect	420	52	421	53
rect	420	55	421	56
rect	420	70	421	71
rect	420	73	421	74
rect	420	79	421	80
rect	420	82	421	83
rect	420	85	421	86
rect	420	88	421	89
rect	420	91	421	92
rect	420	94	421	95
rect	420	97	421	98
rect	420	100	421	101
rect	420	103	421	104
rect	420	106	421	107
rect	420	109	421	110
rect	420	112	421	113
rect	420	115	421	116
rect	420	118	421	119
rect	420	121	421	122
rect	420	124	421	125
rect	420	127	421	128
rect	420	136	421	137
rect	420	145	421	146
rect	420	148	421	149
rect	420	154	421	155
rect	420	157	421	158
rect	420	160	421	161
rect	420	163	421	164
rect	420	166	421	167
rect	420	169	421	170
rect	420	172	421	173
rect	420	175	421	176
rect	420	178	421	179
rect	420	187	421	188
rect	420	190	421	191
rect	420	199	421	200
rect	420	205	421	206
rect	420	214	421	215
rect	420	217	421	218
rect	420	226	421	227
rect	420	229	421	230
rect	420	232	421	233
rect	420	238	421	239
rect	420	241	421	242
rect	420	244	421	245
rect	420	247	421	248
rect	420	250	421	251
rect	420	253	421	254
rect	420	256	421	257
rect	420	259	421	260
rect	420	262	421	263
rect	420	265	421	266
rect	420	268	421	269
rect	420	277	421	278
rect	420	280	421	281
rect	420	283	421	284
rect	420	286	421	287
rect	420	292	421	293
rect	420	301	421	302
rect	420	307	421	308
rect	420	310	421	311
rect	420	313	421	314
rect	420	319	421	320
rect	420	322	421	323
rect	420	325	421	326
rect	420	334	421	335
rect	420	349	421	350
rect	420	355	421	356
rect	420	361	421	362
rect	420	364	421	365
rect	420	367	421	368
rect	427	4	428	5
rect	427	7	428	8
rect	427	10	428	11
rect	427	13	428	14
rect	427	22	428	23
rect	427	25	428	26
rect	427	28	428	29
rect	427	31	428	32
rect	427	34	428	35
rect	427	37	428	38
rect	427	40	428	41
rect	427	43	428	44
rect	427	52	428	53
rect	427	55	428	56
rect	427	70	428	71
rect	427	73	428	74
rect	427	76	428	77
rect	427	82	428	83
rect	427	85	428	86
rect	427	88	428	89
rect	427	91	428	92
rect	427	94	428	95
rect	427	97	428	98
rect	427	100	428	101
rect	427	103	428	104
rect	427	106	428	107
rect	427	109	428	110
rect	427	112	428	113
rect	427	115	428	116
rect	427	118	428	119
rect	427	121	428	122
rect	427	124	428	125
rect	427	127	428	128
rect	427	130	428	131
rect	427	136	428	137
rect	427	145	428	146
rect	427	148	428	149
rect	427	157	428	158
rect	427	160	428	161
rect	427	163	428	164
rect	427	166	428	167
rect	427	169	428	170
rect	427	172	428	173
rect	427	175	428	176
rect	427	178	428	179
rect	427	184	428	185
rect	427	187	428	188
rect	427	190	428	191
rect	427	199	428	200
rect	427	202	428	203
rect	427	214	428	215
rect	427	217	428	218
rect	427	226	428	227
rect	427	229	428	230
rect	427	235	428	236
rect	427	238	428	239
rect	427	241	428	242
rect	427	244	428	245
rect	427	247	428	248
rect	427	250	428	251
rect	427	253	428	254
rect	427	256	428	257
rect	427	259	428	260
rect	427	262	428	263
rect	427	265	428	266
rect	427	268	428	269
rect	427	271	428	272
rect	427	277	428	278
rect	427	280	428	281
rect	427	283	428	284
rect	427	286	428	287
rect	427	292	428	293
rect	427	301	428	302
rect	427	310	428	311
rect	427	313	428	314
rect	427	322	428	323
rect	427	325	428	326
rect	427	331	428	332
rect	427	334	428	335
rect	427	349	428	350
rect	427	355	428	356
rect	427	358	428	359
rect	427	364	428	365
rect	427	367	428	368
rect	428	4	429	5
rect	428	7	429	8
rect	428	10	429	11
rect	428	13	429	14
rect	428	22	429	23
rect	428	25	429	26
rect	428	28	429	29
rect	428	31	429	32
rect	428	34	429	35
rect	428	37	429	38
rect	428	40	429	41
rect	428	43	429	44
rect	428	52	429	53
rect	428	55	429	56
rect	428	70	429	71
rect	428	73	429	74
rect	428	76	429	77
rect	428	82	429	83
rect	428	85	429	86
rect	428	88	429	89
rect	428	91	429	92
rect	428	94	429	95
rect	428	100	429	101
rect	428	103	429	104
rect	428	106	429	107
rect	428	109	429	110
rect	428	112	429	113
rect	428	115	429	116
rect	428	118	429	119
rect	428	121	429	122
rect	428	124	429	125
rect	428	127	429	128
rect	428	130	429	131
rect	428	136	429	137
rect	428	145	429	146
rect	428	148	429	149
rect	428	157	429	158
rect	428	160	429	161
rect	428	163	429	164
rect	428	166	429	167
rect	428	169	429	170
rect	428	172	429	173
rect	428	175	429	176
rect	428	178	429	179
rect	428	184	429	185
rect	428	187	429	188
rect	428	190	429	191
rect	428	199	429	200
rect	428	202	429	203
rect	428	214	429	215
rect	428	217	429	218
rect	428	226	429	227
rect	428	229	429	230
rect	428	235	429	236
rect	428	238	429	239
rect	428	241	429	242
rect	428	244	429	245
rect	428	247	429	248
rect	428	250	429	251
rect	428	253	429	254
rect	428	256	429	257
rect	428	259	429	260
rect	428	262	429	263
rect	428	265	429	266
rect	428	268	429	269
rect	428	271	429	272
rect	428	277	429	278
rect	428	280	429	281
rect	428	283	429	284
rect	428	286	429	287
rect	428	292	429	293
rect	428	301	429	302
rect	428	310	429	311
rect	428	313	429	314
rect	428	322	429	323
rect	428	325	429	326
rect	428	331	429	332
rect	428	334	429	335
rect	428	349	429	350
rect	428	355	429	356
rect	428	358	429	359
rect	428	364	429	365
rect	428	367	429	368
rect	429	4	430	5
rect	429	7	430	8
rect	429	10	430	11
rect	429	13	430	14
rect	429	22	430	23
rect	429	25	430	26
rect	429	28	430	29
rect	429	31	430	32
rect	429	34	430	35
rect	429	37	430	38
rect	429	40	430	41
rect	429	43	430	44
rect	429	52	430	53
rect	429	55	430	56
rect	429	70	430	71
rect	429	73	430	74
rect	429	76	430	77
rect	429	79	430	80
rect	429	82	430	83
rect	429	85	430	86
rect	429	88	430	89
rect	429	91	430	92
rect	429	94	430	95
rect	429	100	430	101
rect	429	103	430	104
rect	429	106	430	107
rect	429	109	430	110
rect	429	112	430	113
rect	429	115	430	116
rect	429	118	430	119
rect	429	121	430	122
rect	429	124	430	125
rect	429	127	430	128
rect	429	130	430	131
rect	429	136	430	137
rect	429	145	430	146
rect	429	148	430	149
rect	429	157	430	158
rect	429	160	430	161
rect	429	163	430	164
rect	429	166	430	167
rect	429	169	430	170
rect	429	172	430	173
rect	429	175	430	176
rect	429	178	430	179
rect	429	184	430	185
rect	429	187	430	188
rect	429	190	430	191
rect	429	199	430	200
rect	429	202	430	203
rect	429	214	430	215
rect	429	217	430	218
rect	429	226	430	227
rect	429	229	430	230
rect	429	235	430	236
rect	429	238	430	239
rect	429	241	430	242
rect	429	244	430	245
rect	429	247	430	248
rect	429	250	430	251
rect	429	253	430	254
rect	429	256	430	257
rect	429	259	430	260
rect	429	262	430	263
rect	429	265	430	266
rect	429	268	430	269
rect	429	271	430	272
rect	429	277	430	278
rect	429	280	430	281
rect	429	283	430	284
rect	429	286	430	287
rect	429	292	430	293
rect	429	301	430	302
rect	429	310	430	311
rect	429	313	430	314
rect	429	322	430	323
rect	429	325	430	326
rect	429	331	430	332
rect	429	334	430	335
rect	429	349	430	350
rect	429	355	430	356
rect	429	358	430	359
rect	429	364	430	365
rect	429	367	430	368
rect	430	4	431	5
rect	430	7	431	8
rect	430	10	431	11
rect	430	13	431	14
rect	430	22	431	23
rect	430	25	431	26
rect	430	28	431	29
rect	430	31	431	32
rect	430	34	431	35
rect	430	37	431	38
rect	430	40	431	41
rect	430	43	431	44
rect	430	52	431	53
rect	430	55	431	56
rect	430	70	431	71
rect	430	73	431	74
rect	430	79	431	80
rect	430	82	431	83
rect	430	85	431	86
rect	430	88	431	89
rect	430	91	431	92
rect	430	94	431	95
rect	430	100	431	101
rect	430	103	431	104
rect	430	106	431	107
rect	430	109	431	110
rect	430	112	431	113
rect	430	115	431	116
rect	430	118	431	119
rect	430	121	431	122
rect	430	124	431	125
rect	430	127	431	128
rect	430	130	431	131
rect	430	136	431	137
rect	430	145	431	146
rect	430	148	431	149
rect	430	157	431	158
rect	430	160	431	161
rect	430	163	431	164
rect	430	166	431	167
rect	430	169	431	170
rect	430	172	431	173
rect	430	175	431	176
rect	430	178	431	179
rect	430	184	431	185
rect	430	187	431	188
rect	430	190	431	191
rect	430	199	431	200
rect	430	202	431	203
rect	430	214	431	215
rect	430	217	431	218
rect	430	226	431	227
rect	430	229	431	230
rect	430	235	431	236
rect	430	238	431	239
rect	430	241	431	242
rect	430	244	431	245
rect	430	247	431	248
rect	430	250	431	251
rect	430	253	431	254
rect	430	256	431	257
rect	430	259	431	260
rect	430	262	431	263
rect	430	268	431	269
rect	430	271	431	272
rect	430	277	431	278
rect	430	280	431	281
rect	430	283	431	284
rect	430	286	431	287
rect	430	292	431	293
rect	430	301	431	302
rect	430	310	431	311
rect	430	313	431	314
rect	430	322	431	323
rect	430	325	431	326
rect	430	331	431	332
rect	430	334	431	335
rect	430	349	431	350
rect	430	355	431	356
rect	430	358	431	359
rect	430	364	431	365
rect	430	367	431	368
rect	431	4	432	5
rect	431	7	432	8
rect	431	10	432	11
rect	431	13	432	14
rect	431	22	432	23
rect	431	25	432	26
rect	431	28	432	29
rect	431	31	432	32
rect	431	34	432	35
rect	431	37	432	38
rect	431	40	432	41
rect	431	43	432	44
rect	431	52	432	53
rect	431	55	432	56
rect	431	70	432	71
rect	431	73	432	74
rect	431	79	432	80
rect	431	82	432	83
rect	431	85	432	86
rect	431	88	432	89
rect	431	91	432	92
rect	431	94	432	95
rect	431	100	432	101
rect	431	103	432	104
rect	431	106	432	107
rect	431	109	432	110
rect	431	112	432	113
rect	431	115	432	116
rect	431	118	432	119
rect	431	121	432	122
rect	431	124	432	125
rect	431	127	432	128
rect	431	130	432	131
rect	431	136	432	137
rect	431	145	432	146
rect	431	148	432	149
rect	431	157	432	158
rect	431	160	432	161
rect	431	163	432	164
rect	431	166	432	167
rect	431	169	432	170
rect	431	172	432	173
rect	431	175	432	176
rect	431	178	432	179
rect	431	184	432	185
rect	431	187	432	188
rect	431	190	432	191
rect	431	199	432	200
rect	431	202	432	203
rect	431	214	432	215
rect	431	217	432	218
rect	431	226	432	227
rect	431	229	432	230
rect	431	235	432	236
rect	431	238	432	239
rect	431	241	432	242
rect	431	244	432	245
rect	431	247	432	248
rect	431	250	432	251
rect	431	253	432	254
rect	431	256	432	257
rect	431	259	432	260
rect	431	262	432	263
rect	431	268	432	269
rect	431	271	432	272
rect	431	277	432	278
rect	431	280	432	281
rect	431	283	432	284
rect	431	286	432	287
rect	431	292	432	293
rect	431	301	432	302
rect	431	310	432	311
rect	431	313	432	314
rect	431	322	432	323
rect	431	325	432	326
rect	431	331	432	332
rect	431	334	432	335
rect	431	349	432	350
rect	431	355	432	356
rect	431	358	432	359
rect	431	364	432	365
rect	431	367	432	368
rect	432	4	433	5
rect	432	7	433	8
rect	432	10	433	11
rect	432	13	433	14
rect	432	22	433	23
rect	432	25	433	26
rect	432	28	433	29
rect	432	31	433	32
rect	432	34	433	35
rect	432	37	433	38
rect	432	40	433	41
rect	432	43	433	44
rect	432	52	433	53
rect	432	55	433	56
rect	432	70	433	71
rect	432	73	433	74
rect	432	79	433	80
rect	432	82	433	83
rect	432	85	433	86
rect	432	88	433	89
rect	432	91	433	92
rect	432	100	433	101
rect	432	103	433	104
rect	432	106	433	107
rect	432	109	433	110
rect	432	112	433	113
rect	432	115	433	116
rect	432	118	433	119
rect	432	121	433	122
rect	432	124	433	125
rect	432	127	433	128
rect	432	130	433	131
rect	432	136	433	137
rect	432	145	433	146
rect	432	148	433	149
rect	432	157	433	158
rect	432	160	433	161
rect	432	163	433	164
rect	432	166	433	167
rect	432	169	433	170
rect	432	172	433	173
rect	432	175	433	176
rect	432	178	433	179
rect	432	184	433	185
rect	432	187	433	188
rect	432	190	433	191
rect	432	199	433	200
rect	432	202	433	203
rect	432	214	433	215
rect	432	217	433	218
rect	432	226	433	227
rect	432	229	433	230
rect	432	238	433	239
rect	432	244	433	245
rect	432	247	433	248
rect	432	250	433	251
rect	432	253	433	254
rect	432	256	433	257
rect	432	259	433	260
rect	432	262	433	263
rect	432	268	433	269
rect	432	271	433	272
rect	432	277	433	278
rect	432	280	433	281
rect	432	283	433	284
rect	432	286	433	287
rect	432	292	433	293
rect	432	301	433	302
rect	432	310	433	311
rect	432	313	433	314
rect	432	322	433	323
rect	432	325	433	326
rect	432	331	433	332
rect	432	334	433	335
rect	432	349	433	350
rect	432	355	433	356
rect	432	358	433	359
rect	432	364	433	365
rect	432	367	433	368
rect	433	4	434	5
rect	433	7	434	8
rect	433	10	434	11
rect	433	13	434	14
rect	433	22	434	23
rect	433	25	434	26
rect	433	28	434	29
rect	433	31	434	32
rect	433	34	434	35
rect	433	37	434	38
rect	433	40	434	41
rect	433	43	434	44
rect	433	52	434	53
rect	433	55	434	56
rect	433	70	434	71
rect	433	73	434	74
rect	433	76	434	77
rect	433	79	434	80
rect	433	82	434	83
rect	433	85	434	86
rect	433	88	434	89
rect	433	91	434	92
rect	433	100	434	101
rect	433	103	434	104
rect	433	106	434	107
rect	433	109	434	110
rect	433	112	434	113
rect	433	115	434	116
rect	433	118	434	119
rect	433	121	434	122
rect	433	124	434	125
rect	433	127	434	128
rect	433	130	434	131
rect	433	136	434	137
rect	433	145	434	146
rect	433	148	434	149
rect	433	157	434	158
rect	433	160	434	161
rect	433	163	434	164
rect	433	166	434	167
rect	433	169	434	170
rect	433	172	434	173
rect	433	175	434	176
rect	433	178	434	179
rect	433	184	434	185
rect	433	187	434	188
rect	433	190	434	191
rect	433	199	434	200
rect	433	202	434	203
rect	433	214	434	215
rect	433	217	434	218
rect	433	226	434	227
rect	433	229	434	230
rect	433	238	434	239
rect	433	244	434	245
rect	433	247	434	248
rect	433	250	434	251
rect	433	253	434	254
rect	433	256	434	257
rect	433	259	434	260
rect	433	262	434	263
rect	433	268	434	269
rect	433	271	434	272
rect	433	277	434	278
rect	433	280	434	281
rect	433	283	434	284
rect	433	286	434	287
rect	433	292	434	293
rect	433	301	434	302
rect	433	310	434	311
rect	433	313	434	314
rect	433	322	434	323
rect	433	325	434	326
rect	433	331	434	332
rect	433	334	434	335
rect	433	349	434	350
rect	433	355	434	356
rect	433	358	434	359
rect	433	364	434	365
rect	433	367	434	368
rect	434	4	435	5
rect	434	7	435	8
rect	434	10	435	11
rect	434	13	435	14
rect	434	22	435	23
rect	434	25	435	26
rect	434	28	435	29
rect	434	31	435	32
rect	434	34	435	35
rect	434	40	435	41
rect	434	43	435	44
rect	434	52	435	53
rect	434	55	435	56
rect	434	70	435	71
rect	434	73	435	74
rect	434	76	435	77
rect	434	79	435	80
rect	434	82	435	83
rect	434	85	435	86
rect	434	88	435	89
rect	434	91	435	92
rect	434	100	435	101
rect	434	103	435	104
rect	434	106	435	107
rect	434	109	435	110
rect	434	112	435	113
rect	434	115	435	116
rect	434	118	435	119
rect	434	121	435	122
rect	434	124	435	125
rect	434	127	435	128
rect	434	136	435	137
rect	434	145	435	146
rect	434	148	435	149
rect	434	157	435	158
rect	434	163	435	164
rect	434	166	435	167
rect	434	169	435	170
rect	434	172	435	173
rect	434	175	435	176
rect	434	178	435	179
rect	434	184	435	185
rect	434	187	435	188
rect	434	190	435	191
rect	434	199	435	200
rect	434	202	435	203
rect	434	214	435	215
rect	434	217	435	218
rect	434	226	435	227
rect	434	229	435	230
rect	434	238	435	239
rect	434	244	435	245
rect	434	250	435	251
rect	434	253	435	254
rect	434	256	435	257
rect	434	259	435	260
rect	434	262	435	263
rect	434	268	435	269
rect	434	271	435	272
rect	434	277	435	278
rect	434	280	435	281
rect	434	283	435	284
rect	434	286	435	287
rect	434	292	435	293
rect	434	301	435	302
rect	434	310	435	311
rect	434	313	435	314
rect	434	322	435	323
rect	434	325	435	326
rect	434	331	435	332
rect	434	334	435	335
rect	434	349	435	350
rect	434	355	435	356
rect	434	358	435	359
rect	434	364	435	365
rect	434	367	435	368
rect	435	4	436	5
rect	435	7	436	8
rect	435	10	436	11
rect	435	13	436	14
rect	435	22	436	23
rect	435	25	436	26
rect	435	28	436	29
rect	435	31	436	32
rect	435	34	436	35
rect	435	40	436	41
rect	435	43	436	44
rect	435	52	436	53
rect	435	55	436	56
rect	435	70	436	71
rect	435	73	436	74
rect	435	76	436	77
rect	435	79	436	80
rect	435	82	436	83
rect	435	85	436	86
rect	435	88	436	89
rect	435	91	436	92
rect	435	100	436	101
rect	435	103	436	104
rect	435	106	436	107
rect	435	109	436	110
rect	435	112	436	113
rect	435	115	436	116
rect	435	118	436	119
rect	435	121	436	122
rect	435	124	436	125
rect	435	127	436	128
rect	435	136	436	137
rect	435	145	436	146
rect	435	148	436	149
rect	435	154	436	155
rect	435	157	436	158
rect	435	163	436	164
rect	435	166	436	167
rect	435	169	436	170
rect	435	172	436	173
rect	435	175	436	176
rect	435	178	436	179
rect	435	184	436	185
rect	435	187	436	188
rect	435	190	436	191
rect	435	199	436	200
rect	435	202	436	203
rect	435	214	436	215
rect	435	217	436	218
rect	435	226	436	227
rect	435	229	436	230
rect	435	235	436	236
rect	435	238	436	239
rect	435	244	436	245
rect	435	250	436	251
rect	435	253	436	254
rect	435	256	436	257
rect	435	259	436	260
rect	435	262	436	263
rect	435	268	436	269
rect	435	271	436	272
rect	435	277	436	278
rect	435	280	436	281
rect	435	283	436	284
rect	435	286	436	287
rect	435	292	436	293
rect	435	301	436	302
rect	435	310	436	311
rect	435	313	436	314
rect	435	322	436	323
rect	435	325	436	326
rect	435	331	436	332
rect	435	334	436	335
rect	435	349	436	350
rect	435	355	436	356
rect	435	358	436	359
rect	435	364	436	365
rect	435	367	436	368
rect	436	4	437	5
rect	436	7	437	8
rect	436	10	437	11
rect	436	13	437	14
rect	436	25	437	26
rect	436	28	437	29
rect	436	31	437	32
rect	436	34	437	35
rect	436	40	437	41
rect	436	43	437	44
rect	436	52	437	53
rect	436	55	437	56
rect	436	70	437	71
rect	436	73	437	74
rect	436	76	437	77
rect	436	79	437	80
rect	436	85	437	86
rect	436	88	437	89
rect	436	91	437	92
rect	436	100	437	101
rect	436	103	437	104
rect	436	109	437	110
rect	436	112	437	113
rect	436	115	437	116
rect	436	118	437	119
rect	436	121	437	122
rect	436	124	437	125
rect	436	127	437	128
rect	436	136	437	137
rect	436	145	437	146
rect	436	148	437	149
rect	436	154	437	155
rect	436	157	437	158
rect	436	166	437	167
rect	436	169	437	170
rect	436	172	437	173
rect	436	175	437	176
rect	436	178	437	179
rect	436	184	437	185
rect	436	187	437	188
rect	436	190	437	191
rect	436	199	437	200
rect	436	202	437	203
rect	436	214	437	215
rect	436	217	437	218
rect	436	226	437	227
rect	436	229	437	230
rect	436	235	437	236
rect	436	238	437	239
rect	436	250	437	251
rect	436	253	437	254
rect	436	256	437	257
rect	436	259	437	260
rect	436	262	437	263
rect	436	268	437	269
rect	436	271	437	272
rect	436	277	437	278
rect	436	280	437	281
rect	436	283	437	284
rect	436	286	437	287
rect	436	292	437	293
rect	436	301	437	302
rect	436	310	437	311
rect	436	313	437	314
rect	436	322	437	323
rect	436	325	437	326
rect	436	331	437	332
rect	436	334	437	335
rect	436	349	437	350
rect	436	355	437	356
rect	436	358	437	359
rect	436	364	437	365
rect	436	367	437	368
rect	437	4	438	5
rect	437	7	438	8
rect	437	10	438	11
rect	437	13	438	14
rect	437	25	438	26
rect	437	28	438	29
rect	437	31	438	32
rect	437	34	438	35
rect	437	37	438	38
rect	437	40	438	41
rect	437	43	438	44
rect	437	52	438	53
rect	437	55	438	56
rect	437	64	438	65
rect	437	70	438	71
rect	437	73	438	74
rect	437	76	438	77
rect	437	79	438	80
rect	437	85	438	86
rect	437	88	438	89
rect	437	91	438	92
rect	437	100	438	101
rect	437	103	438	104
rect	437	109	438	110
rect	437	112	438	113
rect	437	115	438	116
rect	437	118	438	119
rect	437	121	438	122
rect	437	124	438	125
rect	437	127	438	128
rect	437	130	438	131
rect	437	136	438	137
rect	437	142	438	143
rect	437	145	438	146
rect	437	148	438	149
rect	437	154	438	155
rect	437	157	438	158
rect	437	166	438	167
rect	437	169	438	170
rect	437	172	438	173
rect	437	175	438	176
rect	437	178	438	179
rect	437	184	438	185
rect	437	187	438	188
rect	437	190	438	191
rect	437	199	438	200
rect	437	202	438	203
rect	437	214	438	215
rect	437	217	438	218
rect	437	226	438	227
rect	437	229	438	230
rect	437	235	438	236
rect	437	238	438	239
rect	437	247	438	248
rect	437	250	438	251
rect	437	253	438	254
rect	437	256	438	257
rect	437	259	438	260
rect	437	262	438	263
rect	437	268	438	269
rect	437	271	438	272
rect	437	277	438	278
rect	437	280	438	281
rect	437	283	438	284
rect	437	286	438	287
rect	437	292	438	293
rect	437	301	438	302
rect	437	310	438	311
rect	437	313	438	314
rect	437	322	438	323
rect	437	325	438	326
rect	437	331	438	332
rect	437	334	438	335
rect	437	349	438	350
rect	437	355	438	356
rect	437	358	438	359
rect	437	364	438	365
rect	437	367	438	368
rect	438	4	439	5
rect	438	7	439	8
rect	438	10	439	11
rect	438	13	439	14
rect	438	25	439	26
rect	438	31	439	32
rect	438	34	439	35
rect	438	37	439	38
rect	438	40	439	41
rect	438	43	439	44
rect	438	52	439	53
rect	438	55	439	56
rect	438	64	439	65
rect	438	70	439	71
rect	438	76	439	77
rect	438	79	439	80
rect	438	85	439	86
rect	438	88	439	89
rect	438	91	439	92
rect	438	100	439	101
rect	438	103	439	104
rect	438	109	439	110
rect	438	112	439	113
rect	438	115	439	116
rect	438	118	439	119
rect	438	121	439	122
rect	438	127	439	128
rect	438	130	439	131
rect	438	136	439	137
rect	438	142	439	143
rect	438	148	439	149
rect	438	154	439	155
rect	438	157	439	158
rect	438	166	439	167
rect	438	169	439	170
rect	438	172	439	173
rect	438	175	439	176
rect	438	184	439	185
rect	438	187	439	188
rect	438	190	439	191
rect	438	199	439	200
rect	438	202	439	203
rect	438	214	439	215
rect	438	217	439	218
rect	438	226	439	227
rect	438	229	439	230
rect	438	235	439	236
rect	438	247	439	248
rect	438	250	439	251
rect	438	253	439	254
rect	438	256	439	257
rect	438	259	439	260
rect	438	262	439	263
rect	438	268	439	269
rect	438	271	439	272
rect	438	280	439	281
rect	438	283	439	284
rect	438	292	439	293
rect	438	301	439	302
rect	438	313	439	314
rect	438	322	439	323
rect	438	325	439	326
rect	438	331	439	332
rect	438	334	439	335
rect	438	349	439	350
rect	438	355	439	356
rect	438	358	439	359
rect	438	364	439	365
rect	438	367	439	368
rect	439	4	440	5
rect	439	7	440	8
rect	439	10	440	11
rect	439	13	440	14
rect	439	22	440	23
rect	439	25	440	26
rect	439	31	440	32
rect	439	34	440	35
rect	439	37	440	38
rect	439	40	440	41
rect	439	43	440	44
rect	439	52	440	53
rect	439	55	440	56
rect	439	64	440	65
rect	439	70	440	71
rect	439	76	440	77
rect	439	79	440	80
rect	439	82	440	83
rect	439	85	440	86
rect	439	88	440	89
rect	439	91	440	92
rect	439	97	440	98
rect	439	100	440	101
rect	439	103	440	104
rect	439	109	440	110
rect	439	112	440	113
rect	439	115	440	116
rect	439	118	440	119
rect	439	121	440	122
rect	439	127	440	128
rect	439	130	440	131
rect	439	136	440	137
rect	439	142	440	143
rect	439	148	440	149
rect	439	154	440	155
rect	439	157	440	158
rect	439	160	440	161
rect	439	163	440	164
rect	439	166	440	167
rect	439	169	440	170
rect	439	172	440	173
rect	439	175	440	176
rect	439	184	440	185
rect	439	187	440	188
rect	439	190	440	191
rect	439	199	440	200
rect	439	202	440	203
rect	439	214	440	215
rect	439	217	440	218
rect	439	226	440	227
rect	439	229	440	230
rect	439	235	440	236
rect	439	244	440	245
rect	439	247	440	248
rect	439	250	440	251
rect	439	253	440	254
rect	439	256	440	257
rect	439	259	440	260
rect	439	262	440	263
rect	439	268	440	269
rect	439	271	440	272
rect	439	280	440	281
rect	439	283	440	284
rect	439	292	440	293
rect	439	298	440	299
rect	439	301	440	302
rect	439	313	440	314
rect	439	322	440	323
rect	439	325	440	326
rect	439	331	440	332
rect	439	334	440	335
rect	439	349	440	350
rect	439	355	440	356
rect	439	358	440	359
rect	439	364	440	365
rect	439	367	440	368
rect	440	4	441	5
rect	440	7	441	8
rect	440	10	441	11
rect	440	13	441	14
rect	440	22	441	23
rect	440	25	441	26
rect	440	31	441	32
rect	440	34	441	35
rect	440	37	441	38
rect	440	40	441	41
rect	440	52	441	53
rect	440	55	441	56
rect	440	64	441	65
rect	440	76	441	77
rect	440	79	441	80
rect	440	82	441	83
rect	440	85	441	86
rect	440	88	441	89
rect	440	97	441	98
rect	440	100	441	101
rect	440	103	441	104
rect	440	109	441	110
rect	440	112	441	113
rect	440	118	441	119
rect	440	121	441	122
rect	440	127	441	128
rect	440	130	441	131
rect	440	136	441	137
rect	440	142	441	143
rect	440	148	441	149
rect	440	154	441	155
rect	440	157	441	158
rect	440	160	441	161
rect	440	163	441	164
rect	440	166	441	167
rect	440	169	441	170
rect	440	175	441	176
rect	440	184	441	185
rect	440	187	441	188
rect	440	199	441	200
rect	440	202	441	203
rect	440	214	441	215
rect	440	217	441	218
rect	440	226	441	227
rect	440	229	441	230
rect	440	235	441	236
rect	440	244	441	245
rect	440	247	441	248
rect	440	250	441	251
rect	440	256	441	257
rect	440	259	441	260
rect	440	262	441	263
rect	440	268	441	269
rect	440	271	441	272
rect	440	280	441	281
rect	440	283	441	284
rect	440	292	441	293
rect	440	298	441	299
rect	440	313	441	314
rect	440	322	441	323
rect	440	325	441	326
rect	440	331	441	332
rect	440	349	441	350
rect	440	355	441	356
rect	440	358	441	359
rect	440	364	441	365
rect	440	367	441	368
rect	441	4	442	5
rect	441	7	442	8
rect	441	10	442	11
rect	441	13	442	14
rect	441	22	442	23
rect	441	25	442	26
rect	441	28	442	29
rect	441	31	442	32
rect	441	34	442	35
rect	441	37	442	38
rect	441	40	442	41
rect	441	52	442	53
rect	441	55	442	56
rect	441	64	442	65
rect	441	67	442	68
rect	441	73	442	74
rect	441	76	442	77
rect	441	79	442	80
rect	441	82	442	83
rect	441	85	442	86
rect	441	88	442	89
rect	441	94	442	95
rect	441	97	442	98
rect	441	100	442	101
rect	441	103	442	104
rect	441	109	442	110
rect	441	112	442	113
rect	441	118	442	119
rect	441	121	442	122
rect	441	127	442	128
rect	441	130	442	131
rect	441	136	442	137
rect	441	142	442	143
rect	441	145	442	146
rect	441	148	442	149
rect	441	154	442	155
rect	441	157	442	158
rect	441	160	442	161
rect	441	163	442	164
rect	441	166	442	167
rect	441	169	442	170
rect	441	175	442	176
rect	441	178	442	179
rect	441	184	442	185
rect	441	187	442	188
rect	441	199	442	200
rect	441	202	442	203
rect	441	214	442	215
rect	441	217	442	218
rect	441	226	442	227
rect	441	229	442	230
rect	441	235	442	236
rect	441	238	442	239
rect	441	244	442	245
rect	441	247	442	248
rect	441	250	442	251
rect	441	256	442	257
rect	441	259	442	260
rect	441	262	442	263
rect	441	268	442	269
rect	441	271	442	272
rect	441	280	442	281
rect	441	283	442	284
rect	441	286	442	287
rect	441	292	442	293
rect	441	298	442	299
rect	441	310	442	311
rect	441	313	442	314
rect	441	322	442	323
rect	441	325	442	326
rect	441	331	442	332
rect	441	349	442	350
rect	441	355	442	356
rect	441	358	442	359
rect	441	364	442	365
rect	441	367	442	368
rect	442	4	443	5
rect	442	7	443	8
rect	442	10	443	11
rect	442	13	443	14
rect	442	22	443	23
rect	442	25	443	26
rect	442	28	443	29
rect	442	31	443	32
rect	442	34	443	35
rect	442	37	443	38
rect	442	40	443	41
rect	442	52	443	53
rect	442	64	443	65
rect	442	67	443	68
rect	442	73	443	74
rect	442	76	443	77
rect	442	79	443	80
rect	442	82	443	83
rect	442	85	443	86
rect	442	94	443	95
rect	442	97	443	98
rect	442	100	443	101
rect	442	103	443	104
rect	442	109	443	110
rect	442	118	443	119
rect	442	127	443	128
rect	442	130	443	131
rect	442	136	443	137
rect	442	142	443	143
rect	442	145	443	146
rect	442	148	443	149
rect	442	154	443	155
rect	442	157	443	158
rect	442	160	443	161
rect	442	163	443	164
rect	442	166	443	167
rect	442	169	443	170
rect	442	175	443	176
rect	442	178	443	179
rect	442	184	443	185
rect	442	187	443	188
rect	442	199	443	200
rect	442	202	443	203
rect	442	214	443	215
rect	442	217	443	218
rect	442	226	443	227
rect	442	229	443	230
rect	442	235	443	236
rect	442	238	443	239
rect	442	244	443	245
rect	442	247	443	248
rect	442	250	443	251
rect	442	256	443	257
rect	442	259	443	260
rect	442	262	443	263
rect	442	268	443	269
rect	442	271	443	272
rect	442	280	443	281
rect	442	283	443	284
rect	442	286	443	287
rect	442	292	443	293
rect	442	298	443	299
rect	442	310	443	311
rect	442	313	443	314
rect	442	322	443	323
rect	442	325	443	326
rect	442	331	443	332
rect	442	349	443	350
rect	442	355	443	356
rect	442	358	443	359
rect	442	364	443	365
rect	442	367	443	368
rect	443	4	444	5
rect	443	7	444	8
rect	443	10	444	11
rect	443	13	444	14
rect	443	22	444	23
rect	443	25	444	26
rect	443	28	444	29
rect	443	31	444	32
rect	443	34	444	35
rect	443	37	444	38
rect	443	40	444	41
rect	443	43	444	44
rect	443	52	444	53
rect	443	64	444	65
rect	443	67	444	68
rect	443	70	444	71
rect	443	73	444	74
rect	443	76	444	77
rect	443	79	444	80
rect	443	82	444	83
rect	443	85	444	86
rect	443	91	444	92
rect	443	94	444	95
rect	443	97	444	98
rect	443	100	444	101
rect	443	103	444	104
rect	443	109	444	110
rect	443	118	444	119
rect	443	127	444	128
rect	443	130	444	131
rect	443	136	444	137
rect	443	142	444	143
rect	443	145	444	146
rect	443	148	444	149
rect	443	154	444	155
rect	443	157	444	158
rect	443	160	444	161
rect	443	163	444	164
rect	443	166	444	167
rect	443	169	444	170
rect	443	175	444	176
rect	443	178	444	179
rect	443	184	444	185
rect	443	187	444	188
rect	443	199	444	200
rect	443	202	444	203
rect	443	214	444	215
rect	443	217	444	218
rect	443	226	444	227
rect	443	229	444	230
rect	443	235	444	236
rect	443	238	444	239
rect	443	244	444	245
rect	443	247	444	248
rect	443	250	444	251
rect	443	256	444	257
rect	443	259	444	260
rect	443	262	444	263
rect	443	268	444	269
rect	443	271	444	272
rect	443	280	444	281
rect	443	283	444	284
rect	443	286	444	287
rect	443	292	444	293
rect	443	298	444	299
rect	443	310	444	311
rect	443	313	444	314
rect	443	322	444	323
rect	443	325	444	326
rect	443	331	444	332
rect	443	334	444	335
rect	443	349	444	350
rect	443	355	444	356
rect	443	358	444	359
rect	443	364	444	365
rect	443	367	444	368
rect	444	7	445	8
rect	444	10	445	11
rect	444	13	445	14
rect	444	22	445	23
rect	444	25	445	26
rect	444	28	445	29
rect	444	31	445	32
rect	444	34	445	35
rect	444	37	445	38
rect	444	40	445	41
rect	444	43	445	44
rect	444	52	445	53
rect	444	64	445	65
rect	444	67	445	68
rect	444	70	445	71
rect	444	73	445	74
rect	444	76	445	77
rect	444	79	445	80
rect	444	82	445	83
rect	444	85	445	86
rect	444	91	445	92
rect	444	94	445	95
rect	444	97	445	98
rect	444	100	445	101
rect	444	103	445	104
rect	444	109	445	110
rect	444	118	445	119
rect	444	127	445	128
rect	444	130	445	131
rect	444	136	445	137
rect	444	142	445	143
rect	444	145	445	146
rect	444	148	445	149
rect	444	154	445	155
rect	444	157	445	158
rect	444	160	445	161
rect	444	163	445	164
rect	444	166	445	167
rect	444	169	445	170
rect	444	175	445	176
rect	444	178	445	179
rect	444	184	445	185
rect	444	187	445	188
rect	444	199	445	200
rect	444	202	445	203
rect	444	214	445	215
rect	444	217	445	218
rect	444	226	445	227
rect	444	229	445	230
rect	444	235	445	236
rect	444	238	445	239
rect	444	244	445	245
rect	444	247	445	248
rect	444	250	445	251
rect	444	256	445	257
rect	444	259	445	260
rect	444	262	445	263
rect	444	268	445	269
rect	444	271	445	272
rect	444	280	445	281
rect	444	283	445	284
rect	444	286	445	287
rect	444	292	445	293
rect	444	298	445	299
rect	444	310	445	311
rect	444	313	445	314
rect	444	322	445	323
rect	444	325	445	326
rect	444	331	445	332
rect	444	334	445	335
rect	444	349	445	350
rect	444	355	445	356
rect	444	358	445	359
rect	444	364	445	365
rect	445	7	446	8
rect	445	10	446	11
rect	445	13	446	14
rect	445	22	446	23
rect	445	25	446	26
rect	445	28	446	29
rect	445	31	446	32
rect	445	34	446	35
rect	445	37	446	38
rect	445	40	446	41
rect	445	43	446	44
rect	445	52	446	53
rect	445	64	446	65
rect	445	67	446	68
rect	445	70	446	71
rect	445	73	446	74
rect	445	76	446	77
rect	445	79	446	80
rect	445	82	446	83
rect	445	85	446	86
rect	445	91	446	92
rect	445	94	446	95
rect	445	97	446	98
rect	445	100	446	101
rect	445	103	446	104
rect	445	109	446	110
rect	445	118	446	119
rect	445	127	446	128
rect	445	130	446	131
rect	445	136	446	137
rect	445	142	446	143
rect	445	145	446	146
rect	445	148	446	149
rect	445	154	446	155
rect	445	157	446	158
rect	445	160	446	161
rect	445	163	446	164
rect	445	166	446	167
rect	445	169	446	170
rect	445	175	446	176
rect	445	178	446	179
rect	445	184	446	185
rect	445	187	446	188
rect	445	199	446	200
rect	445	202	446	203
rect	445	214	446	215
rect	445	217	446	218
rect	445	226	446	227
rect	445	229	446	230
rect	445	235	446	236
rect	445	238	446	239
rect	445	244	446	245
rect	445	247	446	248
rect	445	250	446	251
rect	445	256	446	257
rect	445	259	446	260
rect	445	262	446	263
rect	445	268	446	269
rect	445	271	446	272
rect	445	280	446	281
rect	445	283	446	284
rect	445	286	446	287
rect	445	292	446	293
rect	445	298	446	299
rect	445	310	446	311
rect	445	313	446	314
rect	445	322	446	323
rect	445	325	446	326
rect	445	331	446	332
rect	445	334	446	335
rect	445	349	446	350
rect	445	355	446	356
rect	445	358	446	359
rect	445	364	446	365
rect	446	10	447	11
rect	446	13	447	14
rect	446	22	447	23
rect	446	25	447	26
rect	446	28	447	29
rect	446	31	447	32
rect	446	34	447	35
rect	446	37	447	38
rect	446	43	447	44
rect	446	52	447	53
rect	446	64	447	65
rect	446	67	447	68
rect	446	70	447	71
rect	446	73	447	74
rect	446	76	447	77
rect	446	79	447	80
rect	446	82	447	83
rect	446	85	447	86
rect	446	91	447	92
rect	446	94	447	95
rect	446	97	447	98
rect	446	100	447	101
rect	446	103	447	104
rect	446	118	447	119
rect	446	130	447	131
rect	446	136	447	137
rect	446	142	447	143
rect	446	145	447	146
rect	446	154	447	155
rect	446	157	447	158
rect	446	160	447	161
rect	446	163	447	164
rect	446	166	447	167
rect	446	169	447	170
rect	446	178	447	179
rect	446	184	447	185
rect	446	187	447	188
rect	446	202	447	203
rect	446	214	447	215
rect	446	226	447	227
rect	446	235	447	236
rect	446	238	447	239
rect	446	244	447	245
rect	446	247	447	248
rect	446	256	447	257
rect	446	259	447	260
rect	446	262	447	263
rect	446	268	447	269
rect	446	271	447	272
rect	446	280	447	281
rect	446	283	447	284
rect	446	286	447	287
rect	446	298	447	299
rect	446	310	447	311
rect	446	322	447	323
rect	446	331	447	332
rect	446	334	447	335
rect	446	349	447	350
rect	446	355	447	356
rect	446	358	447	359
rect	446	364	447	365
rect	447	4	448	5
rect	447	10	448	11
rect	447	13	448	14
rect	447	22	448	23
rect	447	25	448	26
rect	447	28	448	29
rect	447	31	448	32
rect	447	34	448	35
rect	447	37	448	38
rect	447	43	448	44
rect	447	52	448	53
rect	447	55	448	56
rect	447	64	448	65
rect	447	67	448	68
rect	447	70	448	71
rect	447	73	448	74
rect	447	76	448	77
rect	447	79	448	80
rect	447	82	448	83
rect	447	85	448	86
rect	447	88	448	89
rect	447	91	448	92
rect	447	94	448	95
rect	447	97	448	98
rect	447	100	448	101
rect	447	103	448	104
rect	447	112	448	113
rect	447	118	448	119
rect	447	130	448	131
rect	447	133	448	134
rect	447	136	448	137
rect	447	142	448	143
rect	447	145	448	146
rect	447	154	448	155
rect	447	157	448	158
rect	447	160	448	161
rect	447	163	448	164
rect	447	166	448	167
rect	447	169	448	170
rect	447	178	448	179
rect	447	181	448	182
rect	447	184	448	185
rect	447	187	448	188
rect	447	196	448	197
rect	447	202	448	203
rect	447	214	448	215
rect	447	220	448	221
rect	447	226	448	227
rect	447	232	448	233
rect	447	235	448	236
rect	447	238	448	239
rect	447	244	448	245
rect	447	247	448	248
rect	447	253	448	254
rect	447	256	448	257
rect	447	259	448	260
rect	447	262	448	263
rect	447	268	448	269
rect	447	271	448	272
rect	447	277	448	278
rect	447	280	448	281
rect	447	283	448	284
rect	447	286	448	287
rect	447	298	448	299
rect	447	301	448	302
rect	447	310	448	311
rect	447	316	448	317
rect	447	322	448	323
rect	447	331	448	332
rect	447	334	448	335
rect	447	349	448	350
rect	447	355	448	356
rect	447	358	448	359
rect	447	364	448	365
rect	448	4	449	5
rect	448	13	449	14
rect	448	22	449	23
rect	448	28	449	29
rect	448	34	449	35
rect	448	37	449	38
rect	448	43	449	44
rect	448	52	449	53
rect	448	55	449	56
rect	448	64	449	65
rect	448	67	449	68
rect	448	70	449	71
rect	448	73	449	74
rect	448	76	449	77
rect	448	79	449	80
rect	448	82	449	83
rect	448	88	449	89
rect	448	91	449	92
rect	448	94	449	95
rect	448	97	449	98
rect	448	100	449	101
rect	448	103	449	104
rect	448	112	449	113
rect	448	130	449	131
rect	448	133	449	134
rect	448	136	449	137
rect	448	142	449	143
rect	448	145	449	146
rect	448	154	449	155
rect	448	160	449	161
rect	448	163	449	164
rect	448	169	449	170
rect	448	178	449	179
rect	448	181	449	182
rect	448	196	449	197
rect	448	202	449	203
rect	448	220	449	221
rect	448	232	449	233
rect	448	235	449	236
rect	448	238	449	239
rect	448	244	449	245
rect	448	247	449	248
rect	448	253	449	254
rect	448	256	449	257
rect	448	259	449	260
rect	448	262	449	263
rect	448	268	449	269
rect	448	271	449	272
rect	448	277	449	278
rect	448	280	449	281
rect	448	286	449	287
rect	448	298	449	299
rect	448	301	449	302
rect	448	310	449	311
rect	448	316	449	317
rect	448	322	449	323
rect	448	334	449	335
rect	448	349	449	350
rect	448	355	449	356
rect	448	358	449	359
rect	449	4	450	5
rect	449	7	450	8
rect	449	13	450	14
rect	449	19	450	20
rect	449	22	450	23
rect	449	28	450	29
rect	449	34	450	35
rect	449	37	450	38
rect	449	40	450	41
rect	449	43	450	44
rect	449	52	450	53
rect	449	55	450	56
rect	449	64	450	65
rect	449	67	450	68
rect	449	70	450	71
rect	449	73	450	74
rect	449	76	450	77
rect	449	79	450	80
rect	449	82	450	83
rect	449	88	450	89
rect	449	91	450	92
rect	449	94	450	95
rect	449	97	450	98
rect	449	100	450	101
rect	449	103	450	104
rect	449	106	450	107
rect	449	109	450	110
rect	449	112	450	113
rect	449	121	450	122
rect	449	130	450	131
rect	449	133	450	134
rect	449	136	450	137
rect	449	142	450	143
rect	449	145	450	146
rect	449	154	450	155
rect	449	160	450	161
rect	449	163	450	164
rect	449	169	450	170
rect	449	175	450	176
rect	449	178	450	179
rect	449	181	450	182
rect	449	190	450	191
rect	449	196	450	197
rect	449	202	450	203
rect	449	211	450	212
rect	449	217	450	218
rect	449	220	450	221
rect	449	229	450	230
rect	449	232	450	233
rect	449	235	450	236
rect	449	238	450	239
rect	449	244	450	245
rect	449	247	450	248
rect	449	250	450	251
rect	449	253	450	254
rect	449	256	450	257
rect	449	259	450	260
rect	449	262	450	263
rect	449	268	450	269
rect	449	271	450	272
rect	449	277	450	278
rect	449	280	450	281
rect	449	286	450	287
rect	449	295	450	296
rect	449	298	450	299
rect	449	301	450	302
rect	449	304	450	305
rect	449	310	450	311
rect	449	313	450	314
rect	449	316	450	317
rect	449	322	450	323
rect	449	334	450	335
rect	449	346	450	347
rect	449	349	450	350
rect	449	355	450	356
rect	449	358	450	359
rect	450	4	451	5
rect	450	7	451	8
rect	450	19	451	20
rect	450	22	451	23
rect	450	28	451	29
rect	450	37	451	38
rect	450	40	451	41
rect	450	43	451	44
rect	450	52	451	53
rect	450	55	451	56
rect	450	64	451	65
rect	450	67	451	68
rect	450	70	451	71
rect	450	73	451	74
rect	450	76	451	77
rect	450	79	451	80
rect	450	82	451	83
rect	450	88	451	89
rect	450	91	451	92
rect	450	94	451	95
rect	450	97	451	98
rect	450	106	451	107
rect	450	109	451	110
rect	450	112	451	113
rect	450	121	451	122
rect	450	130	451	131
rect	450	133	451	134
rect	450	142	451	143
rect	450	145	451	146
rect	450	154	451	155
rect	450	160	451	161
rect	450	163	451	164
rect	450	175	451	176
rect	450	178	451	179
rect	450	181	451	182
rect	450	190	451	191
rect	450	196	451	197
rect	450	211	451	212
rect	450	217	451	218
rect	450	220	451	221
rect	450	229	451	230
rect	450	232	451	233
rect	450	235	451	236
rect	450	238	451	239
rect	450	244	451	245
rect	450	247	451	248
rect	450	250	451	251
rect	450	253	451	254
rect	450	256	451	257
rect	450	259	451	260
rect	450	268	451	269
rect	450	277	451	278
rect	450	286	451	287
rect	450	295	451	296
rect	450	298	451	299
rect	450	301	451	302
rect	450	304	451	305
rect	450	310	451	311
rect	450	313	451	314
rect	450	316	451	317
rect	450	334	451	335
rect	450	346	451	347
rect	451	4	452	5
rect	451	7	452	8
rect	451	10	452	11
rect	451	19	452	20
rect	451	22	452	23
rect	451	25	452	26
rect	451	28	452	29
rect	451	37	452	38
rect	451	40	452	41
rect	451	43	452	44
rect	451	52	452	53
rect	451	55	452	56
rect	451	64	452	65
rect	451	67	452	68
rect	451	70	452	71
rect	451	73	452	74
rect	451	76	452	77
rect	451	79	452	80
rect	451	82	452	83
rect	451	85	452	86
rect	451	88	452	89
rect	451	91	452	92
rect	451	94	452	95
rect	451	97	452	98
rect	451	106	452	107
rect	451	109	452	110
rect	451	112	452	113
rect	451	121	452	122
rect	451	124	452	125
rect	451	127	452	128
rect	451	130	452	131
rect	451	133	452	134
rect	451	142	452	143
rect	451	145	452	146
rect	451	154	452	155
rect	451	157	452	158
rect	451	160	452	161
rect	451	163	452	164
rect	451	172	452	173
rect	451	175	452	176
rect	451	178	452	179
rect	451	181	452	182
rect	451	190	452	191
rect	451	196	452	197
rect	451	211	452	212
rect	451	214	452	215
rect	451	217	452	218
rect	451	220	452	221
rect	451	229	452	230
rect	451	232	452	233
rect	451	235	452	236
rect	451	238	452	239
rect	451	244	452	245
rect	451	247	452	248
rect	451	250	452	251
rect	451	253	452	254
rect	451	256	452	257
rect	451	259	452	260
rect	451	268	452	269
rect	451	277	452	278
rect	451	286	452	287
rect	451	289	452	290
rect	451	295	452	296
rect	451	298	452	299
rect	451	301	452	302
rect	451	304	452	305
rect	451	310	452	311
rect	451	313	452	314
rect	451	316	452	317
rect	451	331	452	332
rect	451	334	452	335
rect	451	346	452	347
rect	458	4	459	5
rect	458	7	459	8
rect	458	10	459	11
rect	458	16	459	17
rect	458	19	459	20
rect	458	22	459	23
rect	458	25	459	26
rect	458	28	459	29
rect	458	37	459	38
rect	458	40	459	41
rect	458	43	459	44
rect	458	52	459	53
rect	458	55	459	56
rect	458	64	459	65
rect	458	67	459	68
rect	458	70	459	71
rect	458	73	459	74
rect	458	76	459	77
rect	458	79	459	80
rect	458	82	459	83
rect	458	85	459	86
rect	458	88	459	89
rect	458	91	459	92
rect	458	94	459	95
rect	458	97	459	98
rect	458	100	459	101
rect	458	106	459	107
rect	458	109	459	110
rect	458	112	459	113
rect	458	115	459	116
rect	458	121	459	122
rect	458	124	459	125
rect	458	127	459	128
rect	458	130	459	131
rect	458	133	459	134
rect	458	142	459	143
rect	458	145	459	146
rect	458	151	459	152
rect	458	154	459	155
rect	458	157	459	158
rect	458	160	459	161
rect	458	163	459	164
rect	458	169	459	170
rect	458	172	459	173
rect	458	175	459	176
rect	458	178	459	179
rect	458	181	459	182
rect	458	193	459	194
rect	458	196	459	197
rect	458	211	459	212
rect	458	214	459	215
rect	458	217	459	218
rect	458	220	459	221
rect	458	223	459	224
rect	458	229	459	230
rect	458	232	459	233
rect	458	235	459	236
rect	458	238	459	239
rect	458	247	459	248
rect	458	250	459	251
rect	458	253	459	254
rect	458	256	459	257
rect	458	259	459	260
rect	458	268	459	269
rect	458	277	459	278
rect	458	280	459	281
rect	458	286	459	287
rect	458	295	459	296
rect	458	298	459	299
rect	458	301	459	302
rect	458	307	459	308
rect	458	310	459	311
rect	458	313	459	314
rect	458	316	459	317
rect	458	331	459	332
rect	458	343	459	344
rect	458	346	459	347
rect	459	4	460	5
rect	459	7	460	8
rect	459	10	460	11
rect	459	16	460	17
rect	459	19	460	20
rect	459	22	460	23
rect	459	25	460	26
rect	459	28	460	29
rect	459	37	460	38
rect	459	40	460	41
rect	459	43	460	44
rect	459	52	460	53
rect	459	55	460	56
rect	459	64	460	65
rect	459	67	460	68
rect	459	70	460	71
rect	459	73	460	74
rect	459	76	460	77
rect	459	79	460	80
rect	459	82	460	83
rect	459	85	460	86
rect	459	88	460	89
rect	459	91	460	92
rect	459	94	460	95
rect	459	97	460	98
rect	459	100	460	101
rect	459	106	460	107
rect	459	109	460	110
rect	459	112	460	113
rect	459	115	460	116
rect	459	121	460	122
rect	459	124	460	125
rect	459	127	460	128
rect	459	130	460	131
rect	459	133	460	134
rect	459	142	460	143
rect	459	145	460	146
rect	459	151	460	152
rect	459	154	460	155
rect	459	157	460	158
rect	459	160	460	161
rect	459	163	460	164
rect	459	169	460	170
rect	459	172	460	173
rect	459	175	460	176
rect	459	178	460	179
rect	459	181	460	182
rect	459	193	460	194
rect	459	196	460	197
rect	459	211	460	212
rect	459	214	460	215
rect	459	217	460	218
rect	459	220	460	221
rect	459	223	460	224
rect	459	229	460	230
rect	459	232	460	233
rect	459	235	460	236
rect	459	238	460	239
rect	459	247	460	248
rect	459	250	460	251
rect	459	253	460	254
rect	459	256	460	257
rect	459	259	460	260
rect	459	268	460	269
rect	459	277	460	278
rect	459	280	460	281
rect	459	295	460	296
rect	459	298	460	299
rect	459	301	460	302
rect	459	307	460	308
rect	459	310	460	311
rect	459	313	460	314
rect	459	316	460	317
rect	459	331	460	332
rect	459	343	460	344
rect	459	346	460	347
rect	460	4	461	5
rect	460	7	461	8
rect	460	10	461	11
rect	460	16	461	17
rect	460	19	461	20
rect	460	22	461	23
rect	460	25	461	26
rect	460	28	461	29
rect	460	37	461	38
rect	460	40	461	41
rect	460	43	461	44
rect	460	52	461	53
rect	460	55	461	56
rect	460	64	461	65
rect	460	67	461	68
rect	460	70	461	71
rect	460	73	461	74
rect	460	76	461	77
rect	460	79	461	80
rect	460	82	461	83
rect	460	85	461	86
rect	460	88	461	89
rect	460	91	461	92
rect	460	94	461	95
rect	460	97	461	98
rect	460	100	461	101
rect	460	106	461	107
rect	460	109	461	110
rect	460	112	461	113
rect	460	115	461	116
rect	460	121	461	122
rect	460	124	461	125
rect	460	127	461	128
rect	460	130	461	131
rect	460	133	461	134
rect	460	142	461	143
rect	460	145	461	146
rect	460	151	461	152
rect	460	154	461	155
rect	460	157	461	158
rect	460	160	461	161
rect	460	163	461	164
rect	460	169	461	170
rect	460	172	461	173
rect	460	175	461	176
rect	460	178	461	179
rect	460	181	461	182
rect	460	193	461	194
rect	460	196	461	197
rect	460	211	461	212
rect	460	214	461	215
rect	460	217	461	218
rect	460	220	461	221
rect	460	223	461	224
rect	460	229	461	230
rect	460	232	461	233
rect	460	235	461	236
rect	460	238	461	239
rect	460	247	461	248
rect	460	250	461	251
rect	460	253	461	254
rect	460	256	461	257
rect	460	259	461	260
rect	460	268	461	269
rect	460	274	461	275
rect	460	277	461	278
rect	460	280	461	281
rect	460	295	461	296
rect	460	298	461	299
rect	460	301	461	302
rect	460	307	461	308
rect	460	310	461	311
rect	460	313	461	314
rect	460	316	461	317
rect	460	331	461	332
rect	460	343	461	344
rect	460	346	461	347
rect	461	4	462	5
rect	461	7	462	8
rect	461	10	462	11
rect	461	16	462	17
rect	461	19	462	20
rect	461	22	462	23
rect	461	25	462	26
rect	461	28	462	29
rect	461	37	462	38
rect	461	40	462	41
rect	461	43	462	44
rect	461	52	462	53
rect	461	55	462	56
rect	461	64	462	65
rect	461	67	462	68
rect	461	70	462	71
rect	461	73	462	74
rect	461	76	462	77
rect	461	79	462	80
rect	461	82	462	83
rect	461	85	462	86
rect	461	88	462	89
rect	461	91	462	92
rect	461	94	462	95
rect	461	97	462	98
rect	461	100	462	101
rect	461	106	462	107
rect	461	109	462	110
rect	461	112	462	113
rect	461	115	462	116
rect	461	121	462	122
rect	461	124	462	125
rect	461	127	462	128
rect	461	130	462	131
rect	461	133	462	134
rect	461	142	462	143
rect	461	145	462	146
rect	461	151	462	152
rect	461	154	462	155
rect	461	157	462	158
rect	461	160	462	161
rect	461	163	462	164
rect	461	169	462	170
rect	461	172	462	173
rect	461	175	462	176
rect	461	178	462	179
rect	461	181	462	182
rect	461	193	462	194
rect	461	196	462	197
rect	461	211	462	212
rect	461	214	462	215
rect	461	217	462	218
rect	461	220	462	221
rect	461	223	462	224
rect	461	229	462	230
rect	461	232	462	233
rect	461	235	462	236
rect	461	238	462	239
rect	461	247	462	248
rect	461	250	462	251
rect	461	253	462	254
rect	461	256	462	257
rect	461	259	462	260
rect	461	268	462	269
rect	461	274	462	275
rect	461	277	462	278
rect	461	280	462	281
rect	461	295	462	296
rect	461	298	462	299
rect	461	301	462	302
rect	461	307	462	308
rect	461	313	462	314
rect	461	316	462	317
rect	461	331	462	332
rect	461	343	462	344
rect	461	346	462	347
rect	462	4	463	5
rect	462	7	463	8
rect	462	10	463	11
rect	462	16	463	17
rect	462	19	463	20
rect	462	22	463	23
rect	462	25	463	26
rect	462	28	463	29
rect	462	37	463	38
rect	462	40	463	41
rect	462	43	463	44
rect	462	52	463	53
rect	462	55	463	56
rect	462	64	463	65
rect	462	67	463	68
rect	462	70	463	71
rect	462	73	463	74
rect	462	76	463	77
rect	462	79	463	80
rect	462	82	463	83
rect	462	85	463	86
rect	462	88	463	89
rect	462	91	463	92
rect	462	94	463	95
rect	462	97	463	98
rect	462	100	463	101
rect	462	106	463	107
rect	462	109	463	110
rect	462	112	463	113
rect	462	115	463	116
rect	462	121	463	122
rect	462	124	463	125
rect	462	127	463	128
rect	462	130	463	131
rect	462	133	463	134
rect	462	142	463	143
rect	462	145	463	146
rect	462	151	463	152
rect	462	154	463	155
rect	462	157	463	158
rect	462	160	463	161
rect	462	163	463	164
rect	462	169	463	170
rect	462	172	463	173
rect	462	175	463	176
rect	462	178	463	179
rect	462	181	463	182
rect	462	193	463	194
rect	462	196	463	197
rect	462	211	463	212
rect	462	214	463	215
rect	462	217	463	218
rect	462	220	463	221
rect	462	223	463	224
rect	462	229	463	230
rect	462	232	463	233
rect	462	235	463	236
rect	462	238	463	239
rect	462	247	463	248
rect	462	250	463	251
rect	462	253	463	254
rect	462	256	463	257
rect	462	259	463	260
rect	462	268	463	269
rect	462	274	463	275
rect	462	277	463	278
rect	462	280	463	281
rect	462	286	463	287
rect	462	295	463	296
rect	462	298	463	299
rect	462	301	463	302
rect	462	307	463	308
rect	462	313	463	314
rect	462	316	463	317
rect	462	331	463	332
rect	462	343	463	344
rect	462	346	463	347
rect	463	4	464	5
rect	463	7	464	8
rect	463	10	464	11
rect	463	16	464	17
rect	463	19	464	20
rect	463	22	464	23
rect	463	25	464	26
rect	463	28	464	29
rect	463	37	464	38
rect	463	40	464	41
rect	463	43	464	44
rect	463	52	464	53
rect	463	55	464	56
rect	463	64	464	65
rect	463	67	464	68
rect	463	70	464	71
rect	463	73	464	74
rect	463	76	464	77
rect	463	79	464	80
rect	463	82	464	83
rect	463	85	464	86
rect	463	88	464	89
rect	463	91	464	92
rect	463	94	464	95
rect	463	97	464	98
rect	463	100	464	101
rect	463	106	464	107
rect	463	109	464	110
rect	463	112	464	113
rect	463	115	464	116
rect	463	121	464	122
rect	463	127	464	128
rect	463	130	464	131
rect	463	133	464	134
rect	463	142	464	143
rect	463	145	464	146
rect	463	151	464	152
rect	463	154	464	155
rect	463	157	464	158
rect	463	160	464	161
rect	463	163	464	164
rect	463	169	464	170
rect	463	172	464	173
rect	463	175	464	176
rect	463	178	464	179
rect	463	181	464	182
rect	463	193	464	194
rect	463	196	464	197
rect	463	211	464	212
rect	463	214	464	215
rect	463	217	464	218
rect	463	220	464	221
rect	463	223	464	224
rect	463	229	464	230
rect	463	232	464	233
rect	463	235	464	236
rect	463	238	464	239
rect	463	247	464	248
rect	463	250	464	251
rect	463	253	464	254
rect	463	256	464	257
rect	463	259	464	260
rect	463	268	464	269
rect	463	274	464	275
rect	463	277	464	278
rect	463	280	464	281
rect	463	286	464	287
rect	463	295	464	296
rect	463	298	464	299
rect	463	301	464	302
rect	463	307	464	308
rect	463	313	464	314
rect	463	316	464	317
rect	463	331	464	332
rect	463	343	464	344
rect	463	346	464	347
rect	464	4	465	5
rect	464	7	465	8
rect	464	10	465	11
rect	464	16	465	17
rect	464	19	465	20
rect	464	22	465	23
rect	464	25	465	26
rect	464	28	465	29
rect	464	37	465	38
rect	464	40	465	41
rect	464	43	465	44
rect	464	52	465	53
rect	464	55	465	56
rect	464	64	465	65
rect	464	67	465	68
rect	464	70	465	71
rect	464	73	465	74
rect	464	76	465	77
rect	464	79	465	80
rect	464	82	465	83
rect	464	85	465	86
rect	464	88	465	89
rect	464	91	465	92
rect	464	94	465	95
rect	464	97	465	98
rect	464	100	465	101
rect	464	106	465	107
rect	464	109	465	110
rect	464	112	465	113
rect	464	115	465	116
rect	464	121	465	122
rect	464	127	465	128
rect	464	130	465	131
rect	464	133	465	134
rect	464	142	465	143
rect	464	145	465	146
rect	464	151	465	152
rect	464	154	465	155
rect	464	157	465	158
rect	464	160	465	161
rect	464	163	465	164
rect	464	169	465	170
rect	464	172	465	173
rect	464	175	465	176
rect	464	178	465	179
rect	464	181	465	182
rect	464	193	465	194
rect	464	196	465	197
rect	464	211	465	212
rect	464	214	465	215
rect	464	217	465	218
rect	464	220	465	221
rect	464	223	465	224
rect	464	229	465	230
rect	464	232	465	233
rect	464	235	465	236
rect	464	238	465	239
rect	464	247	465	248
rect	464	250	465	251
rect	464	253	465	254
rect	464	256	465	257
rect	464	259	465	260
rect	464	268	465	269
rect	464	274	465	275
rect	464	277	465	278
rect	464	280	465	281
rect	464	286	465	287
rect	464	295	465	296
rect	464	298	465	299
rect	464	301	465	302
rect	464	307	465	308
rect	464	310	465	311
rect	464	313	465	314
rect	464	316	465	317
rect	464	331	465	332
rect	464	343	465	344
rect	464	346	465	347
rect	465	4	466	5
rect	465	7	466	8
rect	465	10	466	11
rect	465	16	466	17
rect	465	19	466	20
rect	465	22	466	23
rect	465	25	466	26
rect	465	28	466	29
rect	465	37	466	38
rect	465	40	466	41
rect	465	43	466	44
rect	465	52	466	53
rect	465	55	466	56
rect	465	64	466	65
rect	465	67	466	68
rect	465	70	466	71
rect	465	73	466	74
rect	465	76	466	77
rect	465	79	466	80
rect	465	82	466	83
rect	465	85	466	86
rect	465	88	466	89
rect	465	91	466	92
rect	465	94	466	95
rect	465	97	466	98
rect	465	100	466	101
rect	465	106	466	107
rect	465	109	466	110
rect	465	112	466	113
rect	465	115	466	116
rect	465	121	466	122
rect	465	127	466	128
rect	465	130	466	131
rect	465	142	466	143
rect	465	145	466	146
rect	465	151	466	152
rect	465	154	466	155
rect	465	157	466	158
rect	465	160	466	161
rect	465	163	466	164
rect	465	169	466	170
rect	465	172	466	173
rect	465	175	466	176
rect	465	178	466	179
rect	465	181	466	182
rect	465	193	466	194
rect	465	211	466	212
rect	465	214	466	215
rect	465	217	466	218
rect	465	220	466	221
rect	465	223	466	224
rect	465	229	466	230
rect	465	232	466	233
rect	465	235	466	236
rect	465	247	466	248
rect	465	250	466	251
rect	465	253	466	254
rect	465	256	466	257
rect	465	259	466	260
rect	465	268	466	269
rect	465	274	466	275
rect	465	277	466	278
rect	465	280	466	281
rect	465	286	466	287
rect	465	295	466	296
rect	465	298	466	299
rect	465	301	466	302
rect	465	307	466	308
rect	465	310	466	311
rect	465	313	466	314
rect	465	316	466	317
rect	465	331	466	332
rect	465	343	466	344
rect	465	346	466	347
rect	466	4	467	5
rect	466	7	467	8
rect	466	10	467	11
rect	466	16	467	17
rect	466	19	467	20
rect	466	22	467	23
rect	466	25	467	26
rect	466	28	467	29
rect	466	37	467	38
rect	466	40	467	41
rect	466	43	467	44
rect	466	52	467	53
rect	466	55	467	56
rect	466	64	467	65
rect	466	67	467	68
rect	466	70	467	71
rect	466	73	467	74
rect	466	76	467	77
rect	466	79	467	80
rect	466	82	467	83
rect	466	85	467	86
rect	466	88	467	89
rect	466	91	467	92
rect	466	94	467	95
rect	466	97	467	98
rect	466	100	467	101
rect	466	106	467	107
rect	466	109	467	110
rect	466	112	467	113
rect	466	115	467	116
rect	466	121	467	122
rect	466	124	467	125
rect	466	127	467	128
rect	466	130	467	131
rect	466	142	467	143
rect	466	145	467	146
rect	466	151	467	152
rect	466	154	467	155
rect	466	157	467	158
rect	466	160	467	161
rect	466	163	467	164
rect	466	169	467	170
rect	466	172	467	173
rect	466	175	467	176
rect	466	178	467	179
rect	466	181	467	182
rect	466	187	467	188
rect	466	193	467	194
rect	466	211	467	212
rect	466	214	467	215
rect	466	217	467	218
rect	466	220	467	221
rect	466	223	467	224
rect	466	226	467	227
rect	466	229	467	230
rect	466	232	467	233
rect	466	235	467	236
rect	466	247	467	248
rect	466	250	467	251
rect	466	253	467	254
rect	466	256	467	257
rect	466	259	467	260
rect	466	268	467	269
rect	466	274	467	275
rect	466	277	467	278
rect	466	280	467	281
rect	466	286	467	287
rect	466	295	467	296
rect	466	298	467	299
rect	466	301	467	302
rect	466	307	467	308
rect	466	310	467	311
rect	466	313	467	314
rect	466	316	467	317
rect	466	331	467	332
rect	466	343	467	344
rect	466	346	467	347
rect	467	4	468	5
rect	467	7	468	8
rect	467	10	468	11
rect	467	16	468	17
rect	467	19	468	20
rect	467	22	468	23
rect	467	25	468	26
rect	467	28	468	29
rect	467	37	468	38
rect	467	40	468	41
rect	467	43	468	44
rect	467	52	468	53
rect	467	55	468	56
rect	467	64	468	65
rect	467	67	468	68
rect	467	70	468	71
rect	467	73	468	74
rect	467	76	468	77
rect	467	79	468	80
rect	467	82	468	83
rect	467	85	468	86
rect	467	88	468	89
rect	467	91	468	92
rect	467	94	468	95
rect	467	97	468	98
rect	467	100	468	101
rect	467	106	468	107
rect	467	109	468	110
rect	467	112	468	113
rect	467	115	468	116
rect	467	121	468	122
rect	467	124	468	125
rect	467	127	468	128
rect	467	130	468	131
rect	467	142	468	143
rect	467	145	468	146
rect	467	151	468	152
rect	467	154	468	155
rect	467	157	468	158
rect	467	160	468	161
rect	467	163	468	164
rect	467	169	468	170
rect	467	175	468	176
rect	467	178	468	179
rect	467	181	468	182
rect	467	187	468	188
rect	467	193	468	194
rect	467	214	468	215
rect	467	217	468	218
rect	467	220	468	221
rect	467	223	468	224
rect	467	226	468	227
rect	467	229	468	230
rect	467	232	468	233
rect	467	235	468	236
rect	467	247	468	248
rect	467	250	468	251
rect	467	253	468	254
rect	467	256	468	257
rect	467	268	468	269
rect	467	274	468	275
rect	467	277	468	278
rect	467	280	468	281
rect	467	286	468	287
rect	467	295	468	296
rect	467	298	468	299
rect	467	301	468	302
rect	467	307	468	308
rect	467	310	468	311
rect	467	313	468	314
rect	467	316	468	317
rect	467	331	468	332
rect	467	343	468	344
rect	467	346	468	347
rect	468	4	469	5
rect	468	7	469	8
rect	468	10	469	11
rect	468	16	469	17
rect	468	19	469	20
rect	468	22	469	23
rect	468	25	469	26
rect	468	28	469	29
rect	468	37	469	38
rect	468	40	469	41
rect	468	43	469	44
rect	468	52	469	53
rect	468	55	469	56
rect	468	64	469	65
rect	468	67	469	68
rect	468	70	469	71
rect	468	73	469	74
rect	468	76	469	77
rect	468	79	469	80
rect	468	82	469	83
rect	468	85	469	86
rect	468	88	469	89
rect	468	91	469	92
rect	468	94	469	95
rect	468	97	469	98
rect	468	100	469	101
rect	468	106	469	107
rect	468	109	469	110
rect	468	112	469	113
rect	468	115	469	116
rect	468	121	469	122
rect	468	124	469	125
rect	468	127	469	128
rect	468	130	469	131
rect	468	133	469	134
rect	468	142	469	143
rect	468	145	469	146
rect	468	151	469	152
rect	468	154	469	155
rect	468	157	469	158
rect	468	160	469	161
rect	468	163	469	164
rect	468	169	469	170
rect	468	175	469	176
rect	468	178	469	179
rect	468	181	469	182
rect	468	187	469	188
rect	468	193	469	194
rect	468	196	469	197
rect	468	214	469	215
rect	468	217	469	218
rect	468	220	469	221
rect	468	223	469	224
rect	468	226	469	227
rect	468	229	469	230
rect	468	232	469	233
rect	468	235	469	236
rect	468	238	469	239
rect	468	247	469	248
rect	468	250	469	251
rect	468	253	469	254
rect	468	256	469	257
rect	468	268	469	269
rect	468	274	469	275
rect	468	277	469	278
rect	468	280	469	281
rect	468	286	469	287
rect	468	295	469	296
rect	468	298	469	299
rect	468	301	469	302
rect	468	307	469	308
rect	468	310	469	311
rect	468	313	469	314
rect	468	316	469	317
rect	468	331	469	332
rect	468	343	469	344
rect	468	346	469	347
rect	469	4	470	5
rect	469	7	470	8
rect	469	10	470	11
rect	469	16	470	17
rect	469	19	470	20
rect	469	22	470	23
rect	469	25	470	26
rect	469	28	470	29
rect	469	37	470	38
rect	469	40	470	41
rect	469	43	470	44
rect	469	52	470	53
rect	469	55	470	56
rect	469	67	470	68
rect	469	70	470	71
rect	469	73	470	74
rect	469	76	470	77
rect	469	79	470	80
rect	469	82	470	83
rect	469	85	470	86
rect	469	88	470	89
rect	469	91	470	92
rect	469	94	470	95
rect	469	97	470	98
rect	469	100	470	101
rect	469	106	470	107
rect	469	109	470	110
rect	469	112	470	113
rect	469	115	470	116
rect	469	121	470	122
rect	469	124	470	125
rect	469	127	470	128
rect	469	130	470	131
rect	469	133	470	134
rect	469	142	470	143
rect	469	145	470	146
rect	469	151	470	152
rect	469	154	470	155
rect	469	157	470	158
rect	469	160	470	161
rect	469	169	470	170
rect	469	175	470	176
rect	469	178	470	179
rect	469	181	470	182
rect	469	187	470	188
rect	469	193	470	194
rect	469	196	470	197
rect	469	214	470	215
rect	469	220	470	221
rect	469	226	470	227
rect	469	229	470	230
rect	469	232	470	233
rect	469	235	470	236
rect	469	238	470	239
rect	469	247	470	248
rect	469	250	470	251
rect	469	253	470	254
rect	469	256	470	257
rect	469	268	470	269
rect	469	274	470	275
rect	469	277	470	278
rect	469	280	470	281
rect	469	286	470	287
rect	469	295	470	296
rect	469	298	470	299
rect	469	301	470	302
rect	469	307	470	308
rect	469	310	470	311
rect	469	313	470	314
rect	469	316	470	317
rect	469	331	470	332
rect	469	343	470	344
rect	470	4	471	5
rect	470	7	471	8
rect	470	10	471	11
rect	470	16	471	17
rect	470	19	471	20
rect	470	22	471	23
rect	470	25	471	26
rect	470	28	471	29
rect	470	37	471	38
rect	470	40	471	41
rect	470	43	471	44
rect	470	46	471	47
rect	470	52	471	53
rect	470	55	471	56
rect	470	67	471	68
rect	470	70	471	71
rect	470	73	471	74
rect	470	76	471	77
rect	470	79	471	80
rect	470	82	471	83
rect	470	85	471	86
rect	470	88	471	89
rect	470	91	471	92
rect	470	94	471	95
rect	470	97	471	98
rect	470	100	471	101
rect	470	106	471	107
rect	470	109	471	110
rect	470	112	471	113
rect	470	115	471	116
rect	470	121	471	122
rect	470	124	471	125
rect	470	127	471	128
rect	470	130	471	131
rect	470	133	471	134
rect	470	142	471	143
rect	470	145	471	146
rect	470	151	471	152
rect	470	154	471	155
rect	470	157	471	158
rect	470	160	471	161
rect	470	169	471	170
rect	470	172	471	173
rect	470	175	471	176
rect	470	178	471	179
rect	470	181	471	182
rect	470	187	471	188
rect	470	193	471	194
rect	470	196	471	197
rect	470	211	471	212
rect	470	214	471	215
rect	470	220	471	221
rect	470	226	471	227
rect	470	229	471	230
rect	470	232	471	233
rect	470	235	471	236
rect	470	238	471	239
rect	470	247	471	248
rect	470	250	471	251
rect	470	253	471	254
rect	470	256	471	257
rect	470	268	471	269
rect	470	274	471	275
rect	470	277	471	278
rect	470	280	471	281
rect	470	286	471	287
rect	470	295	471	296
rect	470	298	471	299
rect	470	301	471	302
rect	470	307	471	308
rect	470	310	471	311
rect	470	313	471	314
rect	470	316	471	317
rect	470	331	471	332
rect	470	343	471	344
rect	471	4	472	5
rect	471	7	472	8
rect	471	10	472	11
rect	471	16	472	17
rect	471	19	472	20
rect	471	22	472	23
rect	471	25	472	26
rect	471	28	472	29
rect	471	37	472	38
rect	471	40	472	41
rect	471	43	472	44
rect	471	46	472	47
rect	471	52	472	53
rect	471	55	472	56
rect	471	67	472	68
rect	471	70	472	71
rect	471	73	472	74
rect	471	76	472	77
rect	471	82	472	83
rect	471	85	472	86
rect	471	88	472	89
rect	471	91	472	92
rect	471	94	472	95
rect	471	97	472	98
rect	471	100	472	101
rect	471	106	472	107
rect	471	109	472	110
rect	471	112	472	113
rect	471	115	472	116
rect	471	121	472	122
rect	471	124	472	125
rect	471	127	472	128
rect	471	130	472	131
rect	471	133	472	134
rect	471	142	472	143
rect	471	145	472	146
rect	471	157	472	158
rect	471	160	472	161
rect	471	169	472	170
rect	471	172	472	173
rect	471	178	472	179
rect	471	181	472	182
rect	471	187	472	188
rect	471	193	472	194
rect	471	196	472	197
rect	471	211	472	212
rect	471	214	472	215
rect	471	220	472	221
rect	471	226	472	227
rect	471	229	472	230
rect	471	232	472	233
rect	471	235	472	236
rect	471	238	472	239
rect	471	250	472	251
rect	471	253	472	254
rect	471	256	472	257
rect	471	268	472	269
rect	471	274	472	275
rect	471	277	472	278
rect	471	280	472	281
rect	471	286	472	287
rect	471	295	472	296
rect	471	298	472	299
rect	471	301	472	302
rect	471	307	472	308
rect	471	310	472	311
rect	471	313	472	314
rect	471	316	472	317
rect	471	331	472	332
rect	471	343	472	344
rect	472	4	473	5
rect	472	7	473	8
rect	472	10	473	11
rect	472	16	473	17
rect	472	19	473	20
rect	472	22	473	23
rect	472	25	473	26
rect	472	28	473	29
rect	472	37	473	38
rect	472	40	473	41
rect	472	43	473	44
rect	472	46	473	47
rect	472	52	473	53
rect	472	55	473	56
rect	472	64	473	65
rect	472	67	473	68
rect	472	70	473	71
rect	472	73	473	74
rect	472	76	473	77
rect	472	82	473	83
rect	472	85	473	86
rect	472	88	473	89
rect	472	91	473	92
rect	472	94	473	95
rect	472	97	473	98
rect	472	100	473	101
rect	472	106	473	107
rect	472	109	473	110
rect	472	112	473	113
rect	472	115	473	116
rect	472	121	473	122
rect	472	124	473	125
rect	472	127	473	128
rect	472	130	473	131
rect	472	133	473	134
rect	472	142	473	143
rect	472	145	473	146
rect	472	157	473	158
rect	472	160	473	161
rect	472	163	473	164
rect	472	169	473	170
rect	472	172	473	173
rect	472	178	473	179
rect	472	181	473	182
rect	472	187	473	188
rect	472	193	473	194
rect	472	196	473	197
rect	472	211	473	212
rect	472	214	473	215
rect	472	217	473	218
rect	472	220	473	221
rect	472	226	473	227
rect	472	229	473	230
rect	472	232	473	233
rect	472	235	473	236
rect	472	238	473	239
rect	472	250	473	251
rect	472	253	473	254
rect	472	256	473	257
rect	472	268	473	269
rect	472	274	473	275
rect	472	277	473	278
rect	472	280	473	281
rect	472	286	473	287
rect	472	295	473	296
rect	472	298	473	299
rect	472	301	473	302
rect	472	307	473	308
rect	472	310	473	311
rect	472	313	473	314
rect	472	316	473	317
rect	472	331	473	332
rect	472	343	473	344
rect	473	4	474	5
rect	473	7	474	8
rect	473	10	474	11
rect	473	16	474	17
rect	473	19	474	20
rect	473	22	474	23
rect	473	25	474	26
rect	473	28	474	29
rect	473	37	474	38
rect	473	40	474	41
rect	473	43	474	44
rect	473	46	474	47
rect	473	52	474	53
rect	473	55	474	56
rect	473	64	474	65
rect	473	67	474	68
rect	473	70	474	71
rect	473	76	474	77
rect	473	82	474	83
rect	473	85	474	86
rect	473	88	474	89
rect	473	91	474	92
rect	473	94	474	95
rect	473	106	474	107
rect	473	109	474	110
rect	473	115	474	116
rect	473	121	474	122
rect	473	124	474	125
rect	473	127	474	128
rect	473	130	474	131
rect	473	133	474	134
rect	473	145	474	146
rect	473	157	474	158
rect	473	160	474	161
rect	473	163	474	164
rect	473	172	474	173
rect	473	178	474	179
rect	473	187	474	188
rect	473	193	474	194
rect	473	196	474	197
rect	473	211	474	212
rect	473	217	474	218
rect	473	220	474	221
rect	473	226	474	227
rect	473	229	474	230
rect	473	232	474	233
rect	473	235	474	236
rect	473	238	474	239
rect	473	250	474	251
rect	473	253	474	254
rect	473	274	474	275
rect	473	277	474	278
rect	473	280	474	281
rect	473	286	474	287
rect	473	295	474	296
rect	473	298	474	299
rect	473	307	474	308
rect	473	310	474	311
rect	473	313	474	314
rect	473	316	474	317
rect	473	331	474	332
rect	473	343	474	344
rect	474	4	475	5
rect	474	7	475	8
rect	474	10	475	11
rect	474	16	475	17
rect	474	19	475	20
rect	474	22	475	23
rect	474	25	475	26
rect	474	28	475	29
rect	474	37	475	38
rect	474	40	475	41
rect	474	43	475	44
rect	474	46	475	47
rect	474	52	475	53
rect	474	55	475	56
rect	474	58	475	59
rect	474	64	475	65
rect	474	67	475	68
rect	474	70	475	71
rect	474	76	475	77
rect	474	79	475	80
rect	474	82	475	83
rect	474	85	475	86
rect	474	88	475	89
rect	474	91	475	92
rect	474	94	475	95
rect	474	106	475	107
rect	474	109	475	110
rect	474	115	475	116
rect	474	121	475	122
rect	474	124	475	125
rect	474	127	475	128
rect	474	130	475	131
rect	474	133	475	134
rect	474	139	475	140
rect	474	145	475	146
rect	474	151	475	152
rect	474	157	475	158
rect	474	160	475	161
rect	474	163	475	164
rect	474	172	475	173
rect	474	178	475	179
rect	474	184	475	185
rect	474	187	475	188
rect	474	193	475	194
rect	474	196	475	197
rect	474	211	475	212
rect	474	217	475	218
rect	474	220	475	221
rect	474	223	475	224
rect	474	226	475	227
rect	474	229	475	230
rect	474	232	475	233
rect	474	235	475	236
rect	474	238	475	239
rect	474	247	475	248
rect	474	250	475	251
rect	474	253	475	254
rect	474	259	475	260
rect	474	271	475	272
rect	474	274	475	275
rect	474	277	475	278
rect	474	280	475	281
rect	474	286	475	287
rect	474	295	475	296
rect	474	298	475	299
rect	474	307	475	308
rect	474	310	475	311
rect	474	313	475	314
rect	474	316	475	317
rect	474	331	475	332
rect	474	343	475	344
rect	475	4	476	5
rect	475	7	476	8
rect	475	10	476	11
rect	475	16	476	17
rect	475	19	476	20
rect	475	22	476	23
rect	475	25	476	26
rect	475	28	476	29
rect	475	37	476	38
rect	475	40	476	41
rect	475	43	476	44
rect	475	46	476	47
rect	475	52	476	53
rect	475	58	476	59
rect	475	64	476	65
rect	475	67	476	68
rect	475	70	476	71
rect	475	79	476	80
rect	475	82	476	83
rect	475	85	476	86
rect	475	88	476	89
rect	475	91	476	92
rect	475	94	476	95
rect	475	106	476	107
rect	475	109	476	110
rect	475	124	476	125
rect	475	127	476	128
rect	475	130	476	131
rect	475	133	476	134
rect	475	139	476	140
rect	475	145	476	146
rect	475	151	476	152
rect	475	160	476	161
rect	475	163	476	164
rect	475	172	476	173
rect	475	178	476	179
rect	475	184	476	185
rect	475	187	476	188
rect	475	193	476	194
rect	475	196	476	197
rect	475	211	476	212
rect	475	217	476	218
rect	475	223	476	224
rect	475	226	476	227
rect	475	229	476	230
rect	475	232	476	233
rect	475	235	476	236
rect	475	238	476	239
rect	475	247	476	248
rect	475	250	476	251
rect	475	253	476	254
rect	475	259	476	260
rect	475	271	476	272
rect	475	274	476	275
rect	475	277	476	278
rect	475	280	476	281
rect	475	286	476	287
rect	475	298	476	299
rect	475	307	476	308
rect	475	310	476	311
rect	475	313	476	314
rect	475	316	476	317
rect	475	331	476	332
rect	475	343	476	344
rect	476	4	477	5
rect	476	7	477	8
rect	476	10	477	11
rect	476	16	477	17
rect	476	19	477	20
rect	476	22	477	23
rect	476	25	477	26
rect	476	28	477	29
rect	476	37	477	38
rect	476	40	477	41
rect	476	43	477	44
rect	476	46	477	47
rect	476	52	477	53
rect	476	58	477	59
rect	476	64	477	65
rect	476	67	477	68
rect	476	70	477	71
rect	476	73	477	74
rect	476	79	477	80
rect	476	82	477	83
rect	476	85	477	86
rect	476	88	477	89
rect	476	91	477	92
rect	476	94	477	95
rect	476	100	477	101
rect	476	106	477	107
rect	476	109	477	110
rect	476	124	477	125
rect	476	127	477	128
rect	476	130	477	131
rect	476	133	477	134
rect	476	136	477	137
rect	476	139	477	140
rect	476	145	477	146
rect	476	151	477	152
rect	476	160	477	161
rect	476	163	477	164
rect	476	172	477	173
rect	476	175	477	176
rect	476	178	477	179
rect	476	181	477	182
rect	476	184	477	185
rect	476	187	477	188
rect	476	193	477	194
rect	476	196	477	197
rect	476	211	477	212
rect	476	214	477	215
rect	476	217	477	218
rect	476	223	477	224
rect	476	226	477	227
rect	476	229	477	230
rect	476	232	477	233
rect	476	235	477	236
rect	476	238	477	239
rect	476	247	477	248
rect	476	250	477	251
rect	476	253	477	254
rect	476	256	477	257
rect	476	259	477	260
rect	476	265	477	266
rect	476	268	477	269
rect	476	271	477	272
rect	476	274	477	275
rect	476	277	477	278
rect	476	280	477	281
rect	476	286	477	287
rect	476	298	477	299
rect	476	307	477	308
rect	476	310	477	311
rect	476	313	477	314
rect	476	316	477	317
rect	476	331	477	332
rect	476	343	477	344
rect	477	4	478	5
rect	477	7	478	8
rect	477	10	478	11
rect	477	16	478	17
rect	477	19	478	20
rect	477	22	478	23
rect	477	25	478	26
rect	477	28	478	29
rect	477	37	478	38
rect	477	40	478	41
rect	477	43	478	44
rect	477	46	478	47
rect	477	52	478	53
rect	477	58	478	59
rect	477	64	478	65
rect	477	67	478	68
rect	477	73	478	74
rect	477	79	478	80
rect	477	82	478	83
rect	477	85	478	86
rect	477	88	478	89
rect	477	91	478	92
rect	477	100	478	101
rect	477	106	478	107
rect	477	109	478	110
rect	477	124	478	125
rect	477	133	478	134
rect	477	136	478	137
rect	477	139	478	140
rect	477	145	478	146
rect	477	151	478	152
rect	477	160	478	161
rect	477	163	478	164
rect	477	172	478	173
rect	477	175	478	176
rect	477	181	478	182
rect	477	184	478	185
rect	477	187	478	188
rect	477	193	478	194
rect	477	196	478	197
rect	477	211	478	212
rect	477	214	478	215
rect	477	217	478	218
rect	477	223	478	224
rect	477	226	478	227
rect	477	229	478	230
rect	477	232	478	233
rect	477	238	478	239
rect	477	247	478	248
rect	477	250	478	251
rect	477	253	478	254
rect	477	256	478	257
rect	477	259	478	260
rect	477	265	478	266
rect	477	268	478	269
rect	477	271	478	272
rect	477	274	478	275
rect	477	280	478	281
rect	477	286	478	287
rect	477	298	478	299
rect	477	307	478	308
rect	477	310	478	311
rect	477	313	478	314
rect	477	331	478	332
rect	477	343	478	344
rect	478	4	479	5
rect	478	7	479	8
rect	478	10	479	11
rect	478	16	479	17
rect	478	19	479	20
rect	478	22	479	23
rect	478	25	479	26
rect	478	28	479	29
rect	478	37	479	38
rect	478	40	479	41
rect	478	43	479	44
rect	478	46	479	47
rect	478	52	479	53
rect	478	55	479	56
rect	478	58	479	59
rect	478	64	479	65
rect	478	67	479	68
rect	478	73	479	74
rect	478	76	479	77
rect	478	79	479	80
rect	478	82	479	83
rect	478	85	479	86
rect	478	88	479	89
rect	478	91	479	92
rect	478	100	479	101
rect	478	106	479	107
rect	478	109	479	110
rect	478	121	479	122
rect	478	124	479	125
rect	478	133	479	134
rect	478	136	479	137
rect	478	139	479	140
rect	478	142	479	143
rect	478	145	479	146
rect	478	151	479	152
rect	478	160	479	161
rect	478	163	479	164
rect	478	169	479	170
rect	478	172	479	173
rect	478	175	479	176
rect	478	181	479	182
rect	478	184	479	185
rect	478	187	479	188
rect	478	193	479	194
rect	478	196	479	197
rect	478	208	479	209
rect	478	211	479	212
rect	478	214	479	215
rect	478	217	479	218
rect	478	223	479	224
rect	478	226	479	227
rect	478	229	479	230
rect	478	232	479	233
rect	478	238	479	239
rect	478	244	479	245
rect	478	247	479	248
rect	478	250	479	251
rect	478	253	479	254
rect	478	256	479	257
rect	478	259	479	260
rect	478	265	479	266
rect	478	268	479	269
rect	478	271	479	272
rect	478	274	479	275
rect	478	280	479	281
rect	478	286	479	287
rect	478	292	479	293
rect	478	298	479	299
rect	478	307	479	308
rect	478	310	479	311
rect	478	313	479	314
rect	478	331	479	332
rect	478	343	479	344
rect	479	4	480	5
rect	479	7	480	8
rect	479	10	480	11
rect	479	16	480	17
rect	479	19	480	20
rect	479	22	480	23
rect	479	25	480	26
rect	479	28	480	29
rect	479	40	480	41
rect	479	43	480	44
rect	479	46	480	47
rect	479	52	480	53
rect	479	55	480	56
rect	479	58	480	59
rect	479	64	480	65
rect	479	67	480	68
rect	479	73	480	74
rect	479	76	480	77
rect	479	79	480	80
rect	479	82	480	83
rect	479	85	480	86
rect	479	88	480	89
rect	479	91	480	92
rect	479	100	480	101
rect	479	106	480	107
rect	479	109	480	110
rect	479	121	480	122
rect	479	124	480	125
rect	479	133	480	134
rect	479	136	480	137
rect	479	139	480	140
rect	479	142	480	143
rect	479	145	480	146
rect	479	151	480	152
rect	479	160	480	161
rect	479	163	480	164
rect	479	169	480	170
rect	479	172	480	173
rect	479	175	480	176
rect	479	181	480	182
rect	479	184	480	185
rect	479	187	480	188
rect	479	193	480	194
rect	479	196	480	197
rect	479	208	480	209
rect	479	211	480	212
rect	479	214	480	215
rect	479	217	480	218
rect	479	223	480	224
rect	479	226	480	227
rect	479	229	480	230
rect	479	232	480	233
rect	479	238	480	239
rect	479	244	480	245
rect	479	247	480	248
rect	479	250	480	251
rect	479	253	480	254
rect	479	256	480	257
rect	479	259	480	260
rect	479	265	480	266
rect	479	268	480	269
rect	479	271	480	272
rect	479	274	480	275
rect	479	280	480	281
rect	479	286	480	287
rect	479	292	480	293
rect	479	298	480	299
rect	479	310	480	311
rect	479	313	480	314
rect	479	331	480	332
rect	479	343	480	344
rect	480	4	481	5
rect	480	7	481	8
rect	480	10	481	11
rect	480	16	481	17
rect	480	19	481	20
rect	480	22	481	23
rect	480	25	481	26
rect	480	28	481	29
rect	480	40	481	41
rect	480	43	481	44
rect	480	46	481	47
rect	480	52	481	53
rect	480	55	481	56
rect	480	58	481	59
rect	480	64	481	65
rect	480	67	481	68
rect	480	73	481	74
rect	480	76	481	77
rect	480	79	481	80
rect	480	82	481	83
rect	480	85	481	86
rect	480	88	481	89
rect	480	91	481	92
rect	480	100	481	101
rect	480	106	481	107
rect	480	109	481	110
rect	480	121	481	122
rect	480	124	481	125
rect	480	133	481	134
rect	480	136	481	137
rect	480	139	481	140
rect	480	142	481	143
rect	480	145	481	146
rect	480	151	481	152
rect	480	160	481	161
rect	480	163	481	164
rect	480	169	481	170
rect	480	172	481	173
rect	480	175	481	176
rect	480	181	481	182
rect	480	184	481	185
rect	480	187	481	188
rect	480	193	481	194
rect	480	196	481	197
rect	480	208	481	209
rect	480	211	481	212
rect	480	214	481	215
rect	480	217	481	218
rect	480	223	481	224
rect	480	226	481	227
rect	480	229	481	230
rect	480	232	481	233
rect	480	238	481	239
rect	480	244	481	245
rect	480	247	481	248
rect	480	250	481	251
rect	480	253	481	254
rect	480	256	481	257
rect	480	259	481	260
rect	480	265	481	266
rect	480	268	481	269
rect	480	271	481	272
rect	480	274	481	275
rect	480	280	481	281
rect	480	286	481	287
rect	480	292	481	293
rect	480	298	481	299
rect	480	310	481	311
rect	480	313	481	314
rect	480	331	481	332
rect	480	343	481	344
rect	481	4	482	5
rect	481	7	482	8
rect	481	10	482	11
rect	481	19	482	20
rect	481	22	482	23
rect	481	25	482	26
rect	481	28	482	29
rect	481	40	482	41
rect	481	43	482	44
rect	481	46	482	47
rect	481	52	482	53
rect	481	55	482	56
rect	481	58	482	59
rect	481	64	482	65
rect	481	67	482	68
rect	481	73	482	74
rect	481	76	482	77
rect	481	79	482	80
rect	481	82	482	83
rect	481	85	482	86
rect	481	88	482	89
rect	481	91	482	92
rect	481	100	482	101
rect	481	106	482	107
rect	481	109	482	110
rect	481	121	482	122
rect	481	124	482	125
rect	481	133	482	134
rect	481	136	482	137
rect	481	139	482	140
rect	481	142	482	143
rect	481	145	482	146
rect	481	151	482	152
rect	481	160	482	161
rect	481	163	482	164
rect	481	169	482	170
rect	481	172	482	173
rect	481	175	482	176
rect	481	181	482	182
rect	481	184	482	185
rect	481	187	482	188
rect	481	193	482	194
rect	481	196	482	197
rect	481	208	482	209
rect	481	211	482	212
rect	481	214	482	215
rect	481	217	482	218
rect	481	223	482	224
rect	481	226	482	227
rect	481	229	482	230
rect	481	232	482	233
rect	481	238	482	239
rect	481	244	482	245
rect	481	247	482	248
rect	481	250	482	251
rect	481	253	482	254
rect	481	256	482	257
rect	481	259	482	260
rect	481	265	482	266
rect	481	268	482	269
rect	481	271	482	272
rect	481	274	482	275
rect	481	280	482	281
rect	481	286	482	287
rect	481	292	482	293
rect	481	298	482	299
rect	481	310	482	311
rect	481	331	482	332
rect	481	343	482	344
rect	482	4	483	5
rect	482	7	483	8
rect	482	10	483	11
rect	482	19	483	20
rect	482	22	483	23
rect	482	25	483	26
rect	482	28	483	29
rect	482	40	483	41
rect	482	43	483	44
rect	482	46	483	47
rect	482	52	483	53
rect	482	55	483	56
rect	482	58	483	59
rect	482	64	483	65
rect	482	67	483	68
rect	482	73	483	74
rect	482	76	483	77
rect	482	79	483	80
rect	482	82	483	83
rect	482	85	483	86
rect	482	88	483	89
rect	482	91	483	92
rect	482	100	483	101
rect	482	106	483	107
rect	482	109	483	110
rect	482	121	483	122
rect	482	124	483	125
rect	482	133	483	134
rect	482	136	483	137
rect	482	139	483	140
rect	482	142	483	143
rect	482	145	483	146
rect	482	151	483	152
rect	482	160	483	161
rect	482	163	483	164
rect	482	169	483	170
rect	482	172	483	173
rect	482	175	483	176
rect	482	181	483	182
rect	482	184	483	185
rect	482	187	483	188
rect	482	193	483	194
rect	482	196	483	197
rect	482	208	483	209
rect	482	211	483	212
rect	482	214	483	215
rect	482	217	483	218
rect	482	223	483	224
rect	482	226	483	227
rect	482	229	483	230
rect	482	232	483	233
rect	482	238	483	239
rect	482	244	483	245
rect	482	247	483	248
rect	482	250	483	251
rect	482	253	483	254
rect	482	256	483	257
rect	482	259	483	260
rect	482	265	483	266
rect	482	268	483	269
rect	482	271	483	272
rect	482	274	483	275
rect	482	280	483	281
rect	482	286	483	287
rect	482	292	483	293
rect	482	298	483	299
rect	482	310	483	311
rect	482	331	483	332
rect	482	343	483	344
rect	483	4	484	5
rect	483	7	484	8
rect	483	10	484	11
rect	483	22	484	23
rect	483	25	484	26
rect	483	28	484	29
rect	483	40	484	41
rect	483	46	484	47
rect	483	52	484	53
rect	483	55	484	56
rect	483	58	484	59
rect	483	64	484	65
rect	483	73	484	74
rect	483	76	484	77
rect	483	79	484	80
rect	483	82	484	83
rect	483	88	484	89
rect	483	91	484	92
rect	483	100	484	101
rect	483	109	484	110
rect	483	121	484	122
rect	483	124	484	125
rect	483	133	484	134
rect	483	136	484	137
rect	483	139	484	140
rect	483	142	484	143
rect	483	145	484	146
rect	483	151	484	152
rect	483	160	484	161
rect	483	163	484	164
rect	483	169	484	170
rect	483	172	484	173
rect	483	175	484	176
rect	483	181	484	182
rect	483	184	484	185
rect	483	187	484	188
rect	483	193	484	194
rect	483	196	484	197
rect	483	208	484	209
rect	483	211	484	212
rect	483	214	484	215
rect	483	217	484	218
rect	483	223	484	224
rect	483	226	484	227
rect	483	229	484	230
rect	483	232	484	233
rect	483	238	484	239
rect	483	244	484	245
rect	483	247	484	248
rect	483	250	484	251
rect	483	253	484	254
rect	483	256	484	257
rect	483	259	484	260
rect	483	265	484	266
rect	483	268	484	269
rect	483	271	484	272
rect	483	274	484	275
rect	483	280	484	281
rect	483	286	484	287
rect	483	292	484	293
rect	483	298	484	299
rect	483	310	484	311
rect	483	331	484	332
rect	483	343	484	344
rect	484	4	485	5
rect	484	7	485	8
rect	484	10	485	11
rect	484	16	485	17
rect	484	22	485	23
rect	484	25	485	26
rect	484	28	485	29
rect	484	34	485	35
rect	484	40	485	41
rect	484	46	485	47
rect	484	49	485	50
rect	484	52	485	53
rect	484	55	485	56
rect	484	58	485	59
rect	484	64	485	65
rect	484	70	485	71
rect	484	73	485	74
rect	484	76	485	77
rect	484	79	485	80
rect	484	82	485	83
rect	484	88	485	89
rect	484	91	485	92
rect	484	100	485	101
rect	484	109	485	110
rect	484	121	485	122
rect	484	124	485	125
rect	484	133	485	134
rect	484	136	485	137
rect	484	139	485	140
rect	484	142	485	143
rect	484	145	485	146
rect	484	151	485	152
rect	484	160	485	161
rect	484	163	485	164
rect	484	169	485	170
rect	484	172	485	173
rect	484	175	485	176
rect	484	181	485	182
rect	484	184	485	185
rect	484	187	485	188
rect	484	193	485	194
rect	484	196	485	197
rect	484	208	485	209
rect	484	211	485	212
rect	484	214	485	215
rect	484	217	485	218
rect	484	223	485	224
rect	484	226	485	227
rect	484	229	485	230
rect	484	232	485	233
rect	484	238	485	239
rect	484	244	485	245
rect	484	247	485	248
rect	484	250	485	251
rect	484	253	485	254
rect	484	256	485	257
rect	484	259	485	260
rect	484	265	485	266
rect	484	268	485	269
rect	484	271	485	272
rect	484	274	485	275
rect	484	280	485	281
rect	484	286	485	287
rect	484	292	485	293
rect	484	298	485	299
rect	484	310	485	311
rect	484	316	485	317
rect	484	331	485	332
rect	484	343	485	344
rect	485	10	486	11
rect	485	16	486	17
rect	485	25	486	26
rect	485	28	486	29
rect	485	34	486	35
rect	485	46	486	47
rect	485	49	486	50
rect	485	55	486	56
rect	485	58	486	59
rect	485	64	486	65
rect	485	70	486	71
rect	485	73	486	74
rect	485	76	486	77
rect	485	79	486	80
rect	485	88	486	89
rect	485	91	486	92
rect	485	100	486	101
rect	485	121	486	122
rect	485	124	486	125
rect	485	133	486	134
rect	485	136	486	137
rect	485	139	486	140
rect	485	142	486	143
rect	485	151	486	152
rect	485	163	486	164
rect	485	169	486	170
rect	485	172	486	173
rect	485	175	486	176
rect	485	181	486	182
rect	485	184	486	185
rect	485	187	486	188
rect	485	196	486	197
rect	485	208	486	209
rect	485	211	486	212
rect	485	214	486	215
rect	485	217	486	218
rect	485	223	486	224
rect	485	226	486	227
rect	485	229	486	230
rect	485	238	486	239
rect	485	244	486	245
rect	485	247	486	248
rect	485	256	486	257
rect	485	259	486	260
rect	485	265	486	266
rect	485	268	486	269
rect	485	271	486	272
rect	485	274	486	275
rect	485	280	486	281
rect	485	286	486	287
rect	485	292	486	293
rect	485	298	486	299
rect	485	310	486	311
rect	485	316	486	317
rect	485	331	486	332
rect	486	10	487	11
rect	486	16	487	17
rect	486	19	487	20
rect	486	25	487	26
rect	486	28	487	29
rect	486	31	487	32
rect	486	34	487	35
rect	486	46	487	47
rect	486	49	487	50
rect	486	55	487	56
rect	486	58	487	59
rect	486	61	487	62
rect	486	64	487	65
rect	486	67	487	68
rect	486	70	487	71
rect	486	73	487	74
rect	486	76	487	77
rect	486	79	487	80
rect	486	88	487	89
rect	486	91	487	92
rect	486	100	487	101
rect	486	103	487	104
rect	486	112	487	113
rect	486	121	487	122
rect	486	124	487	125
rect	486	133	487	134
rect	486	136	487	137
rect	486	139	487	140
rect	486	142	487	143
rect	486	151	487	152
rect	486	154	487	155
rect	486	163	487	164
rect	486	166	487	167
rect	486	169	487	170
rect	486	172	487	173
rect	486	175	487	176
rect	486	181	487	182
rect	486	184	487	185
rect	486	187	487	188
rect	486	196	487	197
rect	486	205	487	206
rect	486	208	487	209
rect	486	211	487	212
rect	486	214	487	215
rect	486	217	487	218
rect	486	223	487	224
rect	486	226	487	227
rect	486	229	487	230
rect	486	235	487	236
rect	486	238	487	239
rect	486	244	487	245
rect	486	247	487	248
rect	486	256	487	257
rect	486	259	487	260
rect	486	265	487	266
rect	486	268	487	269
rect	486	271	487	272
rect	486	274	487	275
rect	486	280	487	281
rect	486	286	487	287
rect	486	292	487	293
rect	486	298	487	299
rect	486	310	487	311
rect	486	316	487	317
rect	486	331	487	332
rect	487	16	488	17
rect	487	19	488	20
rect	487	31	488	32
rect	487	34	488	35
rect	487	46	488	47
rect	487	49	488	50
rect	487	55	488	56
rect	487	58	488	59
rect	487	61	488	62
rect	487	64	488	65
rect	487	67	488	68
rect	487	70	488	71
rect	487	73	488	74
rect	487	76	488	77
rect	487	79	488	80
rect	487	88	488	89
rect	487	91	488	92
rect	487	100	488	101
rect	487	103	488	104
rect	487	112	488	113
rect	487	121	488	122
rect	487	124	488	125
rect	487	133	488	134
rect	487	136	488	137
rect	487	139	488	140
rect	487	142	488	143
rect	487	151	488	152
rect	487	154	488	155
rect	487	163	488	164
rect	487	166	488	167
rect	487	169	488	170
rect	487	172	488	173
rect	487	175	488	176
rect	487	181	488	182
rect	487	184	488	185
rect	487	187	488	188
rect	487	196	488	197
rect	487	205	488	206
rect	487	208	488	209
rect	487	211	488	212
rect	487	214	488	215
rect	487	217	488	218
rect	487	223	488	224
rect	487	226	488	227
rect	487	229	488	230
rect	487	235	488	236
rect	487	238	488	239
rect	487	244	488	245
rect	487	247	488	248
rect	487	256	488	257
rect	487	259	488	260
rect	487	265	488	266
rect	487	268	488	269
rect	487	271	488	272
rect	487	274	488	275
rect	487	286	488	287
rect	487	292	488	293
rect	487	310	488	311
rect	487	316	488	317
rect	488	7	489	8
rect	488	16	489	17
rect	488	19	489	20
rect	488	22	489	23
rect	488	31	489	32
rect	488	34	489	35
rect	488	37	489	38
rect	488	46	489	47
rect	488	49	489	50
rect	488	52	489	53
rect	488	55	489	56
rect	488	58	489	59
rect	488	61	489	62
rect	488	64	489	65
rect	488	67	489	68
rect	488	70	489	71
rect	488	73	489	74
rect	488	76	489	77
rect	488	79	489	80
rect	488	88	489	89
rect	488	91	489	92
rect	488	100	489	101
rect	488	103	489	104
rect	488	112	489	113
rect	488	121	489	122
rect	488	124	489	125
rect	488	133	489	134
rect	488	136	489	137
rect	488	139	489	140
rect	488	142	489	143
rect	488	151	489	152
rect	488	154	489	155
rect	488	163	489	164
rect	488	166	489	167
rect	488	169	489	170
rect	488	172	489	173
rect	488	175	489	176
rect	488	181	489	182
rect	488	184	489	185
rect	488	187	489	188
rect	488	196	489	197
rect	488	205	489	206
rect	488	208	489	209
rect	488	211	489	212
rect	488	214	489	215
rect	488	217	489	218
rect	488	223	489	224
rect	488	226	489	227
rect	488	229	489	230
rect	488	235	489	236
rect	488	238	489	239
rect	488	244	489	245
rect	488	247	489	248
rect	488	256	489	257
rect	488	259	489	260
rect	488	265	489	266
rect	488	268	489	269
rect	488	271	489	272
rect	488	274	489	275
rect	488	283	489	284
rect	488	286	489	287
rect	488	292	489	293
rect	488	307	489	308
rect	488	310	489	311
rect	488	316	489	317
rect	495	1	496	2
rect	495	4	496	5
rect	495	7	496	8
rect	495	13	496	14
rect	495	16	496	17
rect	495	19	496	20
rect	495	22	496	23
rect	495	31	496	32
rect	495	34	496	35
rect	495	37	496	38
rect	495	46	496	47
rect	495	49	496	50
rect	495	52	496	53
rect	495	55	496	56
rect	495	58	496	59
rect	495	61	496	62
rect	495	64	496	65
rect	495	67	496	68
rect	495	70	496	71
rect	495	73	496	74
rect	495	76	496	77
rect	495	79	496	80
rect	495	88	496	89
rect	495	91	496	92
rect	495	100	496	101
rect	495	103	496	104
rect	495	106	496	107
rect	495	112	496	113
rect	495	121	496	122
rect	495	124	496	125
rect	495	130	496	131
rect	495	133	496	134
rect	495	136	496	137
rect	495	139	496	140
rect	495	142	496	143
rect	495	145	496	146
rect	495	151	496	152
rect	495	154	496	155
rect	495	163	496	164
rect	495	166	496	167
rect	495	169	496	170
rect	495	172	496	173
rect	495	181	496	182
rect	495	184	496	185
rect	495	187	496	188
rect	495	196	496	197
rect	495	205	496	206
rect	495	208	496	209
rect	495	211	496	212
rect	495	214	496	215
rect	495	223	496	224
rect	495	226	496	227
rect	495	235	496	236
rect	495	238	496	239
rect	495	244	496	245
rect	495	247	496	248
rect	495	256	496	257
rect	495	259	496	260
rect	495	268	496	269
rect	495	271	496	272
rect	495	274	496	275
rect	495	277	496	278
rect	495	283	496	284
rect	495	292	496	293
rect	495	307	496	308
rect	496	1	497	2
rect	496	4	497	5
rect	496	7	497	8
rect	496	13	497	14
rect	496	16	497	17
rect	496	19	497	20
rect	496	22	497	23
rect	496	31	497	32
rect	496	34	497	35
rect	496	37	497	38
rect	496	46	497	47
rect	496	49	497	50
rect	496	52	497	53
rect	496	55	497	56
rect	496	58	497	59
rect	496	61	497	62
rect	496	64	497	65
rect	496	67	497	68
rect	496	70	497	71
rect	496	73	497	74
rect	496	76	497	77
rect	496	79	497	80
rect	496	88	497	89
rect	496	91	497	92
rect	496	100	497	101
rect	496	103	497	104
rect	496	106	497	107
rect	496	112	497	113
rect	496	121	497	122
rect	496	124	497	125
rect	496	130	497	131
rect	496	133	497	134
rect	496	136	497	137
rect	496	139	497	140
rect	496	142	497	143
rect	496	145	497	146
rect	496	151	497	152
rect	496	154	497	155
rect	496	166	497	167
rect	496	169	497	170
rect	496	172	497	173
rect	496	181	497	182
rect	496	184	497	185
rect	496	187	497	188
rect	496	196	497	197
rect	496	205	497	206
rect	496	208	497	209
rect	496	211	497	212
rect	496	214	497	215
rect	496	223	497	224
rect	496	226	497	227
rect	496	235	497	236
rect	496	238	497	239
rect	496	244	497	245
rect	496	247	497	248
rect	496	256	497	257
rect	496	259	497	260
rect	496	268	497	269
rect	496	271	497	272
rect	496	274	497	275
rect	496	277	497	278
rect	496	283	497	284
rect	496	292	497	293
rect	496	307	497	308
rect	497	1	498	2
rect	497	4	498	5
rect	497	7	498	8
rect	497	13	498	14
rect	497	16	498	17
rect	497	19	498	20
rect	497	22	498	23
rect	497	31	498	32
rect	497	34	498	35
rect	497	37	498	38
rect	497	46	498	47
rect	497	49	498	50
rect	497	52	498	53
rect	497	55	498	56
rect	497	58	498	59
rect	497	61	498	62
rect	497	64	498	65
rect	497	67	498	68
rect	497	70	498	71
rect	497	73	498	74
rect	497	76	498	77
rect	497	79	498	80
rect	497	88	498	89
rect	497	91	498	92
rect	497	100	498	101
rect	497	103	498	104
rect	497	106	498	107
rect	497	112	498	113
rect	497	121	498	122
rect	497	124	498	125
rect	497	130	498	131
rect	497	133	498	134
rect	497	136	498	137
rect	497	139	498	140
rect	497	142	498	143
rect	497	145	498	146
rect	497	151	498	152
rect	497	154	498	155
rect	497	160	498	161
rect	497	166	498	167
rect	497	169	498	170
rect	497	172	498	173
rect	497	181	498	182
rect	497	184	498	185
rect	497	187	498	188
rect	497	196	498	197
rect	497	205	498	206
rect	497	208	498	209
rect	497	211	498	212
rect	497	214	498	215
rect	497	223	498	224
rect	497	226	498	227
rect	497	235	498	236
rect	497	238	498	239
rect	497	244	498	245
rect	497	247	498	248
rect	497	256	498	257
rect	497	259	498	260
rect	497	268	498	269
rect	497	271	498	272
rect	497	274	498	275
rect	497	277	498	278
rect	497	283	498	284
rect	497	292	498	293
rect	497	307	498	308
rect	498	1	499	2
rect	498	7	499	8
rect	498	13	499	14
rect	498	16	499	17
rect	498	19	499	20
rect	498	22	499	23
rect	498	31	499	32
rect	498	34	499	35
rect	498	37	499	38
rect	498	46	499	47
rect	498	49	499	50
rect	498	52	499	53
rect	498	55	499	56
rect	498	58	499	59
rect	498	61	499	62
rect	498	64	499	65
rect	498	67	499	68
rect	498	70	499	71
rect	498	73	499	74
rect	498	76	499	77
rect	498	79	499	80
rect	498	88	499	89
rect	498	91	499	92
rect	498	100	499	101
rect	498	103	499	104
rect	498	106	499	107
rect	498	112	499	113
rect	498	121	499	122
rect	498	124	499	125
rect	498	130	499	131
rect	498	133	499	134
rect	498	136	499	137
rect	498	139	499	140
rect	498	142	499	143
rect	498	145	499	146
rect	498	151	499	152
rect	498	154	499	155
rect	498	160	499	161
rect	498	166	499	167
rect	498	169	499	170
rect	498	172	499	173
rect	498	181	499	182
rect	498	184	499	185
rect	498	187	499	188
rect	498	196	499	197
rect	498	205	499	206
rect	498	211	499	212
rect	498	214	499	215
rect	498	223	499	224
rect	498	226	499	227
rect	498	235	499	236
rect	498	238	499	239
rect	498	244	499	245
rect	498	247	499	248
rect	498	256	499	257
rect	498	259	499	260
rect	498	268	499	269
rect	498	271	499	272
rect	498	274	499	275
rect	498	277	499	278
rect	498	283	499	284
rect	498	292	499	293
rect	498	307	499	308
rect	499	1	500	2
rect	499	7	500	8
rect	499	13	500	14
rect	499	16	500	17
rect	499	19	500	20
rect	499	22	500	23
rect	499	31	500	32
rect	499	34	500	35
rect	499	37	500	38
rect	499	46	500	47
rect	499	49	500	50
rect	499	52	500	53
rect	499	55	500	56
rect	499	58	500	59
rect	499	61	500	62
rect	499	64	500	65
rect	499	67	500	68
rect	499	70	500	71
rect	499	73	500	74
rect	499	76	500	77
rect	499	79	500	80
rect	499	88	500	89
rect	499	91	500	92
rect	499	100	500	101
rect	499	103	500	104
rect	499	106	500	107
rect	499	112	500	113
rect	499	121	500	122
rect	499	124	500	125
rect	499	130	500	131
rect	499	133	500	134
rect	499	136	500	137
rect	499	139	500	140
rect	499	142	500	143
rect	499	145	500	146
rect	499	151	500	152
rect	499	154	500	155
rect	499	160	500	161
rect	499	166	500	167
rect	499	169	500	170
rect	499	172	500	173
rect	499	181	500	182
rect	499	184	500	185
rect	499	187	500	188
rect	499	196	500	197
rect	499	205	500	206
rect	499	211	500	212
rect	499	214	500	215
rect	499	223	500	224
rect	499	226	500	227
rect	499	235	500	236
rect	499	238	500	239
rect	499	244	500	245
rect	499	247	500	248
rect	499	256	500	257
rect	499	259	500	260
rect	499	268	500	269
rect	499	271	500	272
rect	499	274	500	275
rect	499	277	500	278
rect	499	283	500	284
rect	499	292	500	293
rect	499	307	500	308
rect	500	1	501	2
rect	500	7	501	8
rect	500	13	501	14
rect	500	16	501	17
rect	500	19	501	20
rect	500	22	501	23
rect	500	31	501	32
rect	500	34	501	35
rect	500	37	501	38
rect	500	46	501	47
rect	500	49	501	50
rect	500	52	501	53
rect	500	55	501	56
rect	500	58	501	59
rect	500	61	501	62
rect	500	64	501	65
rect	500	67	501	68
rect	500	70	501	71
rect	500	73	501	74
rect	500	76	501	77
rect	500	79	501	80
rect	500	88	501	89
rect	500	91	501	92
rect	500	100	501	101
rect	500	103	501	104
rect	500	106	501	107
rect	500	112	501	113
rect	500	121	501	122
rect	500	124	501	125
rect	500	130	501	131
rect	500	133	501	134
rect	500	136	501	137
rect	500	139	501	140
rect	500	142	501	143
rect	500	145	501	146
rect	500	151	501	152
rect	500	154	501	155
rect	500	160	501	161
rect	500	166	501	167
rect	500	169	501	170
rect	500	172	501	173
rect	500	181	501	182
rect	500	184	501	185
rect	500	187	501	188
rect	500	205	501	206
rect	500	211	501	212
rect	500	214	501	215
rect	500	223	501	224
rect	500	226	501	227
rect	500	235	501	236
rect	500	238	501	239
rect	500	244	501	245
rect	500	247	501	248
rect	500	256	501	257
rect	500	259	501	260
rect	500	268	501	269
rect	500	271	501	272
rect	500	274	501	275
rect	500	277	501	278
rect	500	283	501	284
rect	500	292	501	293
rect	500	307	501	308
rect	501	1	502	2
rect	501	7	502	8
rect	501	13	502	14
rect	501	16	502	17
rect	501	19	502	20
rect	501	22	502	23
rect	501	31	502	32
rect	501	34	502	35
rect	501	37	502	38
rect	501	46	502	47
rect	501	49	502	50
rect	501	52	502	53
rect	501	55	502	56
rect	501	58	502	59
rect	501	61	502	62
rect	501	64	502	65
rect	501	67	502	68
rect	501	70	502	71
rect	501	73	502	74
rect	501	76	502	77
rect	501	79	502	80
rect	501	88	502	89
rect	501	91	502	92
rect	501	100	502	101
rect	501	103	502	104
rect	501	106	502	107
rect	501	112	502	113
rect	501	121	502	122
rect	501	124	502	125
rect	501	130	502	131
rect	501	133	502	134
rect	501	136	502	137
rect	501	139	502	140
rect	501	142	502	143
rect	501	145	502	146
rect	501	151	502	152
rect	501	154	502	155
rect	501	160	502	161
rect	501	163	502	164
rect	501	166	502	167
rect	501	169	502	170
rect	501	172	502	173
rect	501	181	502	182
rect	501	184	502	185
rect	501	187	502	188
rect	501	199	502	200
rect	501	205	502	206
rect	501	208	502	209
rect	501	211	502	212
rect	501	214	502	215
rect	501	223	502	224
rect	501	226	502	227
rect	501	235	502	236
rect	501	238	502	239
rect	501	244	502	245
rect	501	247	502	248
rect	501	256	502	257
rect	501	259	502	260
rect	501	268	502	269
rect	501	271	502	272
rect	501	274	502	275
rect	501	277	502	278
rect	501	283	502	284
rect	501	292	502	293
rect	501	307	502	308
rect	502	1	503	2
rect	502	7	503	8
rect	502	13	503	14
rect	502	16	503	17
rect	502	19	503	20
rect	502	22	503	23
rect	502	31	503	32
rect	502	34	503	35
rect	502	37	503	38
rect	502	46	503	47
rect	502	49	503	50
rect	502	52	503	53
rect	502	55	503	56
rect	502	58	503	59
rect	502	61	503	62
rect	502	64	503	65
rect	502	67	503	68
rect	502	70	503	71
rect	502	73	503	74
rect	502	76	503	77
rect	502	79	503	80
rect	502	88	503	89
rect	502	91	503	92
rect	502	100	503	101
rect	502	103	503	104
rect	502	106	503	107
rect	502	112	503	113
rect	502	121	503	122
rect	502	124	503	125
rect	502	130	503	131
rect	502	133	503	134
rect	502	136	503	137
rect	502	139	503	140
rect	502	142	503	143
rect	502	145	503	146
rect	502	151	503	152
rect	502	154	503	155
rect	502	160	503	161
rect	502	163	503	164
rect	502	166	503	167
rect	502	169	503	170
rect	502	172	503	173
rect	502	181	503	182
rect	502	184	503	185
rect	502	187	503	188
rect	502	199	503	200
rect	502	205	503	206
rect	502	208	503	209
rect	502	214	503	215
rect	502	223	503	224
rect	502	226	503	227
rect	502	235	503	236
rect	502	238	503	239
rect	502	244	503	245
rect	502	247	503	248
rect	502	256	503	257
rect	502	259	503	260
rect	502	268	503	269
rect	502	271	503	272
rect	502	274	503	275
rect	502	277	503	278
rect	502	283	503	284
rect	502	292	503	293
rect	502	307	503	308
rect	503	1	504	2
rect	503	7	504	8
rect	503	13	504	14
rect	503	16	504	17
rect	503	19	504	20
rect	503	22	504	23
rect	503	31	504	32
rect	503	34	504	35
rect	503	37	504	38
rect	503	46	504	47
rect	503	49	504	50
rect	503	52	504	53
rect	503	55	504	56
rect	503	58	504	59
rect	503	61	504	62
rect	503	64	504	65
rect	503	67	504	68
rect	503	70	504	71
rect	503	73	504	74
rect	503	76	504	77
rect	503	79	504	80
rect	503	88	504	89
rect	503	91	504	92
rect	503	100	504	101
rect	503	103	504	104
rect	503	106	504	107
rect	503	112	504	113
rect	503	121	504	122
rect	503	124	504	125
rect	503	130	504	131
rect	503	133	504	134
rect	503	136	504	137
rect	503	139	504	140
rect	503	142	504	143
rect	503	145	504	146
rect	503	151	504	152
rect	503	154	504	155
rect	503	160	504	161
rect	503	163	504	164
rect	503	166	504	167
rect	503	169	504	170
rect	503	172	504	173
rect	503	181	504	182
rect	503	184	504	185
rect	503	187	504	188
rect	503	196	504	197
rect	503	199	504	200
rect	503	205	504	206
rect	503	208	504	209
rect	503	214	504	215
rect	503	223	504	224
rect	503	226	504	227
rect	503	235	504	236
rect	503	238	504	239
rect	503	244	504	245
rect	503	247	504	248
rect	503	256	504	257
rect	503	259	504	260
rect	503	268	504	269
rect	503	271	504	272
rect	503	274	504	275
rect	503	277	504	278
rect	503	283	504	284
rect	503	292	504	293
rect	503	307	504	308
rect	504	1	505	2
rect	504	7	505	8
rect	504	13	505	14
rect	504	16	505	17
rect	504	19	505	20
rect	504	22	505	23
rect	504	31	505	32
rect	504	34	505	35
rect	504	37	505	38
rect	504	46	505	47
rect	504	49	505	50
rect	504	52	505	53
rect	504	55	505	56
rect	504	58	505	59
rect	504	61	505	62
rect	504	64	505	65
rect	504	67	505	68
rect	504	70	505	71
rect	504	73	505	74
rect	504	76	505	77
rect	504	79	505	80
rect	504	88	505	89
rect	504	91	505	92
rect	504	100	505	101
rect	504	103	505	104
rect	504	106	505	107
rect	504	112	505	113
rect	504	121	505	122
rect	504	124	505	125
rect	504	130	505	131
rect	504	133	505	134
rect	504	136	505	137
rect	504	139	505	140
rect	504	142	505	143
rect	504	145	505	146
rect	504	151	505	152
rect	504	154	505	155
rect	504	160	505	161
rect	504	163	505	164
rect	504	166	505	167
rect	504	169	505	170
rect	504	172	505	173
rect	504	181	505	182
rect	504	184	505	185
rect	504	187	505	188
rect	504	196	505	197
rect	504	199	505	200
rect	504	205	505	206
rect	504	208	505	209
rect	504	214	505	215
rect	504	223	505	224
rect	504	226	505	227
rect	504	238	505	239
rect	504	244	505	245
rect	504	247	505	248
rect	504	256	505	257
rect	504	259	505	260
rect	504	268	505	269
rect	504	271	505	272
rect	504	274	505	275
rect	504	292	505	293
rect	504	307	505	308
rect	505	1	506	2
rect	505	7	506	8
rect	505	13	506	14
rect	505	16	506	17
rect	505	19	506	20
rect	505	22	506	23
rect	505	31	506	32
rect	505	34	506	35
rect	505	37	506	38
rect	505	46	506	47
rect	505	49	506	50
rect	505	52	506	53
rect	505	55	506	56
rect	505	58	506	59
rect	505	61	506	62
rect	505	64	506	65
rect	505	67	506	68
rect	505	70	506	71
rect	505	73	506	74
rect	505	76	506	77
rect	505	79	506	80
rect	505	88	506	89
rect	505	91	506	92
rect	505	100	506	101
rect	505	103	506	104
rect	505	106	506	107
rect	505	112	506	113
rect	505	121	506	122
rect	505	124	506	125
rect	505	130	506	131
rect	505	133	506	134
rect	505	136	506	137
rect	505	139	506	140
rect	505	142	506	143
rect	505	145	506	146
rect	505	151	506	152
rect	505	154	506	155
rect	505	160	506	161
rect	505	163	506	164
rect	505	166	506	167
rect	505	169	506	170
rect	505	172	506	173
rect	505	181	506	182
rect	505	184	506	185
rect	505	187	506	188
rect	505	190	506	191
rect	505	196	506	197
rect	505	199	506	200
rect	505	205	506	206
rect	505	208	506	209
rect	505	214	506	215
rect	505	223	506	224
rect	505	226	506	227
rect	505	238	506	239
rect	505	244	506	245
rect	505	247	506	248
rect	505	256	506	257
rect	505	259	506	260
rect	505	268	506	269
rect	505	271	506	272
rect	505	274	506	275
rect	505	292	506	293
rect	505	307	506	308
rect	506	1	507	2
rect	506	7	507	8
rect	506	13	507	14
rect	506	16	507	17
rect	506	19	507	20
rect	506	22	507	23
rect	506	31	507	32
rect	506	34	507	35
rect	506	37	507	38
rect	506	46	507	47
rect	506	52	507	53
rect	506	55	507	56
rect	506	58	507	59
rect	506	61	507	62
rect	506	64	507	65
rect	506	67	507	68
rect	506	70	507	71
rect	506	73	507	74
rect	506	76	507	77
rect	506	79	507	80
rect	506	88	507	89
rect	506	91	507	92
rect	506	100	507	101
rect	506	103	507	104
rect	506	106	507	107
rect	506	112	507	113
rect	506	121	507	122
rect	506	124	507	125
rect	506	130	507	131
rect	506	133	507	134
rect	506	136	507	137
rect	506	139	507	140
rect	506	142	507	143
rect	506	145	507	146
rect	506	151	507	152
rect	506	154	507	155
rect	506	160	507	161
rect	506	163	507	164
rect	506	166	507	167
rect	506	169	507	170
rect	506	172	507	173
rect	506	184	507	185
rect	506	187	507	188
rect	506	190	507	191
rect	506	196	507	197
rect	506	199	507	200
rect	506	205	507	206
rect	506	208	507	209
rect	506	214	507	215
rect	506	223	507	224
rect	506	226	507	227
rect	506	238	507	239
rect	506	244	507	245
rect	506	247	507	248
rect	506	256	507	257
rect	506	259	507	260
rect	506	268	507	269
rect	506	271	507	272
rect	506	274	507	275
rect	506	292	507	293
rect	506	307	507	308
rect	507	1	508	2
rect	507	7	508	8
rect	507	13	508	14
rect	507	16	508	17
rect	507	19	508	20
rect	507	22	508	23
rect	507	28	508	29
rect	507	31	508	32
rect	507	34	508	35
rect	507	37	508	38
rect	507	46	508	47
rect	507	52	508	53
rect	507	55	508	56
rect	507	58	508	59
rect	507	61	508	62
rect	507	64	508	65
rect	507	67	508	68
rect	507	70	508	71
rect	507	73	508	74
rect	507	76	508	77
rect	507	79	508	80
rect	507	88	508	89
rect	507	91	508	92
rect	507	100	508	101
rect	507	103	508	104
rect	507	106	508	107
rect	507	112	508	113
rect	507	121	508	122
rect	507	124	508	125
rect	507	130	508	131
rect	507	133	508	134
rect	507	136	508	137
rect	507	139	508	140
rect	507	142	508	143
rect	507	145	508	146
rect	507	151	508	152
rect	507	154	508	155
rect	507	160	508	161
rect	507	163	508	164
rect	507	166	508	167
rect	507	169	508	170
rect	507	172	508	173
rect	507	184	508	185
rect	507	187	508	188
rect	507	190	508	191
rect	507	196	508	197
rect	507	199	508	200
rect	507	205	508	206
rect	507	208	508	209
rect	507	214	508	215
rect	507	223	508	224
rect	507	226	508	227
rect	507	238	508	239
rect	507	244	508	245
rect	507	247	508	248
rect	507	256	508	257
rect	507	259	508	260
rect	507	268	508	269
rect	507	271	508	272
rect	507	274	508	275
rect	507	277	508	278
rect	507	292	508	293
rect	507	307	508	308
rect	508	1	509	2
rect	508	7	509	8
rect	508	13	509	14
rect	508	16	509	17
rect	508	19	509	20
rect	508	22	509	23
rect	508	28	509	29
rect	508	31	509	32
rect	508	34	509	35
rect	508	37	509	38
rect	508	52	509	53
rect	508	55	509	56
rect	508	58	509	59
rect	508	61	509	62
rect	508	64	509	65
rect	508	70	509	71
rect	508	73	509	74
rect	508	76	509	77
rect	508	79	509	80
rect	508	88	509	89
rect	508	91	509	92
rect	508	100	509	101
rect	508	103	509	104
rect	508	106	509	107
rect	508	112	509	113
rect	508	121	509	122
rect	508	124	509	125
rect	508	130	509	131
rect	508	133	509	134
rect	508	136	509	137
rect	508	139	509	140
rect	508	142	509	143
rect	508	154	509	155
rect	508	160	509	161
rect	508	163	509	164
rect	508	166	509	167
rect	508	169	509	170
rect	508	172	509	173
rect	508	184	509	185
rect	508	187	509	188
rect	508	190	509	191
rect	508	196	509	197
rect	508	199	509	200
rect	508	205	509	206
rect	508	208	509	209
rect	508	214	509	215
rect	508	223	509	224
rect	508	244	509	245
rect	508	256	509	257
rect	508	259	509	260
rect	508	268	509	269
rect	508	271	509	272
rect	508	274	509	275
rect	508	277	509	278
rect	508	292	509	293
rect	508	307	509	308
rect	509	1	510	2
rect	509	7	510	8
rect	509	13	510	14
rect	509	16	510	17
rect	509	19	510	20
rect	509	22	510	23
rect	509	25	510	26
rect	509	28	510	29
rect	509	31	510	32
rect	509	34	510	35
rect	509	37	510	38
rect	509	49	510	50
rect	509	52	510	53
rect	509	55	510	56
rect	509	58	510	59
rect	509	61	510	62
rect	509	64	510	65
rect	509	70	510	71
rect	509	73	510	74
rect	509	76	510	77
rect	509	79	510	80
rect	509	88	510	89
rect	509	91	510	92
rect	509	100	510	101
rect	509	103	510	104
rect	509	106	510	107
rect	509	112	510	113
rect	509	121	510	122
rect	509	124	510	125
rect	509	130	510	131
rect	509	133	510	134
rect	509	136	510	137
rect	509	139	510	140
rect	509	142	510	143
rect	509	154	510	155
rect	509	160	510	161
rect	509	163	510	164
rect	509	166	510	167
rect	509	169	510	170
rect	509	172	510	173
rect	509	178	510	179
rect	509	184	510	185
rect	509	187	510	188
rect	509	190	510	191
rect	509	196	510	197
rect	509	199	510	200
rect	509	205	510	206
rect	509	208	510	209
rect	509	214	510	215
rect	509	223	510	224
rect	509	244	510	245
rect	509	256	510	257
rect	509	259	510	260
rect	509	268	510	269
rect	509	271	510	272
rect	509	274	510	275
rect	509	277	510	278
rect	509	292	510	293
rect	509	307	510	308
rect	510	1	511	2
rect	510	7	511	8
rect	510	13	511	14
rect	510	16	511	17
rect	510	19	511	20
rect	510	22	511	23
rect	510	25	511	26
rect	510	28	511	29
rect	510	31	511	32
rect	510	34	511	35
rect	510	37	511	38
rect	510	49	511	50
rect	510	52	511	53
rect	510	55	511	56
rect	510	58	511	59
rect	510	61	511	62
rect	510	70	511	71
rect	510	73	511	74
rect	510	76	511	77
rect	510	79	511	80
rect	510	88	511	89
rect	510	91	511	92
rect	510	100	511	101
rect	510	103	511	104
rect	510	106	511	107
rect	510	112	511	113
rect	510	121	511	122
rect	510	124	511	125
rect	510	130	511	131
rect	510	133	511	134
rect	510	136	511	137
rect	510	139	511	140
rect	510	142	511	143
rect	510	154	511	155
rect	510	160	511	161
rect	510	163	511	164
rect	510	169	511	170
rect	510	172	511	173
rect	510	178	511	179
rect	510	184	511	185
rect	510	187	511	188
rect	510	190	511	191
rect	510	196	511	197
rect	510	199	511	200
rect	510	208	511	209
rect	510	214	511	215
rect	510	223	511	224
rect	510	244	511	245
rect	510	256	511	257
rect	510	259	511	260
rect	510	268	511	269
rect	510	274	511	275
rect	510	277	511	278
rect	510	292	511	293
rect	510	307	511	308
rect	511	1	512	2
rect	511	7	512	8
rect	511	13	512	14
rect	511	16	512	17
rect	511	19	512	20
rect	511	22	512	23
rect	511	25	512	26
rect	511	28	512	29
rect	511	31	512	32
rect	511	34	512	35
rect	511	37	512	38
rect	511	46	512	47
rect	511	49	512	50
rect	511	52	512	53
rect	511	55	512	56
rect	511	58	512	59
rect	511	61	512	62
rect	511	70	512	71
rect	511	73	512	74
rect	511	76	512	77
rect	511	79	512	80
rect	511	88	512	89
rect	511	91	512	92
rect	511	100	512	101
rect	511	103	512	104
rect	511	106	512	107
rect	511	112	512	113
rect	511	121	512	122
rect	511	124	512	125
rect	511	130	512	131
rect	511	133	512	134
rect	511	136	512	137
rect	511	139	512	140
rect	511	142	512	143
rect	511	151	512	152
rect	511	154	512	155
rect	511	160	512	161
rect	511	163	512	164
rect	511	169	512	170
rect	511	172	512	173
rect	511	175	512	176
rect	511	178	512	179
rect	511	184	512	185
rect	511	187	512	188
rect	511	190	512	191
rect	511	196	512	197
rect	511	199	512	200
rect	511	208	512	209
rect	511	214	512	215
rect	511	223	512	224
rect	511	238	512	239
rect	511	244	512	245
rect	511	256	512	257
rect	511	259	512	260
rect	511	268	512	269
rect	511	274	512	275
rect	511	277	512	278
rect	511	292	512	293
rect	511	307	512	308
rect	512	1	513	2
rect	512	7	513	8
rect	512	13	513	14
rect	512	16	513	17
rect	512	19	513	20
rect	512	22	513	23
rect	512	25	513	26
rect	512	28	513	29
rect	512	31	513	32
rect	512	34	513	35
rect	512	37	513	38
rect	512	46	513	47
rect	512	49	513	50
rect	512	52	513	53
rect	512	55	513	56
rect	512	58	513	59
rect	512	70	513	71
rect	512	73	513	74
rect	512	76	513	77
rect	512	79	513	80
rect	512	91	513	92
rect	512	100	513	101
rect	512	103	513	104
rect	512	106	513	107
rect	512	112	513	113
rect	512	121	513	122
rect	512	124	513	125
rect	512	130	513	131
rect	512	133	513	134
rect	512	136	513	137
rect	512	139	513	140
rect	512	142	513	143
rect	512	151	513	152
rect	512	154	513	155
rect	512	160	513	161
rect	512	163	513	164
rect	512	175	513	176
rect	512	178	513	179
rect	512	187	513	188
rect	512	190	513	191
rect	512	196	513	197
rect	512	199	513	200
rect	512	208	513	209
rect	512	214	513	215
rect	512	223	513	224
rect	512	238	513	239
rect	512	256	513	257
rect	512	259	513	260
rect	512	268	513	269
rect	512	277	513	278
rect	512	292	513	293
rect	512	307	513	308
rect	513	1	514	2
rect	513	7	514	8
rect	513	13	514	14
rect	513	16	514	17
rect	513	19	514	20
rect	513	22	514	23
rect	513	25	514	26
rect	513	28	514	29
rect	513	31	514	32
rect	513	34	514	35
rect	513	37	514	38
rect	513	43	514	44
rect	513	46	514	47
rect	513	49	514	50
rect	513	52	514	53
rect	513	55	514	56
rect	513	58	514	59
rect	513	70	514	71
rect	513	73	514	74
rect	513	76	514	77
rect	513	79	514	80
rect	513	85	514	86
rect	513	91	514	92
rect	513	100	514	101
rect	513	103	514	104
rect	513	106	514	107
rect	513	112	514	113
rect	513	121	514	122
rect	513	124	514	125
rect	513	130	514	131
rect	513	133	514	134
rect	513	136	514	137
rect	513	139	514	140
rect	513	142	514	143
rect	513	151	514	152
rect	513	154	514	155
rect	513	160	514	161
rect	513	163	514	164
rect	513	166	514	167
rect	513	175	514	176
rect	513	178	514	179
rect	513	181	514	182
rect	513	187	514	188
rect	513	190	514	191
rect	513	196	514	197
rect	513	199	514	200
rect	513	202	514	203
rect	513	208	514	209
rect	513	211	514	212
rect	513	214	514	215
rect	513	223	514	224
rect	513	238	514	239
rect	513	247	514	248
rect	513	256	514	257
rect	513	259	514	260
rect	513	268	514	269
rect	513	277	514	278
rect	513	292	514	293
rect	513	307	514	308
rect	514	1	515	2
rect	514	7	515	8
rect	514	13	515	14
rect	514	16	515	17
rect	514	19	515	20
rect	514	22	515	23
rect	514	25	515	26
rect	514	28	515	29
rect	514	31	515	32
rect	514	34	515	35
rect	514	37	515	38
rect	514	43	515	44
rect	514	46	515	47
rect	514	49	515	50
rect	514	52	515	53
rect	514	55	515	56
rect	514	70	515	71
rect	514	73	515	74
rect	514	76	515	77
rect	514	79	515	80
rect	514	85	515	86
rect	514	91	515	92
rect	514	103	515	104
rect	514	106	515	107
rect	514	112	515	113
rect	514	121	515	122
rect	514	124	515	125
rect	514	133	515	134
rect	514	136	515	137
rect	514	142	515	143
rect	514	151	515	152
rect	514	160	515	161
rect	514	163	515	164
rect	514	166	515	167
rect	514	175	515	176
rect	514	178	515	179
rect	514	181	515	182
rect	514	190	515	191
rect	514	196	515	197
rect	514	199	515	200
rect	514	202	515	203
rect	514	208	515	209
rect	514	211	515	212
rect	514	214	515	215
rect	514	238	515	239
rect	514	247	515	248
rect	514	259	515	260
rect	514	268	515	269
rect	514	277	515	278
rect	514	292	515	293
rect	514	307	515	308
rect	515	1	516	2
rect	515	7	516	8
rect	515	13	516	14
rect	515	16	516	17
rect	515	19	516	20
rect	515	22	516	23
rect	515	25	516	26
rect	515	28	516	29
rect	515	31	516	32
rect	515	34	516	35
rect	515	37	516	38
rect	515	40	516	41
rect	515	43	516	44
rect	515	46	516	47
rect	515	49	516	50
rect	515	52	516	53
rect	515	55	516	56
rect	515	70	516	71
rect	515	73	516	74
rect	515	76	516	77
rect	515	79	516	80
rect	515	82	516	83
rect	515	85	516	86
rect	515	91	516	92
rect	515	103	516	104
rect	515	106	516	107
rect	515	112	516	113
rect	515	121	516	122
rect	515	124	516	125
rect	515	133	516	134
rect	515	136	516	137
rect	515	142	516	143
rect	515	148	516	149
rect	515	151	516	152
rect	515	160	516	161
rect	515	163	516	164
rect	515	166	516	167
rect	515	169	516	170
rect	515	175	516	176
rect	515	178	516	179
rect	515	181	516	182
rect	515	190	516	191
rect	515	193	516	194
rect	515	196	516	197
rect	515	199	516	200
rect	515	202	516	203
rect	515	208	516	209
rect	515	211	516	212
rect	515	214	516	215
rect	515	235	516	236
rect	515	238	516	239
rect	515	247	516	248
rect	515	259	516	260
rect	515	268	516	269
rect	515	277	516	278
rect	515	292	516	293
rect	515	307	516	308
rect	516	1	517	2
rect	516	7	517	8
rect	516	13	517	14
rect	516	16	517	17
rect	516	19	517	20
rect	516	22	517	23
rect	516	25	517	26
rect	516	28	517	29
rect	516	31	517	32
rect	516	37	517	38
rect	516	40	517	41
rect	516	43	517	44
rect	516	46	517	47
rect	516	49	517	50
rect	516	52	517	53
rect	516	55	517	56
rect	516	70	517	71
rect	516	76	517	77
rect	516	79	517	80
rect	516	82	517	83
rect	516	85	517	86
rect	516	91	517	92
rect	516	103	517	104
rect	516	112	517	113
rect	516	121	517	122
rect	516	124	517	125
rect	516	133	517	134
rect	516	136	517	137
rect	516	142	517	143
rect	516	148	517	149
rect	516	151	517	152
rect	516	160	517	161
rect	516	163	517	164
rect	516	166	517	167
rect	516	169	517	170
rect	516	175	517	176
rect	516	178	517	179
rect	516	181	517	182
rect	516	190	517	191
rect	516	193	517	194
rect	516	196	517	197
rect	516	199	517	200
rect	516	202	517	203
rect	516	208	517	209
rect	516	211	517	212
rect	516	214	517	215
rect	516	235	517	236
rect	516	238	517	239
rect	516	247	517	248
rect	516	259	517	260
rect	516	277	517	278
rect	516	292	517	293
rect	516	307	517	308
rect	517	1	518	2
rect	517	7	518	8
rect	517	13	518	14
rect	517	16	518	17
rect	517	19	518	20
rect	517	22	518	23
rect	517	25	518	26
rect	517	28	518	29
rect	517	31	518	32
rect	517	37	518	38
rect	517	40	518	41
rect	517	43	518	44
rect	517	46	518	47
rect	517	49	518	50
rect	517	52	518	53
rect	517	55	518	56
rect	517	64	518	65
rect	517	70	518	71
rect	517	76	518	77
rect	517	79	518	80
rect	517	82	518	83
rect	517	85	518	86
rect	517	91	518	92
rect	517	103	518	104
rect	517	112	518	113
rect	517	121	518	122
rect	517	124	518	125
rect	517	130	518	131
rect	517	133	518	134
rect	517	136	518	137
rect	517	142	518	143
rect	517	148	518	149
rect	517	151	518	152
rect	517	160	518	161
rect	517	163	518	164
rect	517	166	518	167
rect	517	169	518	170
rect	517	175	518	176
rect	517	178	518	179
rect	517	181	518	182
rect	517	190	518	191
rect	517	193	518	194
rect	517	196	518	197
rect	517	199	518	200
rect	517	202	518	203
rect	517	208	518	209
rect	517	211	518	212
rect	517	214	518	215
rect	517	235	518	236
rect	517	238	518	239
rect	517	247	518	248
rect	517	259	518	260
rect	517	277	518	278
rect	517	292	518	293
rect	517	307	518	308
rect	518	1	519	2
rect	518	7	519	8
rect	518	16	519	17
rect	518	22	519	23
rect	518	25	519	26
rect	518	28	519	29
rect	518	31	519	32
rect	518	37	519	38
rect	518	40	519	41
rect	518	43	519	44
rect	518	46	519	47
rect	518	49	519	50
rect	518	55	519	56
rect	518	64	519	65
rect	518	76	519	77
rect	518	82	519	83
rect	518	85	519	86
rect	518	103	519	104
rect	518	121	519	122
rect	518	124	519	125
rect	518	130	519	131
rect	518	133	519	134
rect	518	148	519	149
rect	518	151	519	152
rect	518	160	519	161
rect	518	163	519	164
rect	518	166	519	167
rect	518	169	519	170
rect	518	175	519	176
rect	518	178	519	179
rect	518	181	519	182
rect	518	190	519	191
rect	518	193	519	194
rect	518	196	519	197
rect	518	199	519	200
rect	518	202	519	203
rect	518	208	519	209
rect	518	211	519	212
rect	518	214	519	215
rect	518	235	519	236
rect	518	238	519	239
rect	518	247	519	248
rect	518	259	519	260
rect	518	277	519	278
rect	518	292	519	293
rect	518	307	519	308
rect	519	1	520	2
rect	519	7	520	8
rect	519	16	520	17
rect	519	22	520	23
rect	519	25	520	26
rect	519	28	520	29
rect	519	31	520	32
rect	519	34	520	35
rect	519	37	520	38
rect	519	40	520	41
rect	519	43	520	44
rect	519	46	520	47
rect	519	49	520	50
rect	519	55	520	56
rect	519	61	520	62
rect	519	64	520	65
rect	519	73	520	74
rect	519	76	520	77
rect	519	82	520	83
rect	519	85	520	86
rect	519	88	520	89
rect	519	100	520	101
rect	519	103	520	104
rect	519	118	520	119
rect	519	121	520	122
rect	519	124	520	125
rect	519	130	520	131
rect	519	133	520	134
rect	519	148	520	149
rect	519	151	520	152
rect	519	160	520	161
rect	519	163	520	164
rect	519	166	520	167
rect	519	169	520	170
rect	519	175	520	176
rect	519	178	520	179
rect	519	181	520	182
rect	519	190	520	191
rect	519	193	520	194
rect	519	196	520	197
rect	519	199	520	200
rect	519	202	520	203
rect	519	208	520	209
rect	519	211	520	212
rect	519	214	520	215
rect	519	235	520	236
rect	519	238	520	239
rect	519	247	520	248
rect	519	250	520	251
rect	519	259	520	260
rect	519	277	520	278
rect	519	292	520	293
rect	519	307	520	308
rect	520	16	521	17
rect	520	25	521	26
rect	520	28	521	29
rect	520	31	521	32
rect	520	34	521	35
rect	520	40	521	41
rect	520	43	521	44
rect	520	46	521	47
rect	520	49	521	50
rect	520	55	521	56
rect	520	61	521	62
rect	520	64	521	65
rect	520	73	521	74
rect	520	76	521	77
rect	520	82	521	83
rect	520	85	521	86
rect	520	88	521	89
rect	520	100	521	101
rect	520	103	521	104
rect	520	118	521	119
rect	520	121	521	122
rect	520	124	521	125
rect	520	130	521	131
rect	520	133	521	134
rect	520	148	521	149
rect	520	151	521	152
rect	520	160	521	161
rect	520	163	521	164
rect	520	166	521	167
rect	520	169	521	170
rect	520	175	521	176
rect	520	178	521	179
rect	520	181	521	182
rect	520	190	521	191
rect	520	193	521	194
rect	520	196	521	197
rect	520	199	521	200
rect	520	202	521	203
rect	520	208	521	209
rect	520	211	521	212
rect	520	214	521	215
rect	520	235	521	236
rect	520	238	521	239
rect	520	247	521	248
rect	520	250	521	251
rect	520	259	521	260
rect	520	277	521	278
rect	520	292	521	293
rect	521	13	522	14
rect	521	16	522	17
rect	521	25	522	26
rect	521	28	522	29
rect	521	31	522	32
rect	521	34	522	35
rect	521	40	522	41
rect	521	43	522	44
rect	521	46	522	47
rect	521	49	522	50
rect	521	52	522	53
rect	521	55	522	56
rect	521	61	522	62
rect	521	64	522	65
rect	521	70	522	71
rect	521	73	522	74
rect	521	76	522	77
rect	521	82	522	83
rect	521	85	522	86
rect	521	88	522	89
rect	521	100	522	101
rect	521	103	522	104
rect	521	118	522	119
rect	521	121	522	122
rect	521	124	522	125
rect	521	130	522	131
rect	521	133	522	134
rect	521	148	522	149
rect	521	151	522	152
rect	521	160	522	161
rect	521	163	522	164
rect	521	166	522	167
rect	521	169	522	170
rect	521	175	522	176
rect	521	178	522	179
rect	521	181	522	182
rect	521	190	522	191
rect	521	193	522	194
rect	521	196	522	197
rect	521	199	522	200
rect	521	202	522	203
rect	521	208	522	209
rect	521	211	522	212
rect	521	214	522	215
rect	521	235	522	236
rect	521	238	522	239
rect	521	241	522	242
rect	521	247	522	248
rect	521	250	522	251
rect	521	259	522	260
rect	521	274	522	275
rect	521	277	522	278
rect	521	292	522	293
rect	522	13	523	14
rect	522	25	523	26
rect	522	28	523	29
rect	522	31	523	32
rect	522	34	523	35
rect	522	40	523	41
rect	522	43	523	44
rect	522	46	523	47
rect	522	49	523	50
rect	522	52	523	53
rect	522	61	523	62
rect	522	64	523	65
rect	522	70	523	71
rect	522	73	523	74
rect	522	82	523	83
rect	522	85	523	86
rect	522	88	523	89
rect	522	100	523	101
rect	522	118	523	119
rect	522	121	523	122
rect	522	124	523	125
rect	522	130	523	131
rect	522	148	523	149
rect	522	151	523	152
rect	522	160	523	161
rect	522	163	523	164
rect	522	166	523	167
rect	522	169	523	170
rect	522	175	523	176
rect	522	178	523	179
rect	522	181	523	182
rect	522	190	523	191
rect	522	193	523	194
rect	522	196	523	197
rect	522	199	523	200
rect	522	202	523	203
rect	522	208	523	209
rect	522	211	523	212
rect	522	214	523	215
rect	522	235	523	236
rect	522	238	523	239
rect	522	241	523	242
rect	522	247	523	248
rect	522	250	523	251
rect	522	274	523	275
rect	522	277	523	278
rect	523	7	524	8
rect	523	13	524	14
rect	523	25	524	26
rect	523	28	524	29
rect	523	31	524	32
rect	523	34	524	35
rect	523	37	524	38
rect	523	40	524	41
rect	523	43	524	44
rect	523	46	524	47
rect	523	49	524	50
rect	523	52	524	53
rect	523	61	524	62
rect	523	64	524	65
rect	523	67	524	68
rect	523	70	524	71
rect	523	73	524	74
rect	523	82	524	83
rect	523	85	524	86
rect	523	88	524	89
rect	523	91	524	92
rect	523	100	524	101
rect	523	115	524	116
rect	523	118	524	119
rect	523	121	524	122
rect	523	124	524	125
rect	523	130	524	131
rect	523	139	524	140
rect	523	148	524	149
rect	523	151	524	152
rect	523	160	524	161
rect	523	163	524	164
rect	523	166	524	167
rect	523	169	524	170
rect	523	175	524	176
rect	523	178	524	179
rect	523	181	524	182
rect	523	190	524	191
rect	523	193	524	194
rect	523	196	524	197
rect	523	199	524	200
rect	523	202	524	203
rect	523	208	524	209
rect	523	211	524	212
rect	523	214	524	215
rect	523	235	524	236
rect	523	238	524	239
rect	523	241	524	242
rect	523	247	524	248
rect	523	250	524	251
rect	523	253	524	254
rect	523	256	524	257
rect	523	265	524	266
rect	523	274	524	275
rect	523	277	524	278
rect	530	7	531	8
rect	530	10	531	11
rect	530	13	531	14
rect	530	25	531	26
rect	530	28	531	29
rect	530	31	531	32
rect	530	34	531	35
rect	530	37	531	38
rect	530	40	531	41
rect	530	43	531	44
rect	530	46	531	47
rect	530	49	531	50
rect	530	52	531	53
rect	530	55	531	56
rect	530	61	531	62
rect	530	64	531	65
rect	530	67	531	68
rect	530	70	531	71
rect	530	73	531	74
rect	530	82	531	83
rect	530	85	531	86
rect	530	88	531	89
rect	530	91	531	92
rect	530	100	531	101
rect	530	115	531	116
rect	530	118	531	119
rect	530	121	531	122
rect	530	124	531	125
rect	530	127	531	128
rect	530	139	531	140
rect	530	148	531	149
rect	530	151	531	152
rect	530	160	531	161
rect	530	163	531	164
rect	530	166	531	167
rect	530	175	531	176
rect	530	178	531	179
rect	530	181	531	182
rect	530	190	531	191
rect	530	193	531	194
rect	530	196	531	197
rect	530	199	531	200
rect	530	202	531	203
rect	530	208	531	209
rect	530	211	531	212
rect	530	214	531	215
rect	530	235	531	236
rect	530	238	531	239
rect	530	247	531	248
rect	530	256	531	257
rect	530	265	531	266
rect	530	274	531	275
rect	531	7	532	8
rect	531	10	532	11
rect	531	13	532	14
rect	531	25	532	26
rect	531	28	532	29
rect	531	31	532	32
rect	531	34	532	35
rect	531	37	532	38
rect	531	40	532	41
rect	531	43	532	44
rect	531	46	532	47
rect	531	49	532	50
rect	531	52	532	53
rect	531	55	532	56
rect	531	61	532	62
rect	531	64	532	65
rect	531	67	532	68
rect	531	70	532	71
rect	531	73	532	74
rect	531	82	532	83
rect	531	85	532	86
rect	531	88	532	89
rect	531	91	532	92
rect	531	100	532	101
rect	531	115	532	116
rect	531	118	532	119
rect	531	121	532	122
rect	531	124	532	125
rect	531	127	532	128
rect	531	139	532	140
rect	531	148	532	149
rect	531	151	532	152
rect	531	163	532	164
rect	531	166	532	167
rect	531	175	532	176
rect	531	178	532	179
rect	531	181	532	182
rect	531	190	532	191
rect	531	193	532	194
rect	531	196	532	197
rect	531	199	532	200
rect	531	202	532	203
rect	531	208	532	209
rect	531	211	532	212
rect	531	214	532	215
rect	531	235	532	236
rect	531	238	532	239
rect	531	247	532	248
rect	531	256	532	257
rect	531	265	532	266
rect	531	274	532	275
rect	532	7	533	8
rect	532	10	533	11
rect	532	13	533	14
rect	532	25	533	26
rect	532	28	533	29
rect	532	31	533	32
rect	532	34	533	35
rect	532	37	533	38
rect	532	40	533	41
rect	532	43	533	44
rect	532	46	533	47
rect	532	49	533	50
rect	532	52	533	53
rect	532	55	533	56
rect	532	61	533	62
rect	532	64	533	65
rect	532	67	533	68
rect	532	70	533	71
rect	532	73	533	74
rect	532	82	533	83
rect	532	85	533	86
rect	532	88	533	89
rect	532	91	533	92
rect	532	100	533	101
rect	532	115	533	116
rect	532	118	533	119
rect	532	121	533	122
rect	532	124	533	125
rect	532	127	533	128
rect	532	139	533	140
rect	532	148	533	149
rect	532	151	533	152
rect	532	154	533	155
rect	532	163	533	164
rect	532	166	533	167
rect	532	175	533	176
rect	532	178	533	179
rect	532	181	533	182
rect	532	190	533	191
rect	532	193	533	194
rect	532	196	533	197
rect	532	199	533	200
rect	532	202	533	203
rect	532	208	533	209
rect	532	211	533	212
rect	532	214	533	215
rect	532	235	533	236
rect	532	238	533	239
rect	532	247	533	248
rect	532	256	533	257
rect	532	265	533	266
rect	532	274	533	275
rect	533	7	534	8
rect	533	10	534	11
rect	533	13	534	14
rect	533	25	534	26
rect	533	28	534	29
rect	533	31	534	32
rect	533	34	534	35
rect	533	37	534	38
rect	533	40	534	41
rect	533	43	534	44
rect	533	46	534	47
rect	533	49	534	50
rect	533	52	534	53
rect	533	55	534	56
rect	533	61	534	62
rect	533	64	534	65
rect	533	67	534	68
rect	533	70	534	71
rect	533	73	534	74
rect	533	82	534	83
rect	533	85	534	86
rect	533	88	534	89
rect	533	91	534	92
rect	533	100	534	101
rect	533	115	534	116
rect	533	118	534	119
rect	533	121	534	122
rect	533	124	534	125
rect	533	127	534	128
rect	533	139	534	140
rect	533	148	534	149
rect	533	151	534	152
rect	533	154	534	155
rect	533	163	534	164
rect	533	175	534	176
rect	533	178	534	179
rect	533	181	534	182
rect	533	190	534	191
rect	533	193	534	194
rect	533	196	534	197
rect	533	199	534	200
rect	533	202	534	203
rect	533	208	534	209
rect	533	211	534	212
rect	533	214	534	215
rect	533	235	534	236
rect	533	238	534	239
rect	533	247	534	248
rect	533	256	534	257
rect	533	265	534	266
rect	533	274	534	275
rect	534	7	535	8
rect	534	10	535	11
rect	534	13	535	14
rect	534	25	535	26
rect	534	28	535	29
rect	534	31	535	32
rect	534	34	535	35
rect	534	37	535	38
rect	534	40	535	41
rect	534	43	535	44
rect	534	46	535	47
rect	534	49	535	50
rect	534	52	535	53
rect	534	55	535	56
rect	534	61	535	62
rect	534	64	535	65
rect	534	67	535	68
rect	534	70	535	71
rect	534	73	535	74
rect	534	82	535	83
rect	534	85	535	86
rect	534	88	535	89
rect	534	91	535	92
rect	534	100	535	101
rect	534	115	535	116
rect	534	118	535	119
rect	534	121	535	122
rect	534	124	535	125
rect	534	127	535	128
rect	534	139	535	140
rect	534	148	535	149
rect	534	151	535	152
rect	534	154	535	155
rect	534	160	535	161
rect	534	163	535	164
rect	534	175	535	176
rect	534	178	535	179
rect	534	181	535	182
rect	534	190	535	191
rect	534	193	535	194
rect	534	196	535	197
rect	534	199	535	200
rect	534	202	535	203
rect	534	208	535	209
rect	534	211	535	212
rect	534	214	535	215
rect	534	235	535	236
rect	534	238	535	239
rect	534	247	535	248
rect	534	256	535	257
rect	534	265	535	266
rect	534	274	535	275
rect	535	7	536	8
rect	535	10	536	11
rect	535	13	536	14
rect	535	34	536	35
rect	535	37	536	38
rect	535	40	536	41
rect	535	43	536	44
rect	535	46	536	47
rect	535	49	536	50
rect	535	52	536	53
rect	535	61	536	62
rect	535	64	536	65
rect	535	67	536	68
rect	535	70	536	71
rect	535	73	536	74
rect	535	82	536	83
rect	535	85	536	86
rect	535	88	536	89
rect	535	91	536	92
rect	535	100	536	101
rect	535	115	536	116
rect	535	118	536	119
rect	535	121	536	122
rect	535	124	536	125
rect	535	127	536	128
rect	535	139	536	140
rect	535	148	536	149
rect	535	151	536	152
rect	535	154	536	155
rect	535	160	536	161
rect	535	175	536	176
rect	535	178	536	179
rect	535	190	536	191
rect	535	193	536	194
rect	535	196	536	197
rect	535	199	536	200
rect	535	202	536	203
rect	535	208	536	209
rect	535	211	536	212
rect	535	214	536	215
rect	535	235	536	236
rect	535	238	536	239
rect	535	247	536	248
rect	535	256	536	257
rect	535	265	536	266
rect	535	274	536	275
rect	536	7	537	8
rect	536	10	537	11
rect	536	13	537	14
rect	536	34	537	35
rect	536	37	537	38
rect	536	40	537	41
rect	536	43	537	44
rect	536	46	537	47
rect	536	49	537	50
rect	536	52	537	53
rect	536	61	537	62
rect	536	64	537	65
rect	536	67	537	68
rect	536	70	537	71
rect	536	73	537	74
rect	536	82	537	83
rect	536	85	537	86
rect	536	88	537	89
rect	536	91	537	92
rect	536	100	537	101
rect	536	115	537	116
rect	536	118	537	119
rect	536	121	537	122
rect	536	124	537	125
rect	536	127	537	128
rect	536	139	537	140
rect	536	148	537	149
rect	536	151	537	152
rect	536	154	537	155
rect	536	157	537	158
rect	536	160	537	161
rect	536	166	537	167
rect	536	175	537	176
rect	536	178	537	179
rect	536	190	537	191
rect	536	193	537	194
rect	536	196	537	197
rect	536	199	537	200
rect	536	202	537	203
rect	536	208	537	209
rect	536	211	537	212
rect	536	214	537	215
rect	536	235	537	236
rect	536	238	537	239
rect	536	247	537	248
rect	536	256	537	257
rect	536	265	537	266
rect	536	274	537	275
rect	537	7	538	8
rect	537	10	538	11
rect	537	13	538	14
rect	537	34	538	35
rect	537	37	538	38
rect	537	40	538	41
rect	537	43	538	44
rect	537	46	538	47
rect	537	49	538	50
rect	537	61	538	62
rect	537	67	538	68
rect	537	70	538	71
rect	537	73	538	74
rect	537	82	538	83
rect	537	88	538	89
rect	537	91	538	92
rect	537	100	538	101
rect	537	115	538	116
rect	537	118	538	119
rect	537	121	538	122
rect	537	124	538	125
rect	537	127	538	128
rect	537	139	538	140
rect	537	148	538	149
rect	537	154	538	155
rect	537	157	538	158
rect	537	160	538	161
rect	537	166	538	167
rect	537	175	538	176
rect	537	190	538	191
rect	537	193	538	194
rect	537	196	538	197
rect	537	211	538	212
rect	537	214	538	215
rect	537	235	538	236
rect	537	238	538	239
rect	537	256	538	257
rect	537	265	538	266
rect	537	274	538	275
rect	538	7	539	8
rect	538	10	539	11
rect	538	13	539	14
rect	538	28	539	29
rect	538	34	539	35
rect	538	37	539	38
rect	538	40	539	41
rect	538	43	539	44
rect	538	46	539	47
rect	538	49	539	50
rect	538	55	539	56
rect	538	61	539	62
rect	538	67	539	68
rect	538	70	539	71
rect	538	73	539	74
rect	538	79	539	80
rect	538	82	539	83
rect	538	88	539	89
rect	538	91	539	92
rect	538	100	539	101
rect	538	115	539	116
rect	538	118	539	119
rect	538	121	539	122
rect	538	124	539	125
rect	538	127	539	128
rect	538	133	539	134
rect	538	139	539	140
rect	538	148	539	149
rect	538	154	539	155
rect	538	157	539	158
rect	538	160	539	161
rect	538	163	539	164
rect	538	166	539	167
rect	538	175	539	176
rect	538	184	539	185
rect	538	190	539	191
rect	538	193	539	194
rect	538	196	539	197
rect	538	211	539	212
rect	538	214	539	215
rect	538	232	539	233
rect	538	235	539	236
rect	538	238	539	239
rect	538	256	539	257
rect	538	265	539	266
rect	538	274	539	275
rect	539	7	540	8
rect	539	10	540	11
rect	539	13	540	14
rect	539	28	540	29
rect	539	34	540	35
rect	539	37	540	38
rect	539	40	540	41
rect	539	43	540	44
rect	539	46	540	47
rect	539	49	540	50
rect	539	55	540	56
rect	539	67	540	68
rect	539	70	540	71
rect	539	79	540	80
rect	539	82	540	83
rect	539	88	540	89
rect	539	91	540	92
rect	539	115	540	116
rect	539	118	540	119
rect	539	124	540	125
rect	539	127	540	128
rect	539	133	540	134
rect	539	139	540	140
rect	539	148	540	149
rect	539	154	540	155
rect	539	157	540	158
rect	539	160	540	161
rect	539	163	540	164
rect	539	166	540	167
rect	539	184	540	185
rect	539	190	540	191
rect	539	196	540	197
rect	539	214	540	215
rect	539	232	540	233
rect	539	235	540	236
rect	539	256	540	257
rect	539	265	540	266
rect	539	274	540	275
rect	540	7	541	8
rect	540	10	541	11
rect	540	13	541	14
rect	540	28	541	29
rect	540	34	541	35
rect	540	37	541	38
rect	540	40	541	41
rect	540	43	541	44
rect	540	46	541	47
rect	540	49	541	50
rect	540	52	541	53
rect	540	55	541	56
rect	540	64	541	65
rect	540	67	541	68
rect	540	70	541	71
rect	540	76	541	77
rect	540	79	541	80
rect	540	82	541	83
rect	540	88	541	89
rect	540	91	541	92
rect	540	112	541	113
rect	540	115	541	116
rect	540	118	541	119
rect	540	124	541	125
rect	540	127	541	128
rect	540	133	541	134
rect	540	139	541	140
rect	540	148	541	149
rect	540	151	541	152
rect	540	154	541	155
rect	540	157	541	158
rect	540	160	541	161
rect	540	163	541	164
rect	540	166	541	167
rect	540	178	541	179
rect	540	184	541	185
rect	540	190	541	191
rect	540	196	541	197
rect	540	202	541	203
rect	540	214	541	215
rect	540	229	541	230
rect	540	232	541	233
rect	540	235	541	236
rect	540	256	541	257
rect	540	265	541	266
rect	540	274	541	275
rect	541	7	542	8
rect	541	10	542	11
rect	541	13	542	14
rect	541	28	542	29
rect	541	34	542	35
rect	541	37	542	38
rect	541	40	542	41
rect	541	43	542	44
rect	541	46	542	47
rect	541	49	542	50
rect	541	52	542	53
rect	541	55	542	56
rect	541	64	542	65
rect	541	67	542	68
rect	541	76	542	77
rect	541	79	542	80
rect	541	88	542	89
rect	541	112	542	113
rect	541	115	542	116
rect	541	124	542	125
rect	541	133	542	134
rect	541	139	542	140
rect	541	148	542	149
rect	541	151	542	152
rect	541	154	542	155
rect	541	157	542	158
rect	541	160	542	161
rect	541	163	542	164
rect	541	166	542	167
rect	541	178	542	179
rect	541	184	542	185
rect	541	190	542	191
rect	541	196	542	197
rect	541	202	542	203
rect	541	214	542	215
rect	541	229	542	230
rect	541	232	542	233
rect	541	235	542	236
rect	541	256	542	257
rect	541	265	542	266
rect	541	274	542	275
rect	542	7	543	8
rect	542	10	543	11
rect	542	13	543	14
rect	542	28	543	29
rect	542	34	543	35
rect	542	37	543	38
rect	542	40	543	41
rect	542	43	543	44
rect	542	46	543	47
rect	542	49	543	50
rect	542	52	543	53
rect	542	55	543	56
rect	542	61	543	62
rect	542	64	543	65
rect	542	67	543	68
rect	542	73	543	74
rect	542	76	543	77
rect	542	79	543	80
rect	542	85	543	86
rect	542	88	543	89
rect	542	109	543	110
rect	542	112	543	113
rect	542	115	543	116
rect	542	124	543	125
rect	542	133	543	134
rect	542	139	543	140
rect	542	148	543	149
rect	542	151	543	152
rect	542	154	543	155
rect	542	157	543	158
rect	542	160	543	161
rect	542	163	543	164
rect	542	166	543	167
rect	542	178	543	179
rect	542	184	543	185
rect	542	190	543	191
rect	542	196	543	197
rect	542	202	543	203
rect	542	214	543	215
rect	542	229	543	230
rect	542	232	543	233
rect	542	235	543	236
rect	542	241	543	242
rect	542	256	543	257
rect	542	265	543	266
rect	542	274	543	275
rect	543	7	544	8
rect	543	13	544	14
rect	543	28	544	29
rect	543	34	544	35
rect	543	37	544	38
rect	543	40	544	41
rect	543	43	544	44
rect	543	46	544	47
rect	543	49	544	50
rect	543	52	544	53
rect	543	55	544	56
rect	543	61	544	62
rect	543	64	544	65
rect	543	67	544	68
rect	543	73	544	74
rect	543	76	544	77
rect	543	79	544	80
rect	543	85	544	86
rect	543	88	544	89
rect	543	109	544	110
rect	543	112	544	113
rect	543	115	544	116
rect	543	124	544	125
rect	543	133	544	134
rect	543	139	544	140
rect	543	148	544	149
rect	543	151	544	152
rect	543	154	544	155
rect	543	157	544	158
rect	543	160	544	161
rect	543	163	544	164
rect	543	166	544	167
rect	543	178	544	179
rect	543	184	544	185
rect	543	190	544	191
rect	543	202	544	203
rect	543	229	544	230
rect	543	232	544	233
rect	543	241	544	242
rect	543	265	544	266
rect	544	7	545	8
rect	544	13	545	14
rect	544	28	545	29
rect	544	34	545	35
rect	544	37	545	38
rect	544	40	545	41
rect	544	43	545	44
rect	544	46	545	47
rect	544	49	545	50
rect	544	52	545	53
rect	544	55	545	56
rect	544	61	545	62
rect	544	64	545	65
rect	544	67	545	68
rect	544	73	545	74
rect	544	76	545	77
rect	544	79	545	80
rect	544	85	545	86
rect	544	88	545	89
rect	544	109	545	110
rect	544	112	545	113
rect	544	115	545	116
rect	544	124	545	125
rect	544	133	545	134
rect	544	139	545	140
rect	544	148	545	149
rect	544	151	545	152
rect	544	154	545	155
rect	544	157	545	158
rect	544	160	545	161
rect	544	163	545	164
rect	544	166	545	167
rect	544	178	545	179
rect	544	181	545	182
rect	544	184	545	185
rect	544	190	545	191
rect	544	199	545	200
rect	544	202	545	203
rect	544	211	545	212
rect	544	220	545	221
rect	544	229	545	230
rect	544	232	545	233
rect	544	241	545	242
rect	544	247	545	248
rect	544	259	545	260
rect	544	265	545	266
rect	545	28	546	29
rect	545	37	546	38
rect	545	40	546	41
rect	545	43	546	44
rect	545	46	546	47
rect	545	49	546	50
rect	545	52	546	53
rect	545	55	546	56
rect	545	61	546	62
rect	545	64	546	65
rect	545	73	546	74
rect	545	76	546	77
rect	545	79	546	80
rect	545	85	546	86
rect	545	109	546	110
rect	545	112	546	113
rect	545	124	546	125
rect	545	133	546	134
rect	545	151	546	152
rect	545	154	546	155
rect	545	157	546	158
rect	545	160	546	161
rect	545	163	546	164
rect	545	166	546	167
rect	545	178	546	179
rect	545	181	546	182
rect	545	184	546	185
rect	545	199	546	200
rect	545	202	546	203
rect	545	211	546	212
rect	545	220	546	221
rect	545	229	546	230
rect	545	232	546	233
rect	545	241	546	242
rect	545	247	546	248
rect	545	259	546	260
rect	546	25	547	26
rect	546	28	547	29
rect	546	37	547	38
rect	546	40	547	41
rect	546	43	547	44
rect	546	46	547	47
rect	546	49	547	50
rect	546	52	547	53
rect	546	55	547	56
rect	546	58	547	59
rect	546	61	547	62
rect	546	64	547	65
rect	546	73	547	74
rect	546	76	547	77
rect	546	79	547	80
rect	546	82	547	83
rect	546	85	547	86
rect	546	100	547	101
rect	546	109	547	110
rect	546	112	547	113
rect	546	121	547	122
rect	546	124	547	125
rect	546	133	547	134
rect	546	142	547	143
rect	546	151	547	152
rect	546	154	547	155
rect	546	157	547	158
rect	546	160	547	161
rect	546	163	547	164
rect	546	166	547	167
rect	546	175	547	176
rect	546	178	547	179
rect	546	181	547	182
rect	546	184	547	185
rect	546	196	547	197
rect	546	199	547	200
rect	546	202	547	203
rect	546	211	547	212
rect	546	220	547	221
rect	546	229	547	230
rect	546	232	547	233
rect	546	241	547	242
rect	546	244	547	245
rect	546	247	547	248
rect	546	256	547	257
rect	546	259	547	260
rect	553	22	554	23
rect	553	25	554	26
rect	553	28	554	29
rect	553	31	554	32
rect	553	37	554	38
rect	553	40	554	41
rect	553	43	554	44
rect	553	46	554	47
rect	553	49	554	50
rect	553	52	554	53
rect	553	55	554	56
rect	553	58	554	59
rect	553	61	554	62
rect	553	64	554	65
rect	553	73	554	74
rect	553	76	554	77
rect	553	79	554	80
rect	553	82	554	83
rect	553	85	554	86
rect	553	100	554	101
rect	553	109	554	110
rect	553	112	554	113
rect	553	118	554	119
rect	553	121	554	122
rect	553	124	554	125
rect	553	133	554	134
rect	553	142	554	143
rect	553	151	554	152
rect	553	154	554	155
rect	553	157	554	158
rect	553	160	554	161
rect	553	163	554	164
rect	553	166	554	167
rect	553	169	554	170
rect	553	172	554	173
rect	553	175	554	176
rect	553	178	554	179
rect	553	181	554	182
rect	553	184	554	185
rect	553	196	554	197
rect	553	199	554	200
rect	553	202	554	203
rect	553	211	554	212
rect	553	220	554	221
rect	553	229	554	230
rect	553	232	554	233
rect	553	235	554	236
rect	553	241	554	242
rect	553	244	554	245
rect	553	247	554	248
rect	553	250	554	251
rect	553	256	554	257
rect	553	259	554	260
rect	554	22	555	23
rect	554	25	555	26
rect	554	28	555	29
rect	554	31	555	32
rect	554	37	555	38
rect	554	40	555	41
rect	554	43	555	44
rect	554	49	555	50
rect	554	52	555	53
rect	554	55	555	56
rect	554	58	555	59
rect	554	61	555	62
rect	554	64	555	65
rect	554	73	555	74
rect	554	76	555	77
rect	554	79	555	80
rect	554	82	555	83
rect	554	85	555	86
rect	554	100	555	101
rect	554	109	555	110
rect	554	112	555	113
rect	554	118	555	119
rect	554	121	555	122
rect	554	124	555	125
rect	554	133	555	134
rect	554	142	555	143
rect	554	154	555	155
rect	554	157	555	158
rect	554	160	555	161
rect	554	163	555	164
rect	554	166	555	167
rect	554	172	555	173
rect	554	175	555	176
rect	554	178	555	179
rect	554	181	555	182
rect	554	184	555	185
rect	554	196	555	197
rect	554	199	555	200
rect	554	202	555	203
rect	554	211	555	212
rect	554	220	555	221
rect	554	229	555	230
rect	554	232	555	233
rect	554	235	555	236
rect	554	241	555	242
rect	554	244	555	245
rect	554	247	555	248
rect	554	250	555	251
rect	554	256	555	257
rect	554	259	555	260
rect	555	22	556	23
rect	555	25	556	26
rect	555	28	556	29
rect	555	31	556	32
rect	555	34	556	35
rect	555	37	556	38
rect	555	40	556	41
rect	555	43	556	44
rect	555	49	556	50
rect	555	52	556	53
rect	555	55	556	56
rect	555	58	556	59
rect	555	61	556	62
rect	555	64	556	65
rect	555	73	556	74
rect	555	76	556	77
rect	555	79	556	80
rect	555	82	556	83
rect	555	85	556	86
rect	555	100	556	101
rect	555	109	556	110
rect	555	112	556	113
rect	555	118	556	119
rect	555	121	556	122
rect	555	124	556	125
rect	555	133	556	134
rect	555	142	556	143
rect	555	154	556	155
rect	555	157	556	158
rect	555	160	556	161
rect	555	163	556	164
rect	555	166	556	167
rect	555	172	556	173
rect	555	175	556	176
rect	555	178	556	179
rect	555	181	556	182
rect	555	184	556	185
rect	555	196	556	197
rect	555	199	556	200
rect	555	202	556	203
rect	555	211	556	212
rect	555	220	556	221
rect	555	229	556	230
rect	555	232	556	233
rect	555	235	556	236
rect	555	241	556	242
rect	555	244	556	245
rect	555	247	556	248
rect	555	250	556	251
rect	555	256	556	257
rect	555	259	556	260
rect	556	22	557	23
rect	556	25	557	26
rect	556	28	557	29
rect	556	34	557	35
rect	556	40	557	41
rect	556	43	557	44
rect	556	49	557	50
rect	556	52	557	53
rect	556	58	557	59
rect	556	61	557	62
rect	556	64	557	65
rect	556	73	557	74
rect	556	76	557	77
rect	556	79	557	80
rect	556	82	557	83
rect	556	85	557	86
rect	556	100	557	101
rect	556	109	557	110
rect	556	112	557	113
rect	556	118	557	119
rect	556	121	557	122
rect	556	124	557	125
rect	556	133	557	134
rect	556	142	557	143
rect	556	154	557	155
rect	556	157	557	158
rect	556	160	557	161
rect	556	163	557	164
rect	556	172	557	173
rect	556	175	557	176
rect	556	178	557	179
rect	556	181	557	182
rect	556	184	557	185
rect	556	196	557	197
rect	556	199	557	200
rect	556	202	557	203
rect	556	211	557	212
rect	556	220	557	221
rect	556	229	557	230
rect	556	232	557	233
rect	556	235	557	236
rect	556	241	557	242
rect	556	244	557	245
rect	556	247	557	248
rect	556	250	557	251
rect	556	256	557	257
rect	556	259	557	260
rect	557	22	558	23
rect	557	25	558	26
rect	557	28	558	29
rect	557	34	558	35
rect	557	40	558	41
rect	557	43	558	44
rect	557	49	558	50
rect	557	52	558	53
rect	557	58	558	59
rect	557	61	558	62
rect	557	64	558	65
rect	557	70	558	71
rect	557	73	558	74
rect	557	76	558	77
rect	557	79	558	80
rect	557	82	558	83
rect	557	85	558	86
rect	557	100	558	101
rect	557	109	558	110
rect	557	112	558	113
rect	557	118	558	119
rect	557	121	558	122
rect	557	124	558	125
rect	557	133	558	134
rect	557	142	558	143
rect	557	154	558	155
rect	557	157	558	158
rect	557	160	558	161
rect	557	163	558	164
rect	557	169	558	170
rect	557	172	558	173
rect	557	175	558	176
rect	557	178	558	179
rect	557	181	558	182
rect	557	184	558	185
rect	557	196	558	197
rect	557	199	558	200
rect	557	202	558	203
rect	557	211	558	212
rect	557	220	558	221
rect	557	229	558	230
rect	557	232	558	233
rect	557	235	558	236
rect	557	241	558	242
rect	557	244	558	245
rect	557	247	558	248
rect	557	250	558	251
rect	557	256	558	257
rect	557	259	558	260
rect	558	22	559	23
rect	558	25	559	26
rect	558	28	559	29
rect	558	34	559	35
rect	558	40	559	41
rect	558	49	559	50
rect	558	52	559	53
rect	558	58	559	59
rect	558	61	559	62
rect	558	70	559	71
rect	558	73	559	74
rect	558	76	559	77
rect	558	79	559	80
rect	558	82	559	83
rect	558	85	559	86
rect	558	100	559	101
rect	558	109	559	110
rect	558	112	559	113
rect	558	118	559	119
rect	558	121	559	122
rect	558	124	559	125
rect	558	133	559	134
rect	558	142	559	143
rect	558	154	559	155
rect	558	157	559	158
rect	558	160	559	161
rect	558	169	559	170
rect	558	172	559	173
rect	558	175	559	176
rect	558	178	559	179
rect	558	181	559	182
rect	558	184	559	185
rect	558	196	559	197
rect	558	199	559	200
rect	558	202	559	203
rect	558	211	559	212
rect	558	220	559	221
rect	558	229	559	230
rect	558	232	559	233
rect	558	235	559	236
rect	558	241	559	242
rect	558	244	559	245
rect	558	247	559	248
rect	558	250	559	251
rect	558	256	559	257
rect	558	259	559	260
rect	559	22	560	23
rect	559	25	560	26
rect	559	28	560	29
rect	559	31	560	32
rect	559	34	560	35
rect	559	40	560	41
rect	559	49	560	50
rect	559	52	560	53
rect	559	55	560	56
rect	559	58	560	59
rect	559	61	560	62
rect	559	70	560	71
rect	559	73	560	74
rect	559	76	560	77
rect	559	79	560	80
rect	559	82	560	83
rect	559	85	560	86
rect	559	100	560	101
rect	559	109	560	110
rect	559	112	560	113
rect	559	118	560	119
rect	559	121	560	122
rect	559	124	560	125
rect	559	133	560	134
rect	559	142	560	143
rect	559	154	560	155
rect	559	157	560	158
rect	559	160	560	161
rect	559	166	560	167
rect	559	169	560	170
rect	559	172	560	173
rect	559	175	560	176
rect	559	178	560	179
rect	559	181	560	182
rect	559	184	560	185
rect	559	196	560	197
rect	559	199	560	200
rect	559	202	560	203
rect	559	211	560	212
rect	559	220	560	221
rect	559	229	560	230
rect	559	232	560	233
rect	559	235	560	236
rect	559	241	560	242
rect	559	244	560	245
rect	559	247	560	248
rect	559	250	560	251
rect	559	256	560	257
rect	559	259	560	260
rect	560	22	561	23
rect	560	25	561	26
rect	560	31	561	32
rect	560	34	561	35
rect	560	40	561	41
rect	560	49	561	50
rect	560	52	561	53
rect	560	55	561	56
rect	560	58	561	59
rect	560	61	561	62
rect	560	70	561	71
rect	560	76	561	77
rect	560	79	561	80
rect	560	82	561	83
rect	560	85	561	86
rect	560	100	561	101
rect	560	109	561	110
rect	560	112	561	113
rect	560	118	561	119
rect	560	121	561	122
rect	560	124	561	125
rect	560	133	561	134
rect	560	142	561	143
rect	560	154	561	155
rect	560	160	561	161
rect	560	166	561	167
rect	560	169	561	170
rect	560	172	561	173
rect	560	175	561	176
rect	560	178	561	179
rect	560	181	561	182
rect	560	196	561	197
rect	560	202	561	203
rect	560	211	561	212
rect	560	220	561	221
rect	560	229	561	230
rect	560	232	561	233
rect	560	235	561	236
rect	560	241	561	242
rect	560	244	561	245
rect	560	247	561	248
rect	560	250	561	251
rect	560	256	561	257
rect	560	259	561	260
rect	561	22	562	23
rect	561	25	562	26
rect	561	31	562	32
rect	561	34	562	35
rect	561	40	562	41
rect	561	43	562	44
rect	561	49	562	50
rect	561	52	562	53
rect	561	55	562	56
rect	561	58	562	59
rect	561	61	562	62
rect	561	64	562	65
rect	561	70	562	71
rect	561	76	562	77
rect	561	79	562	80
rect	561	82	562	83
rect	561	85	562	86
rect	561	100	562	101
rect	561	109	562	110
rect	561	112	562	113
rect	561	118	562	119
rect	561	121	562	122
rect	561	124	562	125
rect	561	133	562	134
rect	561	142	562	143
rect	561	148	562	149
rect	561	154	562	155
rect	561	160	562	161
rect	561	163	562	164
rect	561	166	562	167
rect	561	169	562	170
rect	561	172	562	173
rect	561	175	562	176
rect	561	178	562	179
rect	561	181	562	182
rect	561	196	562	197
rect	561	202	562	203
rect	561	205	562	206
rect	561	211	562	212
rect	561	220	562	221
rect	561	229	562	230
rect	561	232	562	233
rect	561	235	562	236
rect	561	241	562	242
rect	561	244	562	245
rect	561	247	562	248
rect	561	250	562	251
rect	561	256	562	257
rect	561	259	562	260
rect	562	22	563	23
rect	562	25	563	26
rect	562	31	563	32
rect	562	34	563	35
rect	562	43	563	44
rect	562	49	563	50
rect	562	52	563	53
rect	562	55	563	56
rect	562	58	563	59
rect	562	61	563	62
rect	562	64	563	65
rect	562	70	563	71
rect	562	76	563	77
rect	562	79	563	80
rect	562	82	563	83
rect	562	85	563	86
rect	562	100	563	101
rect	562	109	563	110
rect	562	112	563	113
rect	562	118	563	119
rect	562	121	563	122
rect	562	124	563	125
rect	562	133	563	134
rect	562	142	563	143
rect	562	148	563	149
rect	562	154	563	155
rect	562	160	563	161
rect	562	163	563	164
rect	562	166	563	167
rect	562	169	563	170
rect	562	172	563	173
rect	562	175	563	176
rect	562	178	563	179
rect	562	181	563	182
rect	562	196	563	197
rect	562	202	563	203
rect	562	205	563	206
rect	562	211	563	212
rect	562	220	563	221
rect	562	229	563	230
rect	562	232	563	233
rect	562	244	563	245
rect	562	247	563	248
rect	562	256	563	257
rect	562	259	563	260
rect	563	22	564	23
rect	563	25	564	26
rect	563	28	564	29
rect	563	31	564	32
rect	563	34	564	35
rect	563	43	564	44
rect	563	46	564	47
rect	563	49	564	50
rect	563	52	564	53
rect	563	55	564	56
rect	563	58	564	59
rect	563	61	564	62
rect	563	64	564	65
rect	563	70	564	71
rect	563	76	564	77
rect	563	79	564	80
rect	563	82	564	83
rect	563	85	564	86
rect	563	100	564	101
rect	563	109	564	110
rect	563	112	564	113
rect	563	118	564	119
rect	563	121	564	122
rect	563	124	564	125
rect	563	133	564	134
rect	563	142	564	143
rect	563	148	564	149
rect	563	154	564	155
rect	563	160	564	161
rect	563	163	564	164
rect	563	166	564	167
rect	563	169	564	170
rect	563	172	564	173
rect	563	175	564	176
rect	563	178	564	179
rect	563	181	564	182
rect	563	196	564	197
rect	563	202	564	203
rect	563	205	564	206
rect	563	211	564	212
rect	563	220	564	221
rect	563	229	564	230
rect	563	232	564	233
rect	563	244	564	245
rect	563	247	564	248
rect	563	256	564	257
rect	563	259	564	260
rect	564	22	565	23
rect	564	25	565	26
rect	564	28	565	29
rect	564	31	565	32
rect	564	34	565	35
rect	564	43	565	44
rect	564	46	565	47
rect	564	49	565	50
rect	564	55	565	56
rect	564	58	565	59
rect	564	61	565	62
rect	564	64	565	65
rect	564	70	565	71
rect	564	76	565	77
rect	564	82	565	83
rect	564	85	565	86
rect	564	100	565	101
rect	564	109	565	110
rect	564	112	565	113
rect	564	118	565	119
rect	564	121	565	122
rect	564	124	565	125
rect	564	133	565	134
rect	564	142	565	143
rect	564	148	565	149
rect	564	154	565	155
rect	564	160	565	161
rect	564	163	565	164
rect	564	166	565	167
rect	564	169	565	170
rect	564	172	565	173
rect	564	175	565	176
rect	564	181	565	182
rect	564	202	565	203
rect	564	205	565	206
rect	564	220	565	221
rect	564	232	565	233
rect	564	244	565	245
rect	564	256	565	257
rect	564	259	565	260
rect	565	22	566	23
rect	565	25	566	26
rect	565	28	566	29
rect	565	31	566	32
rect	565	34	566	35
rect	565	40	566	41
rect	565	43	566	44
rect	565	46	566	47
rect	565	49	566	50
rect	565	55	566	56
rect	565	58	566	59
rect	565	61	566	62
rect	565	64	566	65
rect	565	70	566	71
rect	565	73	566	74
rect	565	76	566	77
rect	565	82	566	83
rect	565	85	566	86
rect	565	100	566	101
rect	565	109	566	110
rect	565	112	566	113
rect	565	118	566	119
rect	565	121	566	122
rect	565	124	566	125
rect	565	133	566	134
rect	565	142	566	143
rect	565	148	566	149
rect	565	154	566	155
rect	565	157	566	158
rect	565	160	566	161
rect	565	163	566	164
rect	565	166	566	167
rect	565	169	566	170
rect	565	172	566	173
rect	565	175	566	176
rect	565	181	566	182
rect	565	202	566	203
rect	565	205	566	206
rect	565	217	566	218
rect	565	220	566	221
rect	565	232	566	233
rect	565	244	566	245
rect	565	250	566	251
rect	565	256	566	257
rect	565	259	566	260
rect	566	22	567	23
rect	566	25	567	26
rect	566	28	567	29
rect	566	31	567	32
rect	566	34	567	35
rect	566	40	567	41
rect	566	43	567	44
rect	566	46	567	47
rect	566	55	567	56
rect	566	58	567	59
rect	566	64	567	65
rect	566	70	567	71
rect	566	73	567	74
rect	566	82	567	83
rect	566	100	567	101
rect	566	109	567	110
rect	566	124	567	125
rect	566	133	567	134
rect	566	142	567	143
rect	566	148	567	149
rect	566	157	567	158
rect	566	160	567	161
rect	566	163	567	164
rect	566	166	567	167
rect	566	169	567	170
rect	566	175	567	176
rect	566	181	567	182
rect	566	205	567	206
rect	566	217	567	218
rect	566	220	567	221
rect	566	232	567	233
rect	566	250	567	251
rect	566	256	567	257
rect	567	22	568	23
rect	567	25	568	26
rect	567	28	568	29
rect	567	31	568	32
rect	567	34	568	35
rect	567	37	568	38
rect	567	40	568	41
rect	567	43	568	44
rect	567	46	568	47
rect	567	52	568	53
rect	567	55	568	56
rect	567	58	568	59
rect	567	64	568	65
rect	567	67	568	68
rect	567	70	568	71
rect	567	73	568	74
rect	567	79	568	80
rect	567	82	568	83
rect	567	100	568	101
rect	567	106	568	107
rect	567	109	568	110
rect	567	124	568	125
rect	567	133	568	134
rect	567	142	568	143
rect	567	148	568	149
rect	567	157	568	158
rect	567	160	568	161
rect	567	163	568	164
rect	567	166	568	167
rect	567	169	568	170
rect	567	175	568	176
rect	567	181	568	182
rect	567	196	568	197
rect	567	205	568	206
rect	567	214	568	215
rect	567	217	568	218
rect	567	220	568	221
rect	567	223	568	224
rect	567	229	568	230
rect	567	232	568	233
rect	567	247	568	248
rect	567	250	568	251
rect	567	256	568	257
rect	568	28	569	29
rect	568	31	569	32
rect	568	34	569	35
rect	568	37	569	38
rect	568	40	569	41
rect	568	43	569	44
rect	568	46	569	47
rect	568	52	569	53
rect	568	55	569	56
rect	568	64	569	65
rect	568	67	569	68
rect	568	70	569	71
rect	568	73	569	74
rect	568	79	569	80
rect	568	106	569	107
rect	568	124	569	125
rect	568	148	569	149
rect	568	157	569	158
rect	568	160	569	161
rect	568	163	569	164
rect	568	166	569	167
rect	568	169	569	170
rect	568	196	569	197
rect	568	205	569	206
rect	568	214	569	215
rect	568	217	569	218
rect	568	223	569	224
rect	568	229	569	230
rect	568	247	569	248
rect	568	250	569	251
rect	569	7	570	8
rect	569	13	570	14
rect	569	28	570	29
rect	569	31	570	32
rect	569	34	570	35
rect	569	37	570	38
rect	569	40	570	41
rect	569	43	570	44
rect	569	46	570	47
rect	569	49	570	50
rect	569	52	570	53
rect	569	55	570	56
rect	569	64	570	65
rect	569	67	570	68
rect	569	70	570	71
rect	569	73	570	74
rect	569	76	570	77
rect	569	79	570	80
rect	569	94	570	95
rect	569	103	570	104
rect	569	106	570	107
rect	569	115	570	116
rect	569	124	570	125
rect	569	145	570	146
rect	569	148	570	149
rect	569	154	570	155
rect	569	157	570	158
rect	569	160	570	161
rect	569	163	570	164
rect	569	166	570	167
rect	569	169	570	170
rect	569	184	570	185
rect	569	193	570	194
rect	569	196	570	197
rect	569	205	570	206
rect	569	214	570	215
rect	569	217	570	218
rect	569	223	570	224
rect	569	226	570	227
rect	569	229	570	230
rect	569	235	570	236
rect	569	238	570	239
rect	569	244	570	245
rect	569	247	570	248
rect	569	250	570	251
rect	576	13	577	14
rect	576	22	577	23
rect	576	28	577	29
rect	576	31	577	32
rect	576	34	577	35
rect	576	37	577	38
rect	576	40	577	41
rect	576	43	577	44
rect	576	46	577	47
rect	576	49	577	50
rect	576	52	577	53
rect	576	55	577	56
rect	576	61	577	62
rect	576	64	577	65
rect	576	67	577	68
rect	576	70	577	71
rect	576	73	577	74
rect	576	76	577	77
rect	576	79	577	80
rect	576	94	577	95
rect	576	103	577	104
rect	576	106	577	107
rect	576	115	577	116
rect	576	118	577	119
rect	576	124	577	125
rect	576	145	577	146
rect	576	151	577	152
rect	576	154	577	155
rect	576	157	577	158
rect	576	160	577	161
rect	576	163	577	164
rect	576	166	577	167
rect	576	169	577	170
rect	576	184	577	185
rect	576	193	577	194
rect	576	196	577	197
rect	576	205	577	206
rect	576	214	577	215
rect	576	217	577	218
rect	576	226	577	227
rect	576	229	577	230
rect	576	238	577	239
rect	576	247	577	248
rect	576	250	577	251
rect	576	256	577	257
rect	577	13	578	14
rect	577	31	578	32
rect	577	34	578	35
rect	577	37	578	38
rect	577	40	578	41
rect	577	43	578	44
rect	577	46	578	47
rect	577	49	578	50
rect	577	52	578	53
rect	577	55	578	56
rect	577	61	578	62
rect	577	64	578	65
rect	577	67	578	68
rect	577	70	578	71
rect	577	73	578	74
rect	577	76	578	77
rect	577	79	578	80
rect	577	94	578	95
rect	577	103	578	104
rect	577	106	578	107
rect	577	115	578	116
rect	577	118	578	119
rect	577	124	578	125
rect	577	145	578	146
rect	577	151	578	152
rect	577	154	578	155
rect	577	157	578	158
rect	577	160	578	161
rect	577	163	578	164
rect	577	166	578	167
rect	577	169	578	170
rect	577	184	578	185
rect	577	193	578	194
rect	577	196	578	197
rect	577	205	578	206
rect	577	214	578	215
rect	577	217	578	218
rect	577	226	578	227
rect	577	229	578	230
rect	577	238	578	239
rect	577	247	578	248
rect	577	250	578	251
rect	577	256	578	257
rect	578	13	579	14
rect	578	31	579	32
rect	578	34	579	35
rect	578	37	579	38
rect	578	40	579	41
rect	578	43	579	44
rect	578	46	579	47
rect	578	49	579	50
rect	578	52	579	53
rect	578	55	579	56
rect	578	61	579	62
rect	578	64	579	65
rect	578	67	579	68
rect	578	70	579	71
rect	578	73	579	74
rect	578	76	579	77
rect	578	79	579	80
rect	578	94	579	95
rect	578	103	579	104
rect	578	106	579	107
rect	578	115	579	116
rect	578	118	579	119
rect	578	124	579	125
rect	578	145	579	146
rect	578	151	579	152
rect	578	154	579	155
rect	578	157	579	158
rect	578	160	579	161
rect	578	163	579	164
rect	578	166	579	167
rect	578	169	579	170
rect	578	184	579	185
rect	578	193	579	194
rect	578	196	579	197
rect	578	205	579	206
rect	578	214	579	215
rect	578	217	579	218
rect	578	226	579	227
rect	578	229	579	230
rect	578	238	579	239
rect	578	247	579	248
rect	578	250	579	251
rect	578	256	579	257
rect	579	13	580	14
rect	579	31	580	32
rect	579	34	580	35
rect	579	37	580	38
rect	579	43	580	44
rect	579	46	580	47
rect	579	49	580	50
rect	579	52	580	53
rect	579	55	580	56
rect	579	61	580	62
rect	579	64	580	65
rect	579	67	580	68
rect	579	70	580	71
rect	579	73	580	74
rect	579	76	580	77
rect	579	79	580	80
rect	579	94	580	95
rect	579	103	580	104
rect	579	106	580	107
rect	579	115	580	116
rect	579	118	580	119
rect	579	124	580	125
rect	579	145	580	146
rect	579	151	580	152
rect	579	154	580	155
rect	579	157	580	158
rect	579	160	580	161
rect	579	163	580	164
rect	579	166	580	167
rect	579	169	580	170
rect	579	184	580	185
rect	579	193	580	194
rect	579	196	580	197
rect	579	205	580	206
rect	579	214	580	215
rect	579	217	580	218
rect	579	226	580	227
rect	579	229	580	230
rect	579	238	580	239
rect	579	247	580	248
rect	579	250	580	251
rect	579	256	580	257
rect	580	13	581	14
rect	580	22	581	23
rect	580	31	581	32
rect	580	34	581	35
rect	580	37	581	38
rect	580	43	581	44
rect	580	46	581	47
rect	580	49	581	50
rect	580	52	581	53
rect	580	55	581	56
rect	580	61	581	62
rect	580	64	581	65
rect	580	67	581	68
rect	580	70	581	71
rect	580	73	581	74
rect	580	76	581	77
rect	580	79	581	80
rect	580	94	581	95
rect	580	103	581	104
rect	580	106	581	107
rect	580	115	581	116
rect	580	118	581	119
rect	580	124	581	125
rect	580	145	581	146
rect	580	151	581	152
rect	580	154	581	155
rect	580	157	581	158
rect	580	160	581	161
rect	580	163	581	164
rect	580	166	581	167
rect	580	169	581	170
rect	580	184	581	185
rect	580	193	581	194
rect	580	196	581	197
rect	580	205	581	206
rect	580	214	581	215
rect	580	217	581	218
rect	580	226	581	227
rect	580	229	581	230
rect	580	238	581	239
rect	580	247	581	248
rect	580	250	581	251
rect	580	256	581	257
rect	581	13	582	14
rect	581	22	582	23
rect	581	31	582	32
rect	581	34	582	35
rect	581	43	582	44
rect	581	46	582	47
rect	581	49	582	50
rect	581	52	582	53
rect	581	55	582	56
rect	581	61	582	62
rect	581	64	582	65
rect	581	67	582	68
rect	581	70	582	71
rect	581	73	582	74
rect	581	76	582	77
rect	581	79	582	80
rect	581	94	582	95
rect	581	103	582	104
rect	581	106	582	107
rect	581	115	582	116
rect	581	118	582	119
rect	581	124	582	125
rect	581	145	582	146
rect	581	151	582	152
rect	581	154	582	155
rect	581	157	582	158
rect	581	160	582	161
rect	581	163	582	164
rect	581	166	582	167
rect	581	169	582	170
rect	581	184	582	185
rect	581	193	582	194
rect	581	196	582	197
rect	581	205	582	206
rect	581	214	582	215
rect	581	217	582	218
rect	581	226	582	227
rect	581	229	582	230
rect	581	238	582	239
rect	581	247	582	248
rect	581	250	582	251
rect	581	256	582	257
rect	582	13	583	14
rect	582	22	583	23
rect	582	31	583	32
rect	582	34	583	35
rect	582	40	583	41
rect	582	43	583	44
rect	582	46	583	47
rect	582	49	583	50
rect	582	52	583	53
rect	582	55	583	56
rect	582	61	583	62
rect	582	64	583	65
rect	582	67	583	68
rect	582	70	583	71
rect	582	73	583	74
rect	582	76	583	77
rect	582	79	583	80
rect	582	94	583	95
rect	582	103	583	104
rect	582	106	583	107
rect	582	115	583	116
rect	582	118	583	119
rect	582	124	583	125
rect	582	145	583	146
rect	582	151	583	152
rect	582	154	583	155
rect	582	157	583	158
rect	582	160	583	161
rect	582	163	583	164
rect	582	166	583	167
rect	582	169	583	170
rect	582	184	583	185
rect	582	193	583	194
rect	582	196	583	197
rect	582	205	583	206
rect	582	214	583	215
rect	582	217	583	218
rect	582	226	583	227
rect	582	229	583	230
rect	582	238	583	239
rect	582	247	583	248
rect	582	250	583	251
rect	582	256	583	257
rect	583	13	584	14
rect	583	22	584	23
rect	583	34	584	35
rect	583	40	584	41
rect	583	43	584	44
rect	583	46	584	47
rect	583	49	584	50
rect	583	52	584	53
rect	583	55	584	56
rect	583	61	584	62
rect	583	64	584	65
rect	583	67	584	68
rect	583	70	584	71
rect	583	73	584	74
rect	583	76	584	77
rect	583	79	584	80
rect	583	94	584	95
rect	583	103	584	104
rect	583	106	584	107
rect	583	115	584	116
rect	583	118	584	119
rect	583	124	584	125
rect	583	145	584	146
rect	583	151	584	152
rect	583	154	584	155
rect	583	157	584	158
rect	583	160	584	161
rect	583	163	584	164
rect	583	166	584	167
rect	583	169	584	170
rect	583	184	584	185
rect	583	193	584	194
rect	583	196	584	197
rect	583	205	584	206
rect	583	214	584	215
rect	583	217	584	218
rect	583	226	584	227
rect	583	229	584	230
rect	583	238	584	239
rect	583	247	584	248
rect	583	250	584	251
rect	583	256	584	257
rect	584	13	585	14
rect	584	22	585	23
rect	584	34	585	35
rect	584	37	585	38
rect	584	40	585	41
rect	584	43	585	44
rect	584	46	585	47
rect	584	49	585	50
rect	584	52	585	53
rect	584	55	585	56
rect	584	61	585	62
rect	584	64	585	65
rect	584	67	585	68
rect	584	70	585	71
rect	584	73	585	74
rect	584	76	585	77
rect	584	79	585	80
rect	584	94	585	95
rect	584	103	585	104
rect	584	106	585	107
rect	584	115	585	116
rect	584	118	585	119
rect	584	124	585	125
rect	584	145	585	146
rect	584	151	585	152
rect	584	154	585	155
rect	584	157	585	158
rect	584	160	585	161
rect	584	163	585	164
rect	584	166	585	167
rect	584	169	585	170
rect	584	184	585	185
rect	584	193	585	194
rect	584	196	585	197
rect	584	205	585	206
rect	584	214	585	215
rect	584	217	585	218
rect	584	226	585	227
rect	584	229	585	230
rect	584	238	585	239
rect	584	247	585	248
rect	584	250	585	251
rect	584	256	585	257
rect	585	13	586	14
rect	585	22	586	23
rect	585	34	586	35
rect	585	37	586	38
rect	585	40	586	41
rect	585	43	586	44
rect	585	46	586	47
rect	585	49	586	50
rect	585	52	586	53
rect	585	61	586	62
rect	585	64	586	65
rect	585	67	586	68
rect	585	70	586	71
rect	585	73	586	74
rect	585	76	586	77
rect	585	79	586	80
rect	585	94	586	95
rect	585	103	586	104
rect	585	106	586	107
rect	585	115	586	116
rect	585	118	586	119
rect	585	124	586	125
rect	585	145	586	146
rect	585	151	586	152
rect	585	154	586	155
rect	585	157	586	158
rect	585	160	586	161
rect	585	163	586	164
rect	585	166	586	167
rect	585	169	586	170
rect	585	184	586	185
rect	585	193	586	194
rect	585	196	586	197
rect	585	205	586	206
rect	585	214	586	215
rect	585	217	586	218
rect	585	226	586	227
rect	585	229	586	230
rect	585	238	586	239
rect	585	247	586	248
rect	585	250	586	251
rect	585	256	586	257
rect	586	13	587	14
rect	586	22	587	23
rect	586	31	587	32
rect	586	34	587	35
rect	586	37	587	38
rect	586	40	587	41
rect	586	43	587	44
rect	586	46	587	47
rect	586	49	587	50
rect	586	52	587	53
rect	586	61	587	62
rect	586	64	587	65
rect	586	67	587	68
rect	586	70	587	71
rect	586	73	587	74
rect	586	76	587	77
rect	586	79	587	80
rect	586	94	587	95
rect	586	103	587	104
rect	586	106	587	107
rect	586	115	587	116
rect	586	118	587	119
rect	586	124	587	125
rect	586	145	587	146
rect	586	151	587	152
rect	586	154	587	155
rect	586	157	587	158
rect	586	160	587	161
rect	586	163	587	164
rect	586	166	587	167
rect	586	169	587	170
rect	586	184	587	185
rect	586	193	587	194
rect	586	196	587	197
rect	586	205	587	206
rect	586	214	587	215
rect	586	217	587	218
rect	586	226	587	227
rect	586	229	587	230
rect	586	238	587	239
rect	586	247	587	248
rect	586	250	587	251
rect	586	256	587	257
rect	587	13	588	14
rect	587	22	588	23
rect	587	31	588	32
rect	587	34	588	35
rect	587	37	588	38
rect	587	40	588	41
rect	587	46	588	47
rect	587	49	588	50
rect	587	52	588	53
rect	587	61	588	62
rect	587	64	588	65
rect	587	70	588	71
rect	587	73	588	74
rect	587	76	588	77
rect	587	79	588	80
rect	587	94	588	95
rect	587	103	588	104
rect	587	106	588	107
rect	587	115	588	116
rect	587	118	588	119
rect	587	124	588	125
rect	587	145	588	146
rect	587	151	588	152
rect	587	154	588	155
rect	587	157	588	158
rect	587	160	588	161
rect	587	163	588	164
rect	587	166	588	167
rect	587	169	588	170
rect	587	184	588	185
rect	587	193	588	194
rect	587	196	588	197
rect	587	205	588	206
rect	587	214	588	215
rect	587	217	588	218
rect	587	226	588	227
rect	587	229	588	230
rect	587	238	588	239
rect	587	247	588	248
rect	587	250	588	251
rect	587	256	588	257
rect	588	13	589	14
rect	588	22	589	23
rect	588	25	589	26
rect	588	31	589	32
rect	588	34	589	35
rect	588	37	589	38
rect	588	40	589	41
rect	588	46	589	47
rect	588	49	589	50
rect	588	52	589	53
rect	588	55	589	56
rect	588	61	589	62
rect	588	64	589	65
rect	588	70	589	71
rect	588	73	589	74
rect	588	76	589	77
rect	588	79	589	80
rect	588	94	589	95
rect	588	103	589	104
rect	588	106	589	107
rect	588	115	589	116
rect	588	118	589	119
rect	588	124	589	125
rect	588	145	589	146
rect	588	151	589	152
rect	588	154	589	155
rect	588	157	589	158
rect	588	160	589	161
rect	588	163	589	164
rect	588	166	589	167
rect	588	169	589	170
rect	588	184	589	185
rect	588	193	589	194
rect	588	196	589	197
rect	588	205	589	206
rect	588	214	589	215
rect	588	217	589	218
rect	588	226	589	227
rect	588	229	589	230
rect	588	238	589	239
rect	588	247	589	248
rect	588	250	589	251
rect	588	256	589	257
rect	589	13	590	14
rect	589	22	590	23
rect	589	25	590	26
rect	589	31	590	32
rect	589	34	590	35
rect	589	37	590	38
rect	589	40	590	41
rect	589	49	590	50
rect	589	52	590	53
rect	589	55	590	56
rect	589	70	590	71
rect	589	73	590	74
rect	589	76	590	77
rect	589	94	590	95
rect	589	103	590	104
rect	589	106	590	107
rect	589	115	590	116
rect	589	118	590	119
rect	589	124	590	125
rect	589	145	590	146
rect	589	151	590	152
rect	589	154	590	155
rect	589	157	590	158
rect	589	160	590	161
rect	589	163	590	164
rect	589	166	590	167
rect	589	169	590	170
rect	589	184	590	185
rect	589	193	590	194
rect	589	196	590	197
rect	589	214	590	215
rect	589	217	590	218
rect	589	226	590	227
rect	589	229	590	230
rect	589	238	590	239
rect	589	247	590	248
rect	589	250	590	251
rect	589	256	590	257
rect	590	13	591	14
rect	590	22	591	23
rect	590	25	591	26
rect	590	31	591	32
rect	590	34	591	35
rect	590	37	591	38
rect	590	40	591	41
rect	590	43	591	44
rect	590	49	591	50
rect	590	52	591	53
rect	590	55	591	56
rect	590	67	591	68
rect	590	70	591	71
rect	590	73	591	74
rect	590	76	591	77
rect	590	94	591	95
rect	590	103	591	104
rect	590	106	591	107
rect	590	115	591	116
rect	590	118	591	119
rect	590	124	591	125
rect	590	145	591	146
rect	590	151	591	152
rect	590	154	591	155
rect	590	157	591	158
rect	590	160	591	161
rect	590	163	591	164
rect	590	166	591	167
rect	590	169	591	170
rect	590	184	591	185
rect	590	193	591	194
rect	590	196	591	197
rect	590	208	591	209
rect	590	214	591	215
rect	590	217	591	218
rect	590	226	591	227
rect	590	229	591	230
rect	590	238	591	239
rect	590	247	591	248
rect	590	250	591	251
rect	590	256	591	257
rect	591	13	592	14
rect	591	22	592	23
rect	591	25	592	26
rect	591	31	592	32
rect	591	34	592	35
rect	591	37	592	38
rect	591	40	592	41
rect	591	43	592	44
rect	591	49	592	50
rect	591	55	592	56
rect	591	67	592	68
rect	591	70	592	71
rect	591	73	592	74
rect	591	94	592	95
rect	591	106	592	107
rect	591	115	592	116
rect	591	118	592	119
rect	591	124	592	125
rect	591	145	592	146
rect	591	157	592	158
rect	591	160	592	161
rect	591	163	592	164
rect	591	166	592	167
rect	591	184	592	185
rect	591	193	592	194
rect	591	196	592	197
rect	591	208	592	209
rect	591	214	592	215
rect	591	226	592	227
rect	591	229	592	230
rect	591	247	592	248
rect	591	250	592	251
rect	591	256	592	257
rect	592	13	593	14
rect	592	22	593	23
rect	592	25	593	26
rect	592	31	593	32
rect	592	34	593	35
rect	592	37	593	38
rect	592	40	593	41
rect	592	43	593	44
rect	592	46	593	47
rect	592	49	593	50
rect	592	55	593	56
rect	592	64	593	65
rect	592	67	593	68
rect	592	70	593	71
rect	592	73	593	74
rect	592	94	593	95
rect	592	97	593	98
rect	592	106	593	107
rect	592	115	593	116
rect	592	118	593	119
rect	592	124	593	125
rect	592	145	593	146
rect	592	157	593	158
rect	592	160	593	161
rect	592	163	593	164
rect	592	166	593	167
rect	592	175	593	176
rect	592	184	593	185
rect	592	193	593	194
rect	592	196	593	197
rect	592	202	593	203
rect	592	208	593	209
rect	592	214	593	215
rect	592	223	593	224
rect	592	226	593	227
rect	592	229	593	230
rect	592	247	593	248
rect	592	250	593	251
rect	592	256	593	257
rect	593	13	594	14
rect	593	22	594	23
rect	593	25	594	26
rect	593	31	594	32
rect	593	34	594	35
rect	593	37	594	38
rect	593	40	594	41
rect	593	43	594	44
rect	593	46	594	47
rect	593	55	594	56
rect	593	64	594	65
rect	593	67	594	68
rect	593	70	594	71
rect	593	94	594	95
rect	593	97	594	98
rect	593	106	594	107
rect	593	118	594	119
rect	593	124	594	125
rect	593	145	594	146
rect	593	160	594	161
rect	593	163	594	164
rect	593	166	594	167
rect	593	175	594	176
rect	593	184	594	185
rect	593	196	594	197
rect	593	202	594	203
rect	593	208	594	209
rect	593	214	594	215
rect	593	223	594	224
rect	593	226	594	227
rect	593	247	594	248
rect	593	250	594	251
rect	593	256	594	257
rect	594	13	595	14
rect	594	22	595	23
rect	594	25	595	26
rect	594	28	595	29
rect	594	31	595	32
rect	594	34	595	35
rect	594	37	595	38
rect	594	40	595	41
rect	594	43	595	44
rect	594	46	595	47
rect	594	55	595	56
rect	594	61	595	62
rect	594	64	595	65
rect	594	67	595	68
rect	594	70	595	71
rect	594	94	595	95
rect	594	97	595	98
rect	594	103	595	104
rect	594	106	595	107
rect	594	118	595	119
rect	594	124	595	125
rect	594	142	595	143
rect	594	145	595	146
rect	594	160	595	161
rect	594	163	595	164
rect	594	166	595	167
rect	594	169	595	170
rect	594	175	595	176
rect	594	184	595	185
rect	594	196	595	197
rect	594	199	595	200
rect	594	202	595	203
rect	594	205	595	206
rect	594	208	595	209
rect	594	211	595	212
rect	594	214	595	215
rect	594	223	595	224
rect	594	226	595	227
rect	594	247	595	248
rect	594	250	595	251
rect	594	256	595	257
rect	595	13	596	14
rect	595	22	596	23
rect	595	25	596	26
rect	595	28	596	29
rect	595	31	596	32
rect	595	37	596	38
rect	595	40	596	41
rect	595	43	596	44
rect	595	46	596	47
rect	595	55	596	56
rect	595	61	596	62
rect	595	64	596	65
rect	595	67	596	68
rect	595	97	596	98
rect	595	103	596	104
rect	595	124	596	125
rect	595	142	596	143
rect	595	160	596	161
rect	595	169	596	170
rect	595	175	596	176
rect	595	184	596	185
rect	595	196	596	197
rect	595	199	596	200
rect	595	202	596	203
rect	595	205	596	206
rect	595	208	596	209
rect	595	211	596	212
rect	595	223	596	224
rect	596	13	597	14
rect	596	22	597	23
rect	596	25	597	26
rect	596	28	597	29
rect	596	31	597	32
rect	596	37	597	38
rect	596	40	597	41
rect	596	43	597	44
rect	596	46	597	47
rect	596	49	597	50
rect	596	55	597	56
rect	596	58	597	59
rect	596	61	597	62
rect	596	64	597	65
rect	596	67	597	68
rect	596	88	597	89
rect	596	97	597	98
rect	596	100	597	101
rect	596	103	597	104
rect	596	109	597	110
rect	596	124	597	125
rect	596	133	597	134
rect	596	142	597	143
rect	596	151	597	152
rect	596	160	597	161
rect	596	169	597	170
rect	596	172	597	173
rect	596	175	597	176
rect	596	184	597	185
rect	596	193	597	194
rect	596	196	597	197
rect	596	199	597	200
rect	596	202	597	203
rect	596	205	597	206
rect	596	208	597	209
rect	596	211	597	212
rect	596	220	597	221
rect	596	223	597	224
rect	596	238	597	239
rect	603	10	604	11
rect	603	13	604	14
rect	603	22	604	23
rect	603	25	604	26
rect	603	28	604	29
rect	603	31	604	32
rect	603	34	604	35
rect	603	40	604	41
rect	603	43	604	44
rect	603	46	604	47
rect	603	55	604	56
rect	603	58	604	59
rect	603	61	604	62
rect	603	64	604	65
rect	603	67	604	68
rect	603	88	604	89
rect	603	97	604	98
rect	603	100	604	101
rect	603	103	604	104
rect	603	106	604	107
rect	603	124	604	125
rect	603	133	604	134
rect	603	136	604	137
rect	603	142	604	143
rect	603	151	604	152
rect	603	160	604	161
rect	603	169	604	170
rect	603	172	604	173
rect	603	175	604	176
rect	603	184	604	185
rect	603	193	604	194
rect	603	196	604	197
rect	603	205	604	206
rect	603	208	604	209
rect	603	211	604	212
rect	603	220	604	221
rect	603	223	604	224
rect	603	226	604	227
rect	603	238	604	239
rect	604	10	605	11
rect	604	13	605	14
rect	604	25	605	26
rect	604	28	605	29
rect	604	31	605	32
rect	604	34	605	35
rect	604	40	605	41
rect	604	46	605	47
rect	604	55	605	56
rect	604	61	605	62
rect	604	64	605	65
rect	604	67	605	68
rect	604	88	605	89
rect	604	97	605	98
rect	604	100	605	101
rect	604	103	605	104
rect	604	106	605	107
rect	604	124	605	125
rect	604	133	605	134
rect	604	136	605	137
rect	604	142	605	143
rect	604	151	605	152
rect	604	160	605	161
rect	604	169	605	170
rect	604	172	605	173
rect	604	184	605	185
rect	604	193	605	194
rect	604	205	605	206
rect	604	208	605	209
rect	604	220	605	221
rect	604	223	605	224
rect	604	226	605	227
rect	604	238	605	239
rect	605	10	606	11
rect	605	13	606	14
rect	605	19	606	20
rect	605	25	606	26
rect	605	28	606	29
rect	605	31	606	32
rect	605	34	606	35
rect	605	37	606	38
rect	605	40	606	41
rect	605	46	606	47
rect	605	49	606	50
rect	605	55	606	56
rect	605	61	606	62
rect	605	64	606	65
rect	605	67	606	68
rect	605	88	606	89
rect	605	97	606	98
rect	605	100	606	101
rect	605	103	606	104
rect	605	106	606	107
rect	605	124	606	125
rect	605	133	606	134
rect	605	136	606	137
rect	605	142	606	143
rect	605	151	606	152
rect	605	160	606	161
rect	605	164	606	165
rect	605	169	606	170
rect	605	172	606	173
rect	605	178	606	179
rect	605	184	606	185
rect	605	193	606	194
rect	605	199	606	200
rect	605	205	606	206
rect	605	208	606	209
rect	605	220	606	221
rect	605	223	606	224
rect	605	226	606	227
rect	605	238	606	239
rect	606	10	607	11
rect	606	13	607	14
rect	606	19	607	20
rect	606	28	607	29
rect	606	31	607	32
rect	606	34	607	35
rect	606	37	607	38
rect	606	40	607	41
rect	606	46	607	47
rect	606	49	607	50
rect	606	61	607	62
rect	606	64	607	65
rect	606	100	607	101
rect	606	103	607	104
rect	606	124	607	125
rect	606	133	607	134
rect	606	136	607	137
rect	606	142	607	143
rect	606	151	607	152
rect	606	160	607	161
rect	606	164	607	165
rect	606	169	607	170
rect	606	172	607	173
rect	606	178	607	179
rect	606	193	607	194
rect	606	199	607	200
rect	606	208	607	209
rect	606	220	607	221
rect	606	223	607	224
rect	606	226	607	227
rect	606	238	607	239
rect	607	10	608	11
rect	607	13	608	14
rect	607	19	608	20
rect	607	22	608	23
rect	607	28	608	29
rect	607	31	608	32
rect	607	34	608	35
rect	607	37	608	38
rect	607	40	608	41
rect	607	43	608	44
rect	607	46	608	47
rect	607	49	608	50
rect	607	58	608	59
rect	607	61	608	62
rect	607	64	608	65
rect	607	85	608	86
rect	607	100	608	101
rect	607	103	608	104
rect	607	124	608	125
rect	607	133	608	134
rect	607	136	608	137
rect	607	142	608	143
rect	607	151	608	152
rect	607	160	608	161
rect	607	164	608	165
rect	607	169	608	170
rect	607	172	608	173
rect	607	175	608	176
rect	607	178	608	179
rect	607	193	608	194
rect	607	196	608	197
rect	607	199	608	200
rect	607	208	608	209
rect	607	220	608	221
rect	607	223	608	224
rect	607	226	608	227
rect	607	238	608	239
rect	608	13	609	14
rect	608	19	609	20
rect	608	22	609	23
rect	608	31	609	32
rect	608	37	609	38
rect	608	43	609	44
rect	608	46	609	47
rect	608	49	609	50
rect	608	58	609	59
rect	608	61	609	62
rect	608	85	609	86
rect	608	100	609	101
rect	608	124	609	125
rect	608	133	609	134
rect	608	151	609	152
rect	608	160	609	161
rect	608	169	609	170
rect	608	172	609	173
rect	608	175	609	176
rect	608	178	609	179
rect	608	196	609	197
rect	608	199	609	200
rect	608	223	609	224
rect	608	238	609	239
rect	609	7	610	8
rect	609	13	610	14
rect	609	19	610	20
rect	609	22	610	23
rect	609	25	610	26
rect	609	31	610	32
rect	609	37	610	38
rect	609	43	610	44
rect	609	46	610	47
rect	609	49	610	50
rect	609	55	610	56
rect	609	58	610	59
rect	609	61	610	62
rect	609	82	610	83
rect	609	85	610	86
rect	609	100	610	101
rect	609	124	610	125
rect	609	133	610	134
rect	609	151	610	152
rect	609	160	610	161
rect	609	169	610	170
rect	609	172	610	173
rect	609	175	610	176
rect	609	178	610	179
rect	609	184	610	185
rect	609	196	610	197
rect	609	199	610	200
rect	609	202	610	203
rect	609	211	610	212
rect	609	223	610	224
rect	609	238	610	239
rect	610	7	611	8
rect	610	19	611	20
rect	610	22	611	23
rect	610	25	611	26
rect	610	37	611	38
rect	610	43	611	44
rect	610	49	611	50
rect	610	55	611	56
rect	610	58	611	59
rect	610	82	611	83
rect	610	85	611	86
rect	610	175	611	176
rect	610	178	611	179
rect	610	184	611	185
rect	610	196	611	197
rect	610	199	611	200
rect	610	202	611	203
rect	610	211	611	212
rect	610	238	611	239
rect	611	7	612	8
rect	611	10	612	11
rect	611	19	612	20
rect	611	22	612	23
rect	611	25	612	26
rect	611	28	612	29
rect	611	37	612	38
rect	611	40	612	41
rect	611	43	612	44
rect	611	49	612	50
rect	611	52	612	53
rect	611	55	612	56
rect	611	58	612	59
rect	611	79	612	80
rect	611	82	612	83
rect	611	85	612	86
rect	611	118	612	119
rect	611	127	612	128
rect	611	142	612	143
rect	611	157	612	158
rect	611	166	612	167
rect	611	175	612	176
rect	611	178	612	179
rect	611	181	612	182
rect	611	184	612	185
rect	611	193	612	194
rect	611	196	612	197
rect	611	199	612	200
rect	611	202	612	203
rect	611	211	612	212
rect	611	238	612	239
rect	618	7	619	8
rect	618	10	619	11
rect	618	13	619	14
rect	618	19	619	20
rect	618	22	619	23
rect	618	25	619	26
rect	618	28	619	29
rect	618	37	619	38
rect	618	40	619	41
rect	618	46	619	47
rect	618	49	619	50
rect	618	52	619	53
rect	618	55	619	56
rect	618	58	619	59
rect	618	79	619	80
rect	618	82	619	83
rect	618	85	619	86
rect	618	103	619	104
rect	618	118	619	119
rect	618	127	619	128
rect	618	142	619	143
rect	618	157	619	158
rect	618	166	619	167
rect	618	175	619	176
rect	618	178	619	179
rect	618	181	619	182
rect	618	184	619	185
rect	618	187	619	188
rect	618	190	619	191
rect	618	193	619	194
rect	618	196	619	197
rect	618	199	619	200
rect	618	202	619	203
rect	618	211	619	212
rect	618	217	619	218
rect	618	238	619	239
rect	619	7	620	8
rect	619	10	620	11
rect	619	13	620	14
rect	619	19	620	20
rect	619	22	620	23
rect	619	25	620	26
rect	619	28	620	29
rect	619	37	620	38
rect	619	40	620	41
rect	619	46	620	47
rect	619	49	620	50
rect	619	52	620	53
rect	619	55	620	56
rect	619	58	620	59
rect	619	79	620	80
rect	619	82	620	83
rect	619	85	620	86
rect	619	103	620	104
rect	619	118	620	119
rect	619	127	620	128
rect	619	142	620	143
rect	619	157	620	158
rect	619	166	620	167
rect	619	178	620	179
rect	619	181	620	182
rect	619	184	620	185
rect	619	187	620	188
rect	619	193	620	194
rect	619	196	620	197
rect	619	199	620	200
rect	619	202	620	203
rect	619	211	620	212
rect	619	217	620	218
rect	619	238	620	239
rect	620	7	621	8
rect	620	10	621	11
rect	620	13	621	14
rect	620	19	621	20
rect	620	22	621	23
rect	620	25	621	26
rect	620	28	621	29
rect	620	37	621	38
rect	620	40	621	41
rect	620	46	621	47
rect	620	49	621	50
rect	620	52	621	53
rect	620	55	621	56
rect	620	58	621	59
rect	620	79	621	80
rect	620	82	621	83
rect	620	85	621	86
rect	620	103	621	104
rect	620	118	621	119
rect	620	127	621	128
rect	620	142	621	143
rect	620	157	621	158
rect	620	166	621	167
rect	620	178	621	179
rect	620	181	621	182
rect	620	184	621	185
rect	620	187	621	188
rect	620	193	621	194
rect	620	196	621	197
rect	620	199	621	200
rect	620	202	621	203
rect	620	211	621	212
rect	620	217	621	218
rect	620	238	621	239
rect	621	10	622	11
rect	621	19	622	20
rect	621	22	622	23
rect	621	25	622	26
rect	621	37	622	38
rect	621	40	622	41
rect	621	49	622	50
rect	621	55	622	56
rect	621	58	622	59
rect	621	79	622	80
rect	621	82	622	83
rect	621	85	622	86
rect	621	103	622	104
rect	621	118	622	119
rect	621	127	622	128
rect	621	142	622	143
rect	621	157	622	158
rect	621	166	622	167
rect	621	178	622	179
rect	621	181	622	182
rect	621	196	622	197
rect	621	199	622	200
rect	621	202	622	203
rect	621	211	622	212
rect	621	217	622	218
rect	621	238	622	239
rect	622	10	623	11
rect	622	16	623	17
rect	622	19	623	20
rect	622	22	623	23
rect	622	25	623	26
rect	622	37	623	38
rect	622	40	623	41
rect	622	49	623	50
rect	622	55	623	56
rect	622	58	623	59
rect	622	79	623	80
rect	622	82	623	83
rect	622	85	623	86
rect	622	103	623	104
rect	622	118	623	119
rect	622	127	623	128
rect	622	142	623	143
rect	622	157	623	158
rect	622	166	623	167
rect	622	175	623	176
rect	622	178	623	179
rect	622	181	623	182
rect	622	196	623	197
rect	622	199	623	200
rect	622	202	623	203
rect	622	211	623	212
rect	622	217	623	218
rect	622	238	623	239
rect	623	10	624	11
rect	623	16	624	17
rect	623	19	624	20
rect	623	22	624	23
rect	623	37	624	38
rect	623	49	624	50
rect	623	55	624	56
rect	623	82	624	83
rect	623	85	624	86
rect	623	103	624	104
rect	623	118	624	119
rect	623	127	624	128
rect	623	142	624	143
rect	623	157	624	158
rect	623	166	624	167
rect	623	175	624	176
rect	623	178	624	179
rect	623	199	624	200
rect	623	202	624	203
rect	623	211	624	212
rect	623	217	624	218
rect	623	238	624	239
rect	624	10	625	11
rect	624	13	625	14
rect	624	16	625	17
rect	624	19	625	20
rect	624	22	625	23
rect	624	28	625	29
rect	624	37	625	38
rect	624	46	625	47
rect	624	49	625	50
rect	624	55	625	56
rect	624	61	625	62
rect	624	82	625	83
rect	624	85	625	86
rect	624	103	625	104
rect	624	118	625	119
rect	624	127	625	128
rect	624	142	625	143
rect	624	157	625	158
rect	624	166	625	167
rect	624	172	625	173
rect	624	175	625	176
rect	624	178	625	179
rect	624	187	625	188
rect	624	199	625	200
rect	624	202	625	203
rect	624	211	625	212
rect	624	217	625	218
rect	624	238	625	239
rect	625	10	626	11
rect	625	13	626	14
rect	625	16	626	17
rect	625	19	626	20
rect	625	22	626	23
rect	625	28	626	29
rect	625	46	626	47
rect	625	49	626	50
rect	625	61	626	62
rect	625	82	626	83
rect	625	103	626	104
rect	625	118	626	119
rect	625	127	626	128
rect	625	142	626	143
rect	625	157	626	158
rect	625	166	626	167
rect	625	172	626	173
rect	625	175	626	176
rect	625	187	626	188
rect	625	199	626	200
rect	625	238	626	239
rect	626	10	627	11
rect	626	13	627	14
rect	626	16	627	17
rect	626	19	627	20
rect	626	22	627	23
rect	626	25	627	26
rect	626	28	627	29
rect	626	43	627	44
rect	626	46	627	47
rect	626	49	627	50
rect	626	61	627	62
rect	626	79	627	80
rect	626	82	627	83
rect	626	103	627	104
rect	626	118	627	119
rect	626	127	627	128
rect	626	142	627	143
rect	626	157	627	158
rect	626	166	627	167
rect	626	169	627	170
rect	626	172	627	173
rect	626	175	627	176
rect	626	187	627	188
rect	626	196	627	197
rect	626	199	627	200
rect	626	238	627	239
rect	627	10	628	11
rect	627	13	628	14
rect	627	16	628	17
rect	627	25	628	26
rect	627	28	628	29
rect	627	43	628	44
rect	627	46	628	47
rect	627	61	628	62
rect	627	79	628	80
rect	627	118	628	119
rect	627	166	628	167
rect	627	169	628	170
rect	627	172	628	173
rect	627	175	628	176
rect	627	187	628	188
rect	627	196	628	197
rect	628	7	629	8
rect	628	10	629	11
rect	628	13	629	14
rect	628	16	629	17
rect	628	25	629	26
rect	628	28	629	29
rect	628	34	629	35
rect	628	40	629	41
rect	628	43	629	44
rect	628	46	629	47
rect	628	61	629	62
rect	628	64	629	65
rect	628	79	629	80
rect	628	88	629	89
rect	628	109	629	110
rect	628	118	629	119
rect	628	133	629	134
rect	628	148	629	149
rect	628	163	629	164
rect	628	166	629	167
rect	628	169	629	170
rect	628	172	629	173
rect	628	175	629	176
rect	628	178	629	179
rect	628	184	629	185
rect	628	187	629	188
rect	628	196	629	197
rect	628	217	629	218
rect	635	13	636	14
rect	635	16	636	17
rect	635	25	636	26
rect	635	28	636	29
rect	635	43	636	44
rect	635	46	636	47
rect	635	52	636	53
rect	635	61	636	62
rect	635	64	636	65
rect	635	79	636	80
rect	635	85	636	86
rect	635	88	636	89
rect	635	109	636	110
rect	635	115	636	116
rect	635	118	636	119
rect	635	133	636	134
rect	635	148	636	149
rect	635	157	636	158
rect	635	163	636	164
rect	635	166	636	167
rect	635	169	636	170
rect	635	172	636	173
rect	635	175	636	176
rect	635	184	636	185
rect	635	187	636	188
rect	635	196	636	197
rect	635	217	636	218
rect	636	13	637	14
rect	636	16	637	17
rect	636	25	637	26
rect	636	28	637	29
rect	636	43	637	44
rect	636	46	637	47
rect	636	52	637	53
rect	636	61	637	62
rect	636	64	637	65
rect	636	79	637	80
rect	636	85	637	86
rect	636	88	637	89
rect	636	109	637	110
rect	636	115	637	116
rect	636	118	637	119
rect	636	133	637	134
rect	636	148	637	149
rect	636	157	637	158
rect	636	163	637	164
rect	636	169	637	170
rect	636	172	637	173
rect	636	184	637	185
rect	636	187	637	188
rect	636	196	637	197
rect	636	217	637	218
rect	637	13	638	14
rect	637	16	638	17
rect	637	25	638	26
rect	637	28	638	29
rect	637	43	638	44
rect	637	46	638	47
rect	637	52	638	53
rect	637	61	638	62
rect	637	64	638	65
rect	637	79	638	80
rect	637	85	638	86
rect	637	88	638	89
rect	637	109	638	110
rect	637	115	638	116
rect	637	118	638	119
rect	637	133	638	134
rect	637	148	638	149
rect	637	157	638	158
rect	637	160	638	161
rect	637	163	638	164
rect	637	169	638	170
rect	637	172	638	173
rect	637	178	638	179
rect	637	184	638	185
rect	637	187	638	188
rect	637	196	638	197
rect	637	217	638	218
rect	638	13	639	14
rect	638	16	639	17
rect	638	25	639	26
rect	638	28	639	29
rect	638	43	639	44
rect	638	46	639	47
rect	638	52	639	53
rect	638	61	639	62
rect	638	64	639	65
rect	638	79	639	80
rect	638	85	639	86
rect	638	88	639	89
rect	638	109	639	110
rect	638	115	639	116
rect	638	118	639	119
rect	638	133	639	134
rect	638	148	639	149
rect	638	160	639	161
rect	638	163	639	164
rect	638	169	639	170
rect	638	172	639	173
rect	638	178	639	179
rect	638	184	639	185
rect	638	187	639	188
rect	638	217	639	218
rect	639	13	640	14
rect	639	16	640	17
rect	639	25	640	26
rect	639	28	640	29
rect	639	43	640	44
rect	639	46	640	47
rect	639	52	640	53
rect	639	61	640	62
rect	639	64	640	65
rect	639	79	640	80
rect	639	85	640	86
rect	639	88	640	89
rect	639	109	640	110
rect	639	115	640	116
rect	639	118	640	119
rect	639	133	640	134
rect	639	148	640	149
rect	639	160	640	161
rect	639	163	640	164
rect	639	169	640	170
rect	639	172	640	173
rect	639	178	640	179
rect	639	184	640	185
rect	639	187	640	188
rect	639	217	640	218
rect	640	13	641	14
rect	640	16	641	17
rect	640	25	641	26
rect	640	28	641	29
rect	640	43	641	44
rect	640	46	641	47
rect	640	52	641	53
rect	640	61	641	62
rect	640	64	641	65
rect	640	85	641	86
rect	640	88	641	89
rect	640	109	641	110
rect	640	115	641	116
rect	640	118	641	119
rect	640	133	641	134
rect	640	148	641	149
rect	640	160	641	161
rect	640	163	641	164
rect	640	169	641	170
rect	640	172	641	173
rect	640	178	641	179
rect	640	184	641	185
rect	640	217	641	218
rect	641	13	642	14
rect	641	16	642	17
rect	641	25	642	26
rect	641	28	642	29
rect	641	43	642	44
rect	641	46	642	47
rect	641	52	642	53
rect	641	55	642	56
rect	641	61	642	62
rect	641	64	642	65
rect	641	85	642	86
rect	641	88	642	89
rect	641	109	642	110
rect	641	115	642	116
rect	641	118	642	119
rect	641	133	642	134
rect	641	148	642	149
rect	641	157	642	158
rect	641	160	642	161
rect	641	163	642	164
rect	641	169	642	170
rect	641	172	642	173
rect	641	178	642	179
rect	641	184	642	185
rect	641	217	642	218
rect	642	13	643	14
rect	642	16	643	17
rect	642	25	643	26
rect	642	28	643	29
rect	642	43	643	44
rect	642	46	643	47
rect	642	55	643	56
rect	642	61	643	62
rect	642	64	643	65
rect	642	85	643	86
rect	642	88	643	89
rect	642	109	643	110
rect	642	115	643	116
rect	642	118	643	119
rect	642	133	643	134
rect	642	148	643	149
rect	642	157	643	158
rect	642	160	643	161
rect	642	163	643	164
rect	642	169	643	170
rect	642	172	643	173
rect	642	178	643	179
rect	642	184	643	185
rect	643	13	644	14
rect	643	16	644	17
rect	643	25	644	26
rect	643	28	644	29
rect	643	43	644	44
rect	643	46	644	47
rect	643	55	644	56
rect	643	61	644	62
rect	643	64	644	65
rect	643	85	644	86
rect	643	88	644	89
rect	643	109	644	110
rect	643	115	644	116
rect	643	118	644	119
rect	643	133	644	134
rect	643	148	644	149
rect	643	157	644	158
rect	643	160	644	161
rect	643	163	644	164
rect	643	169	644	170
rect	643	172	644	173
rect	643	178	644	179
rect	643	184	644	185
rect	644	13	645	14
rect	644	25	645	26
rect	644	43	645	44
rect	644	55	645	56
rect	644	61	645	62
rect	644	85	645	86
rect	644	88	645	89
rect	644	118	645	119
rect	644	133	645	134
rect	644	157	645	158
rect	644	160	645	161
rect	644	169	645	170
rect	644	178	645	179
rect	644	184	645	185
rect	645	10	646	11
rect	645	13	646	14
rect	645	22	646	23
rect	645	25	646	26
rect	645	37	646	38
rect	645	43	646	44
rect	645	49	646	50
rect	645	55	646	56
rect	645	61	646	62
rect	645	85	646	86
rect	645	88	646	89
rect	645	118	646	119
rect	645	133	646	134
rect	645	139	646	140
rect	645	151	646	152
rect	645	157	646	158
rect	645	160	646	161
rect	645	169	646	170
rect	645	175	646	176
rect	645	178	646	179
rect	645	184	646	185
rect	646	10	647	11
rect	646	22	647	23
rect	646	37	647	38
rect	646	49	647	50
rect	646	55	647	56
rect	646	139	647	140
rect	646	151	647	152
rect	646	157	647	158
rect	646	160	647	161
rect	646	169	647	170
rect	646	175	647	176
rect	646	178	647	179
rect	647	7	648	8
rect	647	10	648	11
rect	647	19	648	20
rect	647	22	648	23
rect	647	37	648	38
rect	647	40	648	41
rect	647	46	648	47
rect	647	49	648	50
rect	647	55	648	56
rect	647	79	648	80
rect	647	82	648	83
rect	647	115	648	116
rect	647	124	648	125
rect	647	139	648	140
rect	647	148	648	149
rect	647	151	648	152
rect	647	157	648	158
rect	647	160	648	161
rect	647	169	648	170
rect	647	175	648	176
rect	647	178	648	179
rect	654	4	655	5
rect	654	7	655	8
rect	654	10	655	11
rect	654	13	655	14
rect	654	19	655	20
rect	654	22	655	23
rect	654	37	655	38
rect	654	43	655	44
rect	654	46	655	47
rect	654	49	655	50
rect	654	82	655	83
rect	654	115	655	116
rect	654	124	655	125
rect	654	139	655	140
rect	654	148	655	149
rect	654	151	655	152
rect	654	154	655	155
rect	654	160	655	161
rect	654	169	655	170
rect	655	4	656	5
rect	655	7	656	8
rect	655	10	656	11
rect	655	13	656	14
rect	655	19	656	20
rect	655	22	656	23
rect	655	37	656	38
rect	655	43	656	44
rect	655	46	656	47
rect	655	49	656	50
rect	655	82	656	83
rect	655	115	656	116
rect	655	124	656	125
rect	655	139	656	140
rect	655	151	656	152
rect	655	160	656	161
rect	655	169	656	170
rect	656	4	657	5
rect	656	7	657	8
rect	656	10	657	11
rect	656	13	657	14
rect	656	19	657	20
rect	656	22	657	23
rect	656	37	657	38
rect	656	43	657	44
rect	656	46	657	47
rect	656	49	657	50
rect	656	82	657	83
rect	656	115	657	116
rect	656	124	657	125
rect	656	139	657	140
rect	656	151	657	152
rect	656	160	657	161
rect	656	169	657	170
rect	657	10	658	11
rect	657	22	658	23
rect	657	37	658	38
rect	657	43	658	44
rect	657	46	658	47
rect	657	82	658	83
rect	657	115	658	116
rect	657	124	658	125
rect	657	139	658	140
rect	657	160	658	161
rect	657	169	658	170
rect	658	10	659	11
rect	658	22	659	23
rect	658	31	659	32
rect	658	37	659	38
rect	658	43	659	44
rect	658	46	659	47
rect	658	82	659	83
rect	658	115	659	116
rect	658	124	659	125
rect	658	136	659	137
rect	658	139	659	140
rect	658	160	659	161
rect	658	169	659	170
rect	659	31	660	32
rect	659	115	660	116
rect	659	124	660	125
rect	659	136	660	137
rect	659	139	660	140
rect	660	7	661	8
rect	660	13	661	14
rect	660	28	661	29
rect	660	31	661	32
rect	660	64	661	65
rect	660	85	661	86
rect	660	115	661	116
rect	660	124	661	125
rect	660	136	661	137
rect	660	139	661	140
rect	660	166	661	167
rect	667	4	668	5
rect	667	7	668	8
rect	667	25	668	26
rect	667	28	668	29
rect	667	82	668	83
rect	667	88	668	89
rect	667	115	668	116
rect	667	124	668	125
rect	667	130	668	131
rect	667	139	668	140
rect	667	142	668	143
rect	667	166	668	167
rect	668	4	669	5
rect	668	7	669	8
rect	668	25	669	26
rect	668	28	669	29
rect	668	82	669	83
rect	668	166	669	167
rect	669	4	670	5
rect	669	7	670	8
rect	669	25	670	26
rect	669	28	670	29
rect	669	82	670	83
rect	669	166	670	167
<< via >>
rect	0	121	1	122
rect	0	172	1	173
rect	2	52	3	53
rect	2	58	3	59
rect	2	109	3	110
rect	2	115	3	116
rect	2	118	3	119
rect	2	124	3	125
rect	2	136	3	137
rect	2	145	3	146
rect	4	7	5	8
rect	4	79	5	80
rect	4	85	5	86
rect	4	91	5	92
rect	4	106	5	107
rect	4	142	5	143
rect	13	130	14	131
rect	13	202	14	203
rect	15	121	16	122
rect	15	211	16	212
rect	17	79	18	80
rect	17	85	18	86
rect	17	100	18	101
rect	17	106	18	107
rect	17	118	18	119
rect	17	130	18	131
rect	17	172	18	173
rect	17	178	18	179
rect	19	76	20	77
rect	19	175	20	176
rect	21	25	22	26
rect	21	214	22	215
rect	23	13	24	14
rect	23	172	24	173
rect	25	4	26	5
rect	25	52	26	53
rect	25	73	26	74
rect	25	82	26	83
rect	25	94	26	95
rect	25	106	26	107
rect	25	109	26	110
rect	25	121	26	122
rect	25	124	26	125
rect	25	136	26	137
rect	27	1	28	2
rect	27	7	28	8
rect	27	10	28	11
rect	27	13	28	14
rect	27	16	28	17
rect	27	22	28	23
rect	27	25	28	26
rect	27	28	28	29
rect	27	52	28	53
rect	27	55	28	56
rect	27	67	28	68
rect	27	79	28	80
rect	27	91	28	92
rect	27	109	28	110
rect	27	118	28	119
rect	27	127	28	128
rect	27	133	28	134
rect	27	139	28	140
rect	27	145	28	146
rect	27	163	28	164
rect	27	187	28	188
rect	27	190	28	191
rect	36	130	37	131
rect	36	142	37	143
rect	38	130	39	131
rect	38	136	39	137
rect	40	118	41	119
rect	40	154	41	155
rect	40	157	41	158
rect	40	199	41	200
rect	42	82	43	83
rect	42	103	43	104
rect	42	112	43	113
rect	42	169	43	170
rect	44	52	45	53
rect	44	55	45	56
rect	44	61	45	62
rect	44	67	45	68
rect	44	79	45	80
rect	44	100	45	101
rect	44	109	45	110
rect	44	124	45	125
rect	44	127	45	128
rect	44	133	45	134
rect	44	145	45	146
rect	44	157	45	158
rect	44	187	45	188
rect	44	208	45	209
rect	46	13	47	14
rect	46	16	47	17
rect	46	22	47	23
rect	46	31	47	32
rect	46	34	47	35
rect	46	193	47	194
rect	48	10	49	11
rect	48	145	49	146
rect	48	175	49	176
rect	48	190	49	191
rect	48	211	49	212
rect	48	238	49	239
rect	50	7	51	8
rect	50	13	51	14
rect	50	19	51	20
rect	50	25	51	26
rect	50	28	51	29
rect	50	40	51	41
rect	50	46	51	47
rect	50	64	51	65
rect	50	76	51	77
rect	50	85	51	86
rect	50	91	51	92
rect	50	97	51	98
rect	50	106	51	107
rect	50	139	51	140
rect	50	163	51	164
rect	50	166	51	167
rect	50	172	51	173
rect	50	187	51	188
rect	50	202	51	203
rect	50	211	51	212
rect	50	214	51	215
rect	50	241	51	242
rect	59	199	60	200
rect	59	232	60	233
rect	61	106	62	107
rect	61	121	62	122
rect	61	190	62	191
rect	61	199	62	200
rect	63	103	64	104
rect	63	205	64	206
rect	65	5	66	6
rect	65	28	66	29
rect	65	103	66	104
rect	65	112	66	113
rect	65	154	66	155
rect	65	166	66	167
rect	65	175	66	176
rect	65	196	66	197
rect	65	211	66	212
rect	65	217	66	218
rect	67	16	68	17
rect	67	28	68	29
rect	67	40	68	41
rect	67	49	68	50
rect	67	100	68	101
rect	67	118	68	119
rect	67	121	68	122
rect	67	127	68	128
rect	67	139	68	140
rect	67	154	68	155
rect	67	175	68	176
rect	67	178	68	179
rect	67	187	68	188
rect	67	211	68	212
rect	69	13	70	14
rect	69	25	70	26
rect	69	31	70	32
rect	69	40	70	41
rect	69	67	70	68
rect	69	73	70	74
rect	69	100	70	101
rect	69	112	70	113
rect	69	127	70	128
rect	69	130	70	131
rect	69	139	70	140
rect	69	142	70	143
rect	69	178	70	179
rect	69	181	70	182
rect	69	184	70	185
rect	69	190	70	191
rect	69	241	70	242
rect	69	289	70	290
rect	71	7	72	8
rect	71	16	72	17
rect	71	19	72	20
rect	71	31	72	32
rect	71	64	72	65
rect	71	82	72	83
rect	71	85	72	86
rect	71	91	72	92
rect	71	97	72	98
rect	71	115	72	116
rect	71	130	72	131
rect	71	136	72	137
rect	71	142	72	143
rect	71	145	72	146
rect	71	172	72	173
rect	71	193	72	194
rect	71	208	72	209
rect	71	214	72	215
rect	71	223	72	224
rect	71	229	72	230
rect	71	238	72	239
rect	71	286	72	287
rect	73	5	74	6
rect	73	7	74	8
rect	73	10	74	11
rect	73	19	74	20
rect	73	22	74	23
rect	73	34	74	35
rect	73	55	74	56
rect	73	58	74	59
rect	73	61	74	62
rect	73	67	74	68
rect	73	70	74	71
rect	73	76	74	77
rect	73	79	74	80
rect	73	145	74	146
rect	73	163	74	164
rect	73	187	74	188
rect	73	208	74	209
rect	73	226	74	227
rect	73	238	74	239
rect	73	241	74	242
rect	82	118	83	119
rect	82	130	83	131
rect	82	208	83	209
rect	82	226	83	227
rect	84	118	85	119
rect	84	127	85	128
rect	84	208	85	209
rect	84	214	85	215
rect	86	115	87	116
rect	86	127	87	128
rect	86	196	87	197
rect	86	214	87	215
rect	86	217	87	218
rect	86	235	87	236
rect	88	40	89	41
rect	88	46	89	47
rect	88	73	89	74
rect	88	76	89	77
rect	88	106	89	107
rect	88	115	89	116
rect	88	196	89	197
rect	88	205	89	206
rect	88	211	89	212
rect	88	250	89	251
rect	90	25	91	26
rect	90	43	91	44
rect	90	49	91	50
rect	90	61	91	62
rect	90	67	91	68
rect	90	85	91	86
rect	90	91	91	92
rect	90	109	91	110
rect	90	145	91	146
rect	90	148	91	149
rect	90	202	91	203
rect	90	205	91	206
rect	90	211	91	212
rect	90	220	91	221
rect	90	268	91	269
rect	90	277	91	278
rect	92	19	93	20
rect	92	25	93	26
rect	92	28	93	29
rect	92	49	93	50
rect	92	67	93	68
rect	92	181	93	182
rect	92	199	93	200
rect	92	217	93	218
rect	92	232	93	233
rect	92	238	93	239
rect	92	253	93	254
rect	92	268	93	269
rect	94	10	95	11
rect	94	22	95	23
rect	94	28	95	29
rect	94	31	95	32
rect	94	34	95	35
rect	94	40	95	41
rect	94	58	95	59
rect	94	73	95	74
rect	94	82	95	83
rect	94	94	95	95
rect	94	103	95	104
rect	94	106	95	107
rect	94	142	95	143
rect	94	145	95	146
rect	94	157	95	158
rect	94	163	95	164
rect	94	187	95	188
rect	94	220	95	221
rect	94	229	95	230
rect	94	253	95	254
rect	94	292	95	293
rect	94	298	95	299
rect	96	7	97	8
rect	96	13	97	14
rect	96	16	97	17
rect	96	22	97	23
rect	96	31	97	32
rect	96	34	97	35
rect	96	55	97	56
rect	96	58	97	59
rect	96	64	97	65
rect	96	70	97	71
rect	96	79	97	80
rect	96	103	97	104
rect	96	139	97	140
rect	96	142	97	143
rect	96	154	97	155
rect	96	160	97	161
rect	96	178	97	179
rect	96	187	97	188
rect	96	193	97	194
rect	96	232	97	233
rect	96	289	97	290
rect	96	310	97	311
rect	98	7	99	8
rect	98	100	99	101
rect	98	112	99	113
rect	98	121	99	122
rect	98	124	99	125
rect	98	133	99	134
rect	98	136	99	137
rect	98	157	99	158
rect	98	166	99	167
rect	98	172	99	173
rect	98	175	99	176
rect	98	184	99	185
rect	98	190	99	191
rect	98	229	99	230
rect	98	286	99	287
rect	98	307	99	308
rect	107	101	108	102
rect	107	148	108	149
rect	109	148	110	149
rect	109	154	110	155
rect	111	101	112	102
rect	111	154	112	155
rect	113	103	114	104
rect	113	121	114	122
rect	113	244	114	245
rect	113	250	114	251
rect	115	103	116	104
rect	115	112	116	113
rect	115	115	116	116
rect	115	124	116	125
rect	115	235	116	236
rect	115	250	116	251
rect	117	112	118	113
rect	117	175	118	176
rect	117	217	118	218
rect	117	235	118	236
rect	117	274	118	275
rect	117	277	118	278
rect	119	58	120	59
rect	119	166	120	167
rect	119	205	120	206
rect	119	217	120	218
rect	119	253	120	254
rect	119	277	120	278
rect	121	109	122	110
rect	121	115	122	116
rect	121	145	122	146
rect	121	151	122	152
rect	121	157	122	158
rect	121	166	122	167
rect	121	181	122	182
rect	121	205	122	206
rect	121	247	122	248
rect	121	271	122	272
rect	123	85	124	86
rect	123	91	124	92
rect	123	109	124	110
rect	123	118	124	119
rect	123	136	124	137
rect	123	157	124	158
rect	123	172	124	173
rect	123	181	124	182
rect	123	208	124	209
rect	123	223	124	224
rect	123	232	124	233
rect	123	256	124	257
rect	125	55	126	56
rect	125	64	126	65
rect	125	73	126	74
rect	125	85	126	86
rect	125	106	126	107
rect	125	118	126	119
rect	125	133	126	134
rect	125	145	126	146
rect	125	169	126	170
rect	125	208	126	209
rect	125	214	126	215
rect	125	232	126	233
rect	125	241	126	242
rect	125	262	126	263
rect	127	49	128	50
rect	127	58	128	59
rect	127	70	128	71
rect	127	292	128	293
rect	129	37	130	38
rect	129	88	130	89
rect	129	94	130	95
rect	129	106	130	107
rect	129	130	130	131
rect	129	139	130	140
rect	129	163	130	164
rect	129	175	130	176
rect	129	214	130	215
rect	129	226	130	227
rect	129	238	130	239
rect	129	259	130	260
rect	131	31	132	32
rect	131	37	132	38
rect	131	46	132	47
rect	131	52	132	53
rect	131	64	132	65
rect	131	286	132	287
rect	133	28	134	29
rect	133	34	134	35
rect	133	43	134	44
rect	133	49	134	50
rect	133	61	134	62
rect	133	73	134	74
rect	133	94	134	95
rect	133	97	134	98
rect	133	127	134	128
rect	133	136	134	137
rect	133	160	134	161
rect	133	178	134	179
rect	133	211	134	212
rect	133	220	134	221
rect	133	229	134	230
rect	133	253	134	254
rect	133	310	134	311
rect	133	316	134	317
rect	135	13	136	14
rect	135	16	136	17
rect	135	25	136	26
rect	135	31	136	32
rect	135	40	136	41
rect	135	46	136	47
rect	135	61	136	62
rect	135	271	136	272
rect	135	298	136	299
rect	135	301	136	302
rect	135	307	136	308
rect	135	313	136	314
rect	137	10	138	11
rect	137	13	138	14
rect	137	22	138	23
rect	137	265	138	266
rect	137	292	138	293
rect	137	310	138	311
rect	146	130	147	131
rect	146	157	147	158
rect	148	151	149	152
rect	148	157	149	158
rect	150	142	151	143
rect	150	151	151	152
rect	152	127	153	128
rect	152	142	153	143
rect	152	286	153	287
rect	152	292	153	293
rect	154	61	155	62
rect	154	70	155	71
rect	154	106	155	107
rect	154	127	155	128
rect	154	277	155	278
rect	154	292	155	293
rect	156	58	157	59
rect	156	61	157	62
rect	156	91	157	92
rect	156	106	157	107
rect	156	259	157	260
rect	156	277	157	278
rect	158	52	159	53
rect	158	58	159	59
rect	158	73	159	74
rect	158	91	159	92
rect	158	154	159	155
rect	158	160	159	161
rect	158	214	159	215
rect	158	217	159	218
rect	158	253	159	254
rect	158	259	159	260
rect	160	34	161	35
rect	160	40	161	41
rect	160	52	161	53
rect	160	55	161	56
rect	160	73	161	74
rect	160	76	161	77
rect	160	83	161	84
rect	160	88	161	89
rect	160	148	161	149
rect	160	154	161	155
rect	160	172	161	173
rect	160	175	161	176
rect	160	205	161	206
rect	160	214	161	215
rect	160	244	161	245
rect	160	253	161	254
rect	162	34	163	35
rect	162	163	163	164
rect	162	166	163	167
rect	162	175	163	176
rect	162	178	163	179
rect	162	205	163	206
rect	162	217	163	218
rect	162	220	163	221
rect	162	241	163	242
rect	162	247	163	248
rect	164	19	165	20
rect	164	76	165	77
rect	164	88	165	89
rect	164	103	165	104
rect	164	139	165	140
rect	164	307	165	308
rect	166	16	167	17
rect	166	19	167	20
rect	166	31	167	32
rect	166	199	167	200
rect	166	208	167	209
rect	166	220	167	221
rect	166	232	167	233
rect	166	265	167	266
rect	166	289	167	290
rect	166	304	167	305
rect	166	313	167	314
rect	166	322	167	323
rect	168	13	169	14
rect	168	16	169	17
rect	168	28	169	29
rect	168	37	169	38
rect	168	49	169	50
rect	168	55	169	56
rect	168	83	169	84
rect	168	103	169	104
rect	168	112	169	113
rect	168	115	169	116
rect	168	136	169	137
rect	168	178	169	179
rect	168	181	169	182
rect	168	208	169	209
rect	168	229	169	230
rect	168	250	169	251
rect	168	262	169	263
rect	168	289	169	290
rect	168	295	169	296
rect	168	301	169	302
rect	168	310	169	311
rect	168	328	169	329
rect	170	10	171	11
rect	170	13	171	14
rect	170	25	171	26
rect	170	37	171	38
rect	170	46	171	47
rect	170	49	171	50
rect	170	97	171	98
rect	170	118	171	119
rect	170	121	171	122
rect	170	139	171	140
rect	170	145	171	146
rect	170	181	171	182
rect	170	223	171	224
rect	170	232	171	233
rect	170	235	171	236
rect	170	244	171	245
rect	170	256	171	257
rect	170	262	171	263
rect	170	271	171	272
rect	170	283	171	284
rect	170	286	171	287
rect	170	298	171	299
rect	170	307	171	308
rect	170	313	171	314
rect	170	316	171	317
rect	170	325	171	326
rect	179	181	180	182
rect	179	199	180	200
rect	181	85	182	86
rect	181	100	182	101
rect	181	160	182	161
rect	181	181	182	182
rect	181	313	182	314
rect	181	319	182	320
rect	183	16	184	17
rect	183	268	184	269
rect	183	304	184	305
rect	183	316	184	317
rect	185	91	186	92
rect	185	100	186	101
rect	185	106	186	107
rect	185	124	186	125
rect	185	157	186	158
rect	185	160	186	161
rect	185	268	186	269
rect	185	274	186	275
rect	185	301	186	302
rect	185	313	186	314
rect	187	44	188	45
rect	187	49	188	50
rect	187	82	188	83
rect	187	304	188	305
rect	189	37	190	38
rect	189	46	190	47
rect	189	61	190	62
rect	189	67	190	68
rect	189	76	190	77
rect	189	91	190	92
rect	189	106	190	107
rect	189	112	190	113
rect	189	139	190	140
rect	189	157	190	158
rect	189	175	190	176
rect	189	193	190	194
rect	189	211	190	212
rect	189	277	190	278
rect	189	292	190	293
rect	189	301	190	302
rect	191	19	192	20
rect	191	25	192	26
rect	191	31	192	32
rect	191	121	192	122
rect	191	127	192	128
rect	191	139	192	140
rect	191	166	192	167
rect	191	187	192	188
rect	191	190	192	191
rect	191	196	192	197
rect	191	214	192	215
rect	191	226	192	227
rect	191	265	192	266
rect	191	277	192	278
rect	191	289	192	290
rect	191	298	192	299
rect	191	328	192	329
rect	191	334	192	335
rect	193	16	194	17
rect	193	19	194	20
rect	193	28	194	29
rect	193	37	194	38
rect	193	49	194	50
rect	193	52	194	53
rect	193	58	194	59
rect	193	64	194	65
rect	193	73	194	74
rect	193	79	194	80
rect	193	82	194	83
rect	193	88	194	89
rect	193	103	194	104
rect	193	115	194	116
rect	193	118	194	119
rect	193	136	194	137
rect	193	154	194	155
rect	193	175	194	176
rect	193	178	194	179
rect	193	196	194	197
rect	193	214	194	215
rect	193	217	194	218
rect	193	223	194	224
rect	193	229	194	230
rect	193	238	194	239
rect	193	241	194	242
rect	193	259	194	260
rect	193	271	194	272
rect	193	286	194	287
rect	193	295	194	296
rect	193	325	194	326
rect	193	331	194	332
rect	195	13	196	14
rect	195	22	196	23
rect	195	28	196	29
rect	195	40	196	41
rect	195	44	196	45
rect	195	52	196	53
rect	195	55	196	56
rect	195	61	196	62
rect	195	70	196	71
rect	195	76	196	77
rect	195	88	196	89
rect	195	94	196	95
rect	195	103	196	104
rect	195	109	196	110
rect	195	127	196	128
rect	195	130	196	131
rect	195	133	196	134
rect	195	136	196	137
rect	195	145	196	146
rect	195	151	196	152
rect	195	154	196	155
rect	195	172	196	173
rect	195	178	196	179
rect	195	184	196	185
rect	195	205	196	206
rect	195	217	196	218
rect	195	229	196	230
rect	195	232	196	233
rect	195	235	196	236
rect	195	241	196	242
rect	195	253	196	254
rect	195	259	196	260
rect	195	262	196	263
rect	195	274	196	275
rect	195	286	196	287
rect	195	292	196	293
rect	195	322	196	323
rect	195	328	196	329
rect	204	142	205	143
rect	204	151	205	152
rect	206	127	207	128
rect	206	142	207	143
rect	208	94	209	95
rect	208	100	209	101
rect	208	124	209	125
rect	208	127	209	128
rect	208	199	209	200
rect	208	205	209	206
rect	210	91	211	92
rect	210	100	211	101
rect	210	121	211	122
rect	210	124	211	125
rect	210	181	211	182
rect	210	187	211	188
rect	210	196	211	197
rect	210	202	211	203
rect	212	61	213	62
rect	212	256	213	257
rect	214	61	215	62
rect	214	229	215	230
rect	216	22	217	23
rect	216	265	217	266
rect	218	19	219	20
rect	218	31	219	32
rect	218	37	219	38
rect	218	40	219	41
rect	218	79	219	80
rect	218	82	219	83
rect	218	91	219	92
rect	218	103	219	104
rect	218	106	219	107
rect	218	112	219	113
rect	218	121	219	122
rect	218	154	219	155
rect	218	157	219	158
rect	218	169	219	170
rect	218	181	219	182
rect	218	190	219	191
rect	218	196	219	197
rect	218	214	219	215
rect	218	217	219	218
rect	218	229	219	230
rect	218	244	219	245
rect	218	250	219	251
rect	218	274	219	275
rect	218	280	219	281
rect	220	19	221	20
rect	220	28	221	29
rect	220	34	221	35
rect	220	49	221	50
rect	220	67	221	68
rect	220	106	221	107
rect	220	109	221	110
rect	220	118	221	119
rect	220	139	221	140
rect	220	154	221	155
rect	220	157	221	158
rect	220	160	221	161
rect	220	163	221	164
rect	220	172	221	173
rect	220	178	221	179
rect	220	184	221	185
rect	220	193	221	194
rect	220	217	221	218
rect	220	241	221	242
rect	220	244	221	245
rect	220	247	221	248
rect	220	268	221	269
rect	220	274	221	275
rect	220	277	221	278
rect	220	292	221	293
rect	220	295	221	296
rect	222	10	223	11
rect	222	238	223	239
rect	222	241	223	242
rect	222	262	223	263
rect	222	271	223	272
rect	222	277	223	278
rect	222	283	223	284
rect	222	289	223	290
rect	222	295	223	296
rect	222	304	223	305
rect	222	313	223	314
rect	222	325	223	326
rect	224	28	225	29
rect	224	211	225	212
rect	224	238	225	239
rect	224	253	225	254
rect	224	259	225	260
rect	224	265	225	266
rect	224	271	225	272
rect	224	298	225	299
rect	224	304	225	305
rect	224	316	225	317
rect	226	4	227	5
rect	226	7	227	8
rect	226	10	227	11
rect	226	16	227	17
rect	226	25	227	26
rect	226	37	227	38
rect	226	46	227	47
rect	226	49	227	50
rect	226	52	227	53
rect	226	58	227	59
rect	226	64	227	65
rect	226	67	227	68
rect	226	70	227	71
rect	226	79	227	80
rect	226	88	227	89
rect	226	97	227	98
rect	226	115	227	116
rect	226	118	227	119
rect	226	139	227	140
rect	226	145	227	146
rect	226	160	227	161
rect	226	166	227	167
rect	226	175	227	176
rect	226	199	227	200
rect	226	232	227	233
rect	226	253	227	254
rect	226	256	227	257
rect	226	262	227	263
rect	226	268	227	269
rect	226	286	227	287
rect	226	301	227	302
rect	226	313	227	314
rect	235	94	236	95
rect	235	118	236	119
rect	235	193	236	194
rect	235	217	236	218
rect	237	5	238	6
rect	237	19	238	20
rect	237	76	238	77
rect	237	94	238	95
rect	237	169	238	170
rect	237	193	238	194
rect	239	19	240	20
rect	239	37	240	38
rect	239	67	240	68
rect	239	76	240	77
rect	239	154	240	155
rect	239	175	240	176
rect	241	16	242	17
rect	241	37	242	38
rect	241	67	242	68
rect	241	73	242	74
rect	241	136	242	137
rect	241	169	242	170
rect	241	181	242	182
rect	241	190	242	191
rect	241	277	242	278
rect	241	283	242	284
rect	241	289	242	290
rect	241	310	242	311
rect	241	334	242	335
rect	241	337	242	338
rect	243	5	244	6
rect	243	16	244	17
rect	243	22	244	23
rect	243	40	244	41
rect	243	61	244	62
rect	243	73	244	74
rect	243	103	244	104
rect	243	115	244	116
rect	243	127	244	128
rect	243	136	244	137
rect	243	154	244	155
rect	243	157	244	158
rect	243	172	244	173
rect	243	181	244	182
rect	243	205	244	206
rect	243	208	244	209
rect	243	229	244	230
rect	243	232	244	233
rect	243	262	244	263
rect	243	298	244	299
rect	243	331	244	332
rect	243	355	244	356
rect	245	13	246	14
rect	245	133	246	134
rect	245	151	246	152
rect	245	172	246	173
rect	245	202	246	203
rect	245	214	246	215
rect	245	220	246	221
rect	245	229	246	230
rect	245	253	246	254
rect	245	262	246	263
rect	245	274	246	275
rect	245	277	246	278
rect	245	280	246	281
rect	245	286	246	287
rect	245	289	246	290
rect	245	295	246	296
rect	245	322	246	323
rect	245	352	246	353
rect	247	7	248	8
rect	247	13	248	14
rect	247	31	248	32
rect	247	40	248	41
rect	247	61	248	62
rect	247	64	248	65
rect	247	100	248	101
rect	247	103	248	104
rect	247	106	248	107
rect	247	112	248	113
rect	247	124	248	125
rect	247	151	248	152
rect	247	157	248	158
rect	247	160	248	161
rect	247	196	248	197
rect	247	220	248	221
rect	247	241	248	242
rect	247	256	248	257
rect	247	268	248	269
rect	247	274	248	275
rect	247	280	248	281
rect	247	292	248	293
rect	247	319	248	320
rect	247	325	248	326
rect	247	328	248	329
rect	247	364	248	365
rect	249	1	250	2
rect	249	7	250	8
rect	249	10	250	11
rect	249	109	250	110
rect	249	121	250	122
rect	249	127	250	128
rect	249	145	250	146
rect	249	166	250	167
rect	249	178	250	179
rect	249	184	250	185
rect	249	187	250	188
rect	249	196	250	197
rect	249	199	250	200
rect	249	205	250	206
rect	249	223	250	224
rect	249	226	250	227
rect	249	238	250	239
rect	249	241	250	242
rect	249	250	250	251
rect	249	259	250	260
rect	249	265	250	266
rect	249	301	250	302
rect	249	304	250	305
rect	249	319	250	320
rect	249	322	250	323
rect	249	349	250	350
rect	251	1	252	2
rect	251	10	252	11
rect	251	28	252	29
rect	251	31	252	32
rect	251	49	252	50
rect	251	55	252	56
rect	251	58	252	59
rect	251	70	252	71
rect	251	88	252	89
rect	251	100	252	101
rect	251	112	252	113
rect	251	334	252	335
rect	260	298	261	299
rect	260	304	261	305
rect	262	286	263	287
rect	262	298	263	299
rect	264	280	265	281
rect	264	286	265	287
rect	266	226	267	227
rect	266	280	267	281
rect	268	217	269	218
rect	268	226	269	227
rect	270	193	271	194
rect	270	217	271	218
rect	272	175	273	176
rect	272	193	273	194
rect	274	58	275	59
rect	274	82	275	83
rect	274	172	275	173
rect	274	187	275	188
rect	276	79	277	80
rect	276	82	277	83
rect	276	151	277	152
rect	276	184	277	185
rect	278	28	279	29
rect	278	37	279	38
rect	278	76	279	77
rect	278	85	279	86
rect	278	136	279	137
rect	278	151	279	152
rect	278	169	279	170
rect	278	211	279	212
rect	278	262	279	263
rect	278	268	279	269
rect	278	289	279	290
rect	278	292	279	293
rect	278	310	279	311
rect	278	316	279	317
rect	280	28	281	29
rect	280	34	281	35
rect	280	70	281	71
rect	280	79	281	80
rect	280	118	281	119
rect	280	124	281	125
rect	280	136	281	137
rect	280	139	281	140
rect	280	154	281	155
rect	280	172	281	173
rect	280	175	281	176
rect	280	178	281	179
rect	280	199	281	200
rect	280	208	281	209
rect	280	259	281	260
rect	280	265	281	266
rect	280	283	281	284
rect	280	289	281	290
rect	280	307	281	308
rect	280	313	281	314
rect	282	16	283	17
rect	282	34	283	35
rect	282	67	283	68
rect	282	70	283	71
rect	282	73	283	74
rect	282	76	283	77
rect	282	115	283	116
rect	282	118	283	119
rect	282	139	283	140
rect	282	328	283	329
rect	282	352	283	353
rect	282	361	283	362
rect	284	10	285	11
rect	284	16	285	17
rect	284	22	285	23
rect	284	37	285	38
rect	284	67	285	68
rect	284	88	285	89
rect	284	94	285	95
rect	284	121	285	122
rect	284	133	285	134
rect	284	148	285	149
rect	284	154	285	155
rect	284	157	285	158
rect	284	166	285	167
rect	284	208	285	209
rect	284	235	285	236
rect	284	241	285	242
rect	284	247	285	248
rect	284	250	285	251
rect	284	253	285	254
rect	284	316	285	317
rect	284	325	285	326
rect	284	331	285	332
rect	284	334	285	335
rect	284	349	285	350
rect	284	352	285	353
rect	284	355	285	356
rect	286	10	287	11
rect	286	31	287	32
rect	286	64	287	65
rect	286	115	287	116
rect	286	130	287	131
rect	286	169	287	170
rect	286	178	287	179
rect	286	181	287	182
rect	286	232	287	233
rect	286	355	287	356
rect	288	19	289	20
rect	288	22	289	23
rect	288	31	289	32
rect	288	238	289	239
rect	288	247	289	248
rect	288	253	289	254
rect	288	256	289	257
rect	288	262	289	263
rect	288	271	289	272
rect	288	307	289	308
rect	288	319	289	320
rect	288	346	289	347
rect	290	13	291	14
rect	290	19	291	20
rect	290	55	291	56
rect	290	73	291	74
rect	290	91	291	92
rect	290	94	291	95
rect	290	127	291	128
rect	290	181	291	182
rect	290	205	291	206
rect	290	214	291	215
rect	290	229	291	230
rect	290	238	291	239
rect	290	244	291	245
rect	290	259	291	260
rect	290	271	291	272
rect	290	274	291	275
rect	290	277	291	278
rect	290	283	291	284
rect	290	301	291	302
rect	290	319	291	320
rect	290	322	291	323
rect	290	340	291	341
rect	292	7	293	8
rect	292	13	293	14
rect	292	40	293	41
rect	292	46	293	47
rect	292	49	293	50
rect	292	295	293	296
rect	292	301	293	302
rect	292	310	293	311
rect	292	322	293	323
rect	292	337	293	338
rect	301	238	302	239
rect	301	253	302	254
rect	303	226	304	227
rect	303	241	304	242
rect	305	208	306	209
rect	305	238	306	239
rect	307	196	308	197
rect	307	208	308	209
rect	307	211	308	212
rect	307	226	308	227
rect	309	193	310	194
rect	309	211	310	212
rect	311	151	312	152
rect	311	166	312	167
rect	311	175	312	176
rect	311	196	312	197
rect	313	124	314	125
rect	313	130	314	131
rect	313	148	314	149
rect	313	175	314	176
rect	313	178	314	179
rect	313	184	314	185
rect	313	187	314	188
rect	313	205	314	206
rect	315	61	316	62
rect	315	286	316	287
rect	317	118	318	119
rect	317	157	318	158
rect	317	172	318	173
rect	317	178	318	179
rect	317	181	318	182
rect	317	199	318	200
rect	317	217	318	218
rect	317	229	318	230
rect	317	268	318	269
rect	317	286	318	287
rect	317	331	318	332
rect	317	343	318	344
rect	319	106	320	107
rect	319	109	320	110
rect	319	115	320	116
rect	319	160	320	161
rect	319	169	320	170
rect	319	220	320	221
rect	319	265	320	266
rect	319	268	320	269
rect	319	316	320	317
rect	319	331	320	332
rect	321	11	322	12
rect	321	19	322	20
rect	321	106	322	107
rect	321	136	322	137
rect	321	145	322	146
rect	321	274	322	275
rect	321	280	322	281
rect	321	316	322	317
rect	323	16	324	17
rect	323	25	324	26
rect	323	79	324	80
rect	323	280	324	281
rect	323	301	324	302
rect	323	310	324	311
rect	325	16	326	17
rect	325	31	326	32
rect	325	61	326	62
rect	325	82	326	83
rect	325	97	326	98
rect	325	124	326	125
rect	325	136	326	137
rect	325	139	326	140
rect	325	148	326	149
rect	325	154	326	155
rect	325	163	326	164
rect	325	223	326	224
rect	325	235	326	236
rect	325	244	326	245
rect	325	247	326	248
rect	325	265	326	266
rect	325	271	326	272
rect	325	274	326	275
rect	325	292	326	293
rect	325	301	326	302
rect	325	307	326	308
rect	325	313	326	314
rect	325	349	326	350
rect	325	373	326	374
rect	327	13	328	14
rect	327	19	328	20
rect	327	58	328	59
rect	327	64	328	65
rect	327	73	328	74
rect	327	79	328	80
rect	327	91	328	92
rect	327	94	328	95
rect	327	97	328	98
rect	327	133	328	134
rect	327	139	328	140
rect	327	187	328	188
rect	327	190	328	191
rect	327	193	328	194
rect	327	214	328	215
rect	327	223	328	224
rect	327	232	328	233
rect	327	256	328	257
rect	327	262	328	263
rect	327	271	328	272
rect	327	283	328	284
rect	327	313	328	314
rect	327	340	328	341
rect	327	349	328	350
rect	329	13	330	14
rect	329	28	330	29
rect	329	44	330	45
rect	329	49	330	50
rect	329	58	330	59
rect	329	76	330	77
rect	329	88	330	89
rect	329	94	330	95
rect	329	115	330	116
rect	329	118	330	119
rect	329	133	330	134
rect	329	346	330	347
rect	331	11	332	12
rect	331	28	332	29
rect	331	31	332	32
rect	331	34	332	35
rect	331	46	332	47
rect	331	49	332	50
rect	331	70	332	71
rect	331	76	332	77
rect	331	82	332	83
rect	331	85	332	86
rect	331	88	332	89
rect	331	295	332	296
rect	331	319	332	320
rect	331	340	332	341
rect	331	364	332	365
rect	331	376	332	377
rect	333	22	334	23
rect	333	34	334	35
rect	333	44	334	45
rect	333	46	334	47
rect	333	67	334	68
rect	333	73	334	74
rect	333	85	334	86
rect	333	250	334	251
rect	333	259	334	260
rect	333	283	334	284
rect	333	289	334	290
rect	333	298	334	299
rect	333	304	334	305
rect	333	319	334	320
rect	333	352	334	353
rect	333	364	334	365
rect	335	22	336	23
rect	335	358	336	359
rect	335	361	336	362
rect	335	385	336	386
rect	344	233	345	234
rect	344	295	345	296
rect	346	295	347	296
rect	346	310	347	311
rect	348	86	349	87
rect	348	109	349	110
rect	348	112	349	113
rect	348	133	349	134
rect	348	233	349	234
rect	348	310	349	311
rect	350	10	351	11
rect	350	16	351	17
rect	350	109	351	110
rect	350	127	351	128
rect	350	244	351	245
rect	350	247	351	248
rect	352	16	353	17
rect	352	22	353	23
rect	352	86	353	87
rect	352	127	353	128
rect	352	133	353	134
rect	352	145	353	146
rect	352	238	353	239
rect	352	244	353	245
rect	354	19	355	20
rect	354	22	355	23
rect	354	118	355	119
rect	354	151	355	152
rect	354	238	355	239
rect	354	241	355	242
rect	356	19	357	20
rect	356	43	357	44
rect	356	82	357	83
rect	356	280	357	281
rect	358	28	359	29
rect	358	43	359	44
rect	358	115	359	116
rect	358	136	359	137
rect	358	145	359	146
rect	358	157	359	158
rect	358	241	359	242
rect	358	265	359	266
rect	358	280	359	281
rect	358	298	359	299
rect	358	319	359	320
rect	358	349	359	350
rect	360	28	361	29
rect	360	37	361	38
rect	360	88	361	89
rect	360	97	361	98
rect	360	118	361	119
rect	360	130	361	131
rect	360	136	361	137
rect	360	148	361	149
rect	360	157	361	158
rect	360	160	361	161
rect	360	265	361	266
rect	360	268	361	269
rect	360	298	361	299
rect	360	322	361	323
rect	360	355	361	356
rect	360	364	361	365
rect	360	367	361	368
rect	360	385	361	386
rect	362	4	363	5
rect	362	73	363	74
rect	362	97	363	98
rect	362	106	363	107
rect	362	130	363	131
rect	362	142	363	143
rect	362	154	363	155
rect	362	163	363	164
rect	362	175	363	176
rect	362	190	363	191
rect	362	268	363	269
rect	362	274	363	275
rect	362	292	363	293
rect	362	313	363	314
rect	362	316	363	317
rect	362	322	363	323
rect	362	364	363	365
rect	362	379	363	380
rect	364	25	365	26
rect	364	40	365	41
rect	364	64	365	65
rect	364	67	365	68
rect	364	73	365	74
rect	364	91	365	92
rect	364	106	365	107
rect	364	121	365	122
rect	364	124	365	125
rect	364	160	365	161
rect	364	163	365	164
rect	364	166	365	167
rect	364	172	365	173
rect	364	178	365	179
rect	364	187	365	188
rect	364	196	365	197
rect	364	199	365	200
rect	364	211	365	212
rect	364	218	365	219
rect	364	220	365	221
rect	364	250	365	251
rect	364	271	365	272
rect	364	277	365	278
rect	364	286	365	287
rect	364	313	365	314
rect	364	319	365	320
rect	364	325	365	326
rect	364	343	365	344
rect	364	358	365	359
rect	364	373	365	374
rect	366	25	367	26
rect	366	31	367	32
rect	366	37	367	38
rect	366	46	367	47
rect	366	58	367	59
rect	366	64	367	65
rect	366	91	367	92
rect	366	94	367	95
rect	366	121	367	122
rect	366	139	367	140
rect	366	142	367	143
rect	366	169	367	170
rect	366	178	367	179
rect	366	181	367	182
rect	366	184	367	185
rect	366	190	367	191
rect	366	208	367	209
rect	366	211	367	212
rect	366	220	367	221
rect	366	223	367	224
rect	366	226	367	227
rect	366	349	367	350
rect	366	352	367	353
rect	366	376	367	377
rect	368	31	369	32
rect	368	34	369	35
rect	368	46	369	47
rect	368	49	369	50
rect	368	55	369	56
rect	368	61	369	62
rect	368	94	369	95
rect	368	100	369	101
rect	368	103	369	104
rect	368	124	369	125
rect	368	148	369	149
rect	368	169	369	170
rect	368	175	369	176
rect	368	193	369	194
rect	368	205	369	206
rect	368	208	369	209
rect	368	218	369	219
rect	368	223	369	224
rect	368	226	369	227
rect	368	229	369	230
rect	368	235	369	236
rect	368	259	369	260
rect	368	262	369	263
rect	368	283	369	284
rect	368	289	369	290
rect	368	328	369	329
rect	368	331	369	332
rect	368	337	369	338
rect	368	340	369	341
rect	368	370	369	371
rect	377	169	378	170
rect	377	172	378	173
rect	379	172	380	173
rect	379	187	380	188
rect	381	148	382	149
rect	381	187	382	188
rect	383	148	384	149
rect	383	175	384	176
rect	383	203	384	204
rect	383	268	384	269
rect	385	163	386	164
rect	385	175	386	176
rect	385	268	386	269
rect	385	280	386	281
rect	387	157	388	158
rect	387	163	388	164
rect	387	277	388	278
rect	387	280	388	281
rect	389	154	390	155
rect	389	157	390	158
rect	389	265	390	266
rect	389	277	390	278
rect	391	145	392	146
rect	391	154	392	155
rect	391	203	392	204
rect	391	265	392	266
rect	393	124	394	125
rect	393	145	394	146
rect	393	256	394	257
rect	393	262	394	263
rect	395	100	396	101
rect	395	112	396	113
rect	395	124	396	125
rect	395	136	396	137
rect	395	247	396	248
rect	395	256	396	257
rect	397	112	398	113
rect	397	121	398	122
rect	397	127	398	128
rect	397	136	398	137
rect	397	241	398	242
rect	397	247	398	248
rect	399	97	400	98
rect	399	127	400	128
rect	399	238	400	239
rect	399	241	400	242
rect	399	250	400	251
rect	399	259	400	260
rect	401	85	402	86
rect	401	88	402	89
rect	401	97	402	98
rect	401	109	402	110
rect	401	118	402	119
rect	401	121	402	122
rect	401	223	402	224
rect	401	250	402	251
rect	403	85	404	86
rect	403	91	404	92
rect	403	109	404	110
rect	403	115	404	116
rect	403	118	404	119
rect	403	133	404	134
rect	403	160	404	161
rect	403	166	404	167
rect	403	220	404	221
rect	403	238	404	239
rect	405	25	406	26
rect	405	31	406	32
rect	405	91	406	92
rect	405	307	406	308
rect	407	25	408	26
rect	407	37	408	38
rect	407	43	408	44
rect	407	229	408	230
rect	409	22	410	23
rect	409	37	410	38
rect	409	52	410	53
rect	409	55	410	56
rect	409	64	410	65
rect	409	70	410	71
rect	409	79	410	80
rect	409	103	410	104
rect	409	115	410	116
rect	409	130	410	131
rect	409	151	410	152
rect	409	160	410	161
rect	409	211	410	212
rect	409	214	410	215
rect	409	217	410	218
rect	409	226	410	227
rect	409	229	410	230
rect	409	253	410	254
rect	409	322	410	323
rect	409	361	410	362
rect	411	10	412	11
rect	411	22	412	23
rect	411	55	412	56
rect	411	67	412	68
rect	411	73	412	74
rect	411	79	412	80
rect	411	88	412	89
rect	411	271	412	272
rect	411	286	412	287
rect	411	292	412	293
rect	411	319	412	320
rect	411	322	412	323
rect	413	10	414	11
rect	413	19	414	20
rect	413	28	414	29
rect	413	43	414	44
rect	413	46	414	47
rect	413	358	414	359
rect	415	7	416	8
rect	415	16	416	17
rect	415	19	416	20
rect	415	28	416	29
rect	415	34	416	35
rect	415	232	416	233
rect	415	244	416	245
rect	415	253	416	254
rect	415	289	416	290
rect	415	292	416	293
rect	415	313	416	314
rect	415	325	416	326
rect	417	4	418	5
rect	417	76	418	77
rect	417	82	418	83
rect	417	205	418	206
rect	417	208	418	209
rect	417	226	418	227
rect	417	235	418	236
rect	417	244	418	245
rect	417	283	418	284
rect	417	298	418	299
rect	417	310	418	311
rect	417	325	418	326
rect	419	1	420	2
rect	419	295	420	296
rect	419	310	420	311
rect	419	319	420	320
rect	419	331	420	332
rect	419	334	420	335
rect	419	349	420	350
rect	419	352	420	353
rect	428	79	429	80
rect	428	97	429	98
rect	430	76	431	77
rect	430	265	431	266
rect	432	76	433	77
rect	432	94	433	95
rect	432	235	433	236
rect	432	241	433	242
rect	434	37	435	38
rect	434	130	435	131
rect	434	154	435	155
rect	434	160	435	161
rect	434	235	435	236
rect	434	247	435	248
rect	436	22	437	23
rect	436	37	437	38
rect	436	64	437	65
rect	436	82	437	83
rect	436	106	437	107
rect	436	130	437	131
rect	436	142	437	143
rect	436	163	437	164
rect	436	244	437	245
rect	436	247	437	248
rect	438	22	439	23
rect	438	28	439	29
rect	438	73	439	74
rect	438	82	439	83
rect	438	97	439	98
rect	438	124	439	125
rect	438	145	439	146
rect	438	160	439	161
rect	438	163	439	164
rect	438	178	439	179
rect	438	238	439	239
rect	438	244	439	245
rect	438	277	439	278
rect	438	286	439	287
rect	438	298	439	299
rect	438	310	439	311
rect	440	28	441	29
rect	440	43	441	44
rect	440	67	441	68
rect	440	70	441	71
rect	440	73	441	74
rect	440	91	441	92
rect	440	94	441	95
rect	440	115	441	116
rect	440	145	441	146
rect	440	172	441	173
rect	440	178	441	179
rect	440	190	441	191
rect	440	238	441	239
rect	440	253	441	254
rect	440	286	441	287
rect	440	301	441	302
rect	440	310	441	311
rect	440	334	441	335
rect	442	43	443	44
rect	442	55	443	56
rect	442	70	443	71
rect	442	88	443	89
rect	442	91	443	92
rect	442	112	443	113
rect	442	121	443	122
rect	442	334	443	335
rect	444	4	445	5
rect	444	367	445	368
rect	446	4	447	5
rect	446	7	447	8
rect	446	40	447	41
rect	446	55	447	56
rect	446	88	447	89
rect	446	109	447	110
rect	446	112	447	113
rect	446	127	447	128
rect	446	133	447	134
rect	446	148	447	149
rect	446	175	447	176
rect	446	181	447	182
rect	446	196	447	197
rect	446	199	447	200
rect	446	217	447	218
rect	446	220	447	221
rect	446	229	447	230
rect	446	232	447	233
rect	446	250	447	251
rect	446	253	447	254
rect	446	277	447	278
rect	446	292	447	293
rect	446	301	447	302
rect	446	313	447	314
rect	446	316	447	317
rect	446	325	447	326
rect	448	7	449	8
rect	448	10	449	11
rect	448	19	449	20
rect	448	25	449	26
rect	448	31	449	32
rect	448	40	449	41
rect	448	85	449	86
rect	448	106	449	107
rect	448	109	449	110
rect	448	118	449	119
rect	448	121	449	122
rect	448	157	449	158
rect	448	166	449	167
rect	448	175	449	176
rect	448	184	449	185
rect	448	187	449	188
rect	448	190	449	191
rect	448	211	449	212
rect	448	214	449	215
rect	448	217	449	218
rect	448	226	449	227
rect	448	229	449	230
rect	448	250	449	251
rect	448	283	449	284
rect	448	295	449	296
rect	448	304	449	305
rect	448	313	449	314
rect	448	331	449	332
rect	448	346	449	347
rect	448	364	449	365
rect	450	10	451	11
rect	450	13	451	14
rect	450	25	451	26
rect	450	34	451	35
rect	450	85	451	86
rect	450	100	451	101
rect	450	103	451	104
rect	450	124	451	125
rect	450	127	451	128
rect	450	136	451	137
rect	450	157	451	158
rect	450	169	451	170
rect	450	172	451	173
rect	450	202	451	203
rect	450	214	451	215
rect	450	262	451	263
rect	450	271	451	272
rect	450	280	451	281
rect	450	289	451	290
rect	450	322	451	323
rect	450	331	451	332
rect	450	349	451	350
rect	450	355	451	356
rect	450	358	451	359
rect	459	274	460	275
rect	459	286	460	287
rect	461	286	462	287
rect	461	310	462	311
rect	463	124	464	125
rect	463	310	464	311
rect	465	124	466	125
rect	465	133	466	134
rect	465	187	466	188
rect	465	196	466	197
rect	465	226	466	227
rect	465	238	466	239
rect	467	133	468	134
rect	467	172	468	173
rect	467	196	468	197
rect	467	211	468	212
rect	467	238	468	239
rect	467	259	468	260
rect	469	46	470	47
rect	469	64	470	65
rect	469	163	470	164
rect	469	172	470	173
rect	469	211	470	212
rect	469	217	470	218
rect	469	223	470	224
rect	469	346	470	347
rect	471	64	472	65
rect	471	79	472	80
rect	471	151	472	152
rect	471	154	472	155
rect	471	163	472	164
rect	471	175	472	176
rect	471	217	472	218
rect	471	247	472	248
rect	473	58	474	59
rect	473	73	474	74
rect	473	79	474	80
rect	473	97	474	98
rect	473	100	474	101
rect	473	112	474	113
rect	473	139	474	140
rect	473	142	474	143
rect	473	151	474	152
rect	473	169	474	170
rect	473	181	474	182
rect	473	184	474	185
rect	473	214	474	215
rect	473	223	474	224
rect	473	247	474	248
rect	473	256	474	257
rect	473	259	474	260
rect	473	268	474	269
rect	473	271	474	272
rect	473	301	474	302
rect	475	55	476	56
rect	475	73	476	74
rect	475	76	476	77
rect	475	100	476	101
rect	475	115	476	116
rect	475	121	476	122
rect	475	136	476	137
rect	475	157	476	158
rect	475	175	476	176
rect	475	181	476	182
rect	475	214	476	215
rect	475	220	476	221
rect	475	256	476	257
rect	475	265	476	266
rect	475	268	476	269
rect	475	295	476	296
rect	477	55	478	56
rect	477	70	478	71
rect	477	76	478	77
rect	477	94	478	95
rect	477	121	478	122
rect	477	127	478	128
rect	477	130	478	131
rect	477	142	478	143
rect	477	169	478	170
rect	477	178	478	179
rect	477	208	478	209
rect	477	235	478	236
rect	477	244	478	245
rect	477	277	478	278
rect	477	292	478	293
rect	477	316	478	317
rect	479	37	480	38
rect	479	307	480	308
rect	481	16	482	17
rect	481	313	482	314
rect	483	16	484	17
rect	483	19	484	20
rect	483	34	484	35
rect	483	43	484	44
rect	483	49	484	50
rect	483	67	484	68
rect	483	70	484	71
rect	483	85	484	86
rect	483	106	484	107
rect	483	316	484	317
rect	485	4	486	5
rect	485	7	486	8
rect	485	19	486	20
rect	485	22	486	23
rect	485	31	486	32
rect	485	40	486	41
rect	485	52	486	53
rect	485	61	486	62
rect	485	67	486	68
rect	485	82	486	83
rect	485	103	486	104
rect	485	109	486	110
rect	485	112	486	113
rect	485	145	486	146
rect	485	154	486	155
rect	485	160	486	161
rect	485	166	486	167
rect	485	193	486	194
rect	485	205	486	206
rect	485	232	486	233
rect	485	235	486	236
rect	485	250	486	251
rect	485	253	486	254
rect	485	343	486	344
rect	487	7	488	8
rect	487	10	488	11
rect	487	22	488	23
rect	487	25	488	26
rect	487	28	488	29
rect	487	37	488	38
rect	487	52	488	53
rect	487	280	488	281
rect	487	283	488	284
rect	487	298	488	299
rect	487	307	488	308
rect	487	331	488	332
rect	496	160	497	161
rect	496	163	497	164
rect	498	4	499	5
rect	498	208	499	209
rect	500	163	501	164
rect	500	196	501	197
rect	500	199	501	200
rect	500	208	501	209
rect	502	196	503	197
rect	502	211	503	212
rect	504	190	505	191
rect	504	235	505	236
rect	504	277	505	278
rect	504	283	505	284
rect	506	28	507	29
rect	506	49	507	50
rect	506	181	507	182
rect	506	277	507	278
rect	508	25	509	26
rect	508	46	509	47
rect	508	49	509	50
rect	508	67	509	68
rect	508	145	509	146
rect	508	151	509	152
rect	508	178	509	179
rect	508	226	509	227
rect	508	238	509	239
rect	508	247	509	248
rect	510	46	511	47
rect	510	64	511	65
rect	510	151	511	152
rect	510	166	511	167
rect	510	175	511	176
rect	510	205	511	206
rect	510	238	511	239
rect	510	271	511	272
rect	512	43	513	44
rect	512	61	513	62
rect	512	85	513	86
rect	512	88	513	89
rect	512	166	513	167
rect	512	169	513	170
rect	512	172	513	173
rect	512	181	513	182
rect	512	184	513	185
rect	512	202	513	203
rect	512	211	513	212
rect	512	244	513	245
rect	512	247	513	248
rect	512	274	513	275
rect	514	40	515	41
rect	514	58	515	59
rect	514	82	515	83
rect	514	100	515	101
rect	514	130	515	131
rect	514	139	515	140
rect	514	148	515	149
rect	514	154	515	155
rect	514	169	515	170
rect	514	187	515	188
rect	514	193	515	194
rect	514	223	515	224
rect	514	235	515	236
rect	514	256	515	257
rect	516	34	517	35
rect	516	64	517	65
rect	516	73	517	74
rect	516	106	517	107
rect	516	130	517	131
rect	516	268	517	269
rect	518	13	519	14
rect	518	19	519	20
rect	518	34	519	35
rect	518	52	519	53
rect	518	61	519	62
rect	518	70	519	71
rect	518	73	519	74
rect	518	79	519	80
rect	518	88	519	89
rect	518	91	519	92
rect	518	100	519	101
rect	518	112	519	113
rect	518	118	519	119
rect	518	136	519	137
rect	518	142	519	143
rect	518	250	519	251
rect	520	1	521	2
rect	520	7	521	8
rect	520	13	521	14
rect	520	22	521	23
rect	520	37	521	38
rect	520	52	521	53
rect	520	70	521	71
rect	520	241	521	242
rect	520	274	521	275
rect	520	307	521	308
rect	522	7	523	8
rect	522	16	523	17
rect	522	37	523	38
rect	522	55	523	56
rect	522	67	523	68
rect	522	76	523	77
rect	522	91	523	92
rect	522	103	523	104
rect	522	115	523	116
rect	522	133	523	134
rect	522	139	523	140
rect	522	253	523	254
rect	522	256	523	257
rect	522	259	523	260
rect	522	265	523	266
rect	522	292	523	293
rect	531	154	532	155
rect	531	160	532	161
rect	533	160	534	161
rect	533	166	534	167
rect	535	25	536	26
rect	535	28	536	29
rect	535	31	536	32
rect	535	55	536	56
rect	535	157	536	158
rect	535	163	536	164
rect	535	166	536	167
rect	535	181	536	182
rect	537	28	538	29
rect	537	52	538	53
rect	537	55	538	56
rect	537	64	538	65
rect	537	79	538	80
rect	537	85	538	86
rect	537	133	538	134
rect	537	151	538	152
rect	537	163	538	164
rect	537	178	538	179
rect	537	184	538	185
rect	537	199	538	200
rect	537	202	538	203
rect	537	208	538	209
rect	537	232	538	233
rect	537	247	538	248
rect	539	52	540	53
rect	539	61	540	62
rect	539	64	540	65
rect	539	73	540	74
rect	539	76	540	77
rect	539	100	540	101
rect	539	112	540	113
rect	539	121	540	122
rect	539	151	540	152
rect	539	175	540	176
rect	539	178	540	179
rect	539	193	540	194
rect	539	202	540	203
rect	539	211	540	212
rect	539	229	540	230
rect	539	238	540	239
rect	541	61	542	62
rect	541	70	542	71
rect	541	73	542	74
rect	541	82	542	83
rect	541	85	542	86
rect	541	91	542	92
rect	541	109	542	110
rect	541	118	542	119
rect	541	127	542	128
rect	541	241	542	242
rect	543	10	544	11
rect	543	181	544	182
rect	543	196	544	197
rect	543	199	544	200
rect	543	211	544	212
rect	543	214	544	215
rect	543	220	544	221
rect	543	235	544	236
rect	543	247	544	248
rect	543	256	544	257
rect	543	259	544	260
rect	543	274	544	275
rect	545	7	546	8
rect	545	13	546	14
rect	545	25	546	26
rect	545	34	546	35
rect	545	58	546	59
rect	545	67	546	68
rect	545	82	546	83
rect	545	88	546	89
rect	545	100	546	101
rect	545	115	546	116
rect	545	121	546	122
rect	545	139	546	140
rect	545	142	546	143
rect	545	148	546	149
rect	545	175	546	176
rect	545	190	546	191
rect	545	196	546	197
rect	545	244	546	245
rect	545	256	546	257
rect	545	265	546	266
rect	554	34	555	35
rect	554	46	555	47
rect	554	151	555	152
rect	554	169	555	170
rect	556	31	557	32
rect	556	37	557	38
rect	556	55	557	56
rect	556	70	557	71
rect	556	166	557	167
rect	556	169	557	170
rect	558	31	559	32
rect	558	43	559	44
rect	558	55	559	56
rect	558	64	559	65
rect	558	163	559	164
rect	558	166	559	167
rect	560	28	561	29
rect	560	43	561	44
rect	560	64	561	65
rect	560	73	561	74
rect	560	148	561	149
rect	560	157	561	158
rect	560	163	561	164
rect	560	184	561	185
rect	560	199	561	200
rect	560	205	561	206
rect	562	28	563	29
rect	562	40	563	41
rect	562	46	563	47
rect	562	235	563	236
rect	562	241	563	242
rect	562	250	563	251
rect	564	40	565	41
rect	564	52	565	53
rect	564	73	565	74
rect	564	79	565	80
rect	564	157	565	158
rect	564	178	565	179
rect	564	196	565	197
rect	564	211	565	212
rect	564	217	565	218
rect	564	229	565	230
rect	564	247	565	248
rect	564	250	565	251
rect	566	37	567	38
rect	566	49	567	50
rect	566	52	567	53
rect	566	61	567	62
rect	566	67	567	68
rect	566	76	567	77
rect	566	79	567	80
rect	566	85	567	86
rect	566	106	567	107
rect	566	112	567	113
rect	566	118	567	119
rect	566	121	567	122
rect	566	154	567	155
rect	566	172	567	173
rect	566	196	567	197
rect	566	202	567	203
rect	566	214	567	215
rect	566	223	567	224
rect	566	229	567	230
rect	566	244	567	245
rect	566	247	567	248
rect	566	259	567	260
rect	568	7	569	8
rect	568	13	569	14
rect	568	22	569	23
rect	568	25	569	26
rect	568	49	569	50
rect	568	58	569	59
rect	568	76	569	77
rect	568	82	569	83
rect	568	94	569	95
rect	568	100	569	101
rect	568	103	569	104
rect	568	109	569	110
rect	568	115	569	116
rect	568	133	569	134
rect	568	142	569	143
rect	568	145	569	146
rect	568	154	569	155
rect	568	175	569	176
rect	568	181	569	182
rect	568	184	569	185
rect	568	193	569	194
rect	568	220	569	221
rect	568	226	569	227
rect	568	232	569	233
rect	568	235	569	236
rect	568	238	569	239
rect	568	244	569	245
rect	568	256	569	257
rect	577	22	578	23
rect	577	28	578	29
rect	579	22	580	23
rect	579	40	580	41
rect	581	37	582	38
rect	581	40	582	41
rect	583	31	584	32
rect	583	37	584	38
rect	585	31	586	32
rect	585	55	586	56
rect	587	25	588	26
rect	587	43	588	44
rect	587	55	588	56
rect	587	67	588	68
rect	589	43	590	44
rect	589	46	590	47
rect	589	61	590	62
rect	589	64	590	65
rect	589	67	590	68
rect	589	79	590	80
rect	589	205	590	206
rect	589	208	590	209
rect	591	46	592	47
rect	591	52	592	53
rect	591	64	592	65
rect	591	76	592	77
rect	591	97	592	98
rect	591	103	592	104
rect	591	151	592	152
rect	591	154	592	155
rect	591	169	592	170
rect	591	175	592	176
rect	591	202	592	203
rect	591	217	592	218
rect	591	223	592	224
rect	591	238	592	239
rect	593	28	594	29
rect	593	49	594	50
rect	593	61	594	62
rect	593	73	594	74
rect	593	103	594	104
rect	593	115	594	116
rect	593	142	594	143
rect	593	157	594	158
rect	593	169	594	170
rect	593	193	594	194
rect	593	199	594	200
rect	593	205	594	206
rect	593	211	594	212
rect	593	229	594	230
rect	595	34	596	35
rect	595	49	596	50
rect	595	58	596	59
rect	595	70	596	71
rect	595	88	596	89
rect	595	94	596	95
rect	595	100	596	101
rect	595	106	596	107
rect	595	109	596	110
rect	595	118	596	119
rect	595	133	596	134
rect	595	145	596	146
rect	595	151	596	152
rect	595	163	596	164
rect	595	166	596	167
rect	595	172	596	173
rect	595	193	596	194
rect	595	214	596	215
rect	595	220	596	221
rect	595	226	596	227
rect	595	238	596	239
rect	595	247	596	248
rect	595	250	596	251
rect	595	256	596	257
rect	604	19	605	20
rect	604	22	605	23
rect	604	37	605	38
rect	604	43	605	44
rect	604	49	605	50
rect	604	58	605	59
rect	604	164	605	165
rect	604	175	605	176
rect	604	178	605	179
rect	604	196	605	197
rect	604	199	605	200
rect	604	211	605	212
rect	606	22	607	23
rect	606	25	607	26
rect	606	43	607	44
rect	606	55	607	56
rect	606	58	607	59
rect	606	67	607	68
rect	606	85	607	86
rect	606	88	607	89
rect	606	97	607	98
rect	606	106	607	107
rect	606	175	607	176
rect	606	184	607	185
rect	606	196	607	197
rect	606	205	607	206
rect	608	7	609	8
rect	608	10	609	11
rect	608	25	609	26
rect	608	28	609	29
rect	608	34	609	35
rect	608	40	609	41
rect	608	55	609	56
rect	608	64	609	65
rect	608	82	609	83
rect	608	103	609	104
rect	608	136	609	137
rect	608	142	609	143
rect	608	164	609	165
rect	608	184	609	185
rect	608	193	609	194
rect	608	202	609	203
rect	608	208	609	209
rect	608	211	609	212
rect	608	220	609	221
rect	608	226	609	227
rect	610	10	611	11
rect	610	13	611	14
rect	610	28	611	29
rect	610	31	611	32
rect	610	40	611	41
rect	610	46	611	47
rect	610	52	611	53
rect	610	61	611	62
rect	610	79	611	80
rect	610	100	611	101
rect	610	118	611	119
rect	610	124	611	125
rect	610	127	611	128
rect	610	133	611	134
rect	610	142	611	143
rect	610	151	611	152
rect	610	157	611	158
rect	610	160	611	161
rect	610	166	611	167
rect	610	169	611	170
rect	610	172	611	173
rect	610	181	611	182
rect	610	193	611	194
rect	610	223	611	224
rect	619	175	620	176
rect	619	190	620	191
rect	621	7	622	8
rect	621	13	622	14
rect	621	16	622	17
rect	621	28	622	29
rect	621	46	622	47
rect	621	52	622	53
rect	621	175	622	176
rect	621	184	622	185
rect	621	187	622	188
rect	621	193	622	194
rect	623	13	624	14
rect	623	25	624	26
rect	623	28	624	29
rect	623	40	624	41
rect	623	46	624	47
rect	623	58	624	59
rect	623	61	624	62
rect	623	79	624	80
rect	623	172	624	173
rect	623	181	624	182
rect	623	187	624	188
rect	623	196	624	197
rect	625	25	626	26
rect	625	37	626	38
rect	625	43	626	44
rect	625	55	626	56
rect	625	79	626	80
rect	625	85	626	86
rect	625	169	626	170
rect	625	178	626	179
rect	625	196	626	197
rect	625	202	626	203
rect	625	211	626	212
rect	625	217	626	218
rect	627	7	628	8
rect	627	8	628	9
rect	627	9	628	10
rect	627	11	628	12
rect	627	12	628	13
rect	627	14	628	15
rect	627	15	628	16
rect	627	17	628	18
rect	627	18	628	19
rect	627	19	628	20
rect	627	22	628	23
rect	627	34	628	35
rect	627	40	628	41
rect	627	49	628	50
rect	627	64	628	65
rect	627	82	628	83
rect	627	88	628	89
rect	627	103	628	104
rect	627	109	628	110
rect	627	127	628	128
rect	627	133	628	134
rect	627	142	628	143
rect	627	148	628	149
rect	627	157	628	158
rect	627	163	628	164
rect	627	178	628	179
rect	627	184	628	185
rect	627	199	628	200
rect	627	217	628	218
rect	627	238	628	239
rect	636	160	637	161
rect	636	166	637	167
rect	636	175	637	176
rect	636	178	637	179
rect	638	157	639	158
rect	638	196	639	197
rect	640	55	641	56
rect	640	79	641	80
rect	640	157	641	158
rect	640	187	641	188
rect	642	52	643	53
rect	642	217	643	218
rect	644	10	645	11
rect	644	16	645	17
rect	644	22	645	23
rect	644	28	645	29
rect	644	37	645	38
rect	644	46	645	47
rect	644	49	645	50
rect	644	64	645	65
rect	644	109	645	110
rect	644	115	645	116
rect	644	139	645	140
rect	644	148	645	149
rect	644	151	645	152
rect	644	163	645	164
rect	644	172	645	173
rect	644	175	645	176
rect	646	7	647	8
rect	646	13	647	14
rect	646	19	647	20
rect	646	25	647	26
rect	646	40	647	41
rect	646	43	647	44
rect	646	46	647	47
rect	646	61	647	62
rect	646	79	647	80
rect	646	82	647	83
rect	646	85	647	86
rect	646	88	647	89
rect	646	115	647	116
rect	646	118	647	119
rect	646	124	647	125
rect	646	133	647	134
rect	646	148	647	149
rect	646	184	647	185
rect	655	148	656	149
rect	655	154	656	155
rect	657	4	658	5
rect	657	7	658	8
rect	657	13	658	14
rect	657	19	658	20
rect	657	31	658	32
rect	657	49	658	50
rect	657	136	658	137
rect	657	151	658	152
rect	659	7	660	8
rect	659	10	660	11
rect	659	13	660	14
rect	659	22	660	23
rect	659	28	660	29
rect	659	37	660	38
rect	659	43	660	44
rect	659	46	660	47
rect	659	64	660	65
rect	659	82	660	83
rect	659	85	660	86
rect	659	160	660	161
rect	659	166	660	167
rect	659	169	660	170
rect	668	88	669	89
rect	668	115	669	116
rect	668	124	669	125
rect	668	130	669	131
rect	668	139	669	140
rect	668	142	669	143
rect	670	4	671	5
rect	670	7	671	8
rect	670	25	671	26
rect	670	28	671	29
rect	670	82	671	83
rect	670	166	671	167
