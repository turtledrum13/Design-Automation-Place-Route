magic
tech scmos
timestamp
<< pdiffusion >>
rect	0	9	6	15
rect	0	45	6	51
rect	17	9	23	15
rect	56	45	62	51
rect	0	27	6	33
rect	0	63	6	69
rect	29	27	35	33
rect	20	63	26	69
rect	10	9	16	15
rect	31	45	37	51
rect	27	9	33	15
rect	78	45	84	51
rect	13	27	19	33
rect	10	63	16	69
rect	54	27	60	33
rect	27	63	33	69
rect	0	18	6	24
rect	0	54	6	60
rect	17	18	23	24
rect	35	54	41	60
rect	0	36	6	42
rect	3	72	9	78
rect	35	36	41	42
rect	37	9	43	15
rect	94	45	100	51
rect	60	9	66	15
rect	123	45	129	51
rect	82	27	88	33
rect	37	63	43	69
rect	105	27	111	33
rect	51	63	57	69
rect	47	9	53	15
rect	107	45	113	51
rect	73	9	79	15
rect	130	45	136	51
rect	95	27	101	33
rect	44	63	50	69
rect	112	27	118	33
rect	67	63	73	69
rect	46	18	52	24
rect	82	54	88	60
rect	75	18	81	24
rect	105	54	111	60
rect	67	36	73	42
rect	31	72	37	78
rect	65	18	68	24
rect	6	27	9	33
rect	23	18	26	24
rect	111	54	114	60
rect	6	9	9	15
rect	9	27	12	33
rect	55	54	58	60
rect	41	54	44	60
rect	66	9	69	15
rect	57	63	60	69
rect	53	9	56	15
rect	113	45	116	51
rect	101	54	104	60
rect	31	18	34	24
rect	41	36	44	42
rect	60	27	63	33
rect	116	45	119	51
rect	6	45	9	51
rect	19	27	22	33
rect	23	9	26	15
rect	44	36	47	42
rect	16	63	19	69
rect	88	27	91	33
rect	127	36	130	42
rect	26	18	29	24
rect	14	54	17	60
rect	34	18	37	24
rect	37	45	40	51
rect	33	9	36	15
rect	59	54	62	60
rect	28	54	31	60
rect	100	45	103	51
rect	40	45	43	51
rect	0	72	3	78
rect	69	54	72	60
rect	62	54	65	60
rect	9	45	12	51
rect	33	63	36	69
rect	31	54	34	60
rect	56	9	59	15
rect	6	63	9	69
rect	91	27	94	33
rect	63	27	66	33
rect	66	27	69	33
rect	10	36	13	42
rect	22	27	25	33
rect	136	45	139	51
rect	7	18	10	24
rect	13	36	16	42
rect	62	45	65	51
rect	65	45	68	51
rect	68	18	71	24
rect	88	54	91	60
rect	93	54	96	60
rect	119	45	122	51
rect	35	27	38	33
rect	73	36	76	42
rect	117	36	120	42
rect	7	54	10	60
rect	38	27	41	33
rect	23	54	26	60
rect	107	36	110	42
rect	41	27	44	33
rect	12	45	15	51
rect	44	27	47	33
rect	84	45	87	51
rect	15	45	18	51
rect	72	54	75	60
rect	87	45	90	51
rect	16	36	19	42
rect	44	54	47	60
rect	43	45	46	51
rect	60	18	63	24
rect	10	54	13	60
rect	113	36	116	42
rect	88	36	91	42
rect	91	36	94	42
rect	18	45	21	51
rect	47	36	50	42
rect	140	36	143	42
rect	21	45	24	51
rect	76	36	79	42
rect	69	27	72	33
rect	90	45	93	51
rect	91	63	94	69
rect	123	36	126	42
rect	101	27	104	33
rect	24	45	27	51
rect	57	36	60	42
rect	19	36	22	42
rect	79	36	82	42
rect	6	36	9	42
rect	60	63	63	69
rect	46	45	49	51
rect	50	36	53	42
rect	72	27	75	33
rect	27	45	30	51
rect	103	45	106	51
rect	68	45	71	51
rect	71	45	74	51
rect	19	54	22	60
rect	49	45	52	51
rect	75	27	78	33
rect	82	36	85	42
rect	94	36	97	42
rect	127	27	130	33
rect	102	18	105	24
rect	25	36	28	42
rect	52	45	55	51
rect	25	27	28	33
rect	53	36	56	42
rect	78	27	81	33
rect	28	36	31	42
rect	75	54	78	60
rect	78	54	81	60
rect	50	54	53	60
rect	71	18	74	24
rect	74	45	77	51
rect	131	18	134	24
rect	47	27	50	33
rect	82	18	85	24
rect	50	27	53	33
rect	76	63	79	69
rect	79	63	82	69
rect	69	9	72	15
rect	65	54	68	60
rect	52	18	55	24
rect	42	18	45	24
rect	77	72	80	78
rect	63	63	66	69
rect	43	9	46	15
