magic
tech scmos
timestamp
<< pdiffusion >>
rect	0	6	1	7
rect	1	6	2	7
rect	2	6	3	7
rect	3	6	4	7
rect	4	6	5	7
rect	5	6	6	7
rect	7	6	8	7
rect	8	6	9	7
rect	9	6	10	7
rect	10	6	11	7
rect	11	6	12	7
rect	12	6	13	7
rect	14	6	15	7
rect	15	6	16	7
rect	16	6	17	7
rect	17	6	18	7
rect	18	6	19	7
rect	19	6	20	7
rect	21	6	22	7
rect	22	6	23	7
rect	23	6	24	7
rect	24	6	25	7
rect	25	6	26	7
rect	26	6	27	7
rect	28	6	29	7
rect	29	6	30	7
rect	30	6	31	7
rect	31	6	32	7
rect	32	6	33	7
rect	33	6	34	7
rect	35	6	36	7
rect	36	6	37	7
rect	37	6	38	7
rect	38	6	39	7
rect	39	6	40	7
rect	40	6	41	7
rect	42	6	43	7
rect	43	6	44	7
rect	44	6	45	7
rect	45	6	46	7
rect	46	6	47	7
rect	47	6	48	7
rect	49	6	50	7
rect	50	6	51	7
rect	51	6	52	7
rect	52	6	53	7
rect	53	6	54	7
rect	54	6	55	7
rect	55	6	56	7
rect	56	6	57	7
rect	57	6	58	7
rect	58	6	59	7
rect	59	6	60	7
rect	60	6	61	7
rect	61	6	62	7
rect	62	6	63	7
rect	63	6	64	7
rect	65	6	66	7
rect	66	6	67	7
rect	67	6	68	7
rect	68	6	69	7
rect	69	6	70	7
rect	70	6	71	7
rect	71	6	72	7
rect	72	6	73	7
rect	73	6	74	7
rect	74	6	75	7
rect	75	6	76	7
rect	76	6	77	7
rect	77	6	78	7
rect	78	6	79	7
rect	79	6	80	7
rect	81	6	82	7
rect	82	6	83	7
rect	83	6	84	7
rect	84	6	85	7
rect	85	6	86	7
rect	86	6	87	7
rect	88	6	89	7
rect	89	6	90	7
rect	90	6	91	7
rect	91	6	92	7
rect	92	6	93	7
rect	93	6	94	7
rect	95	6	96	7
rect	96	6	97	7
rect	97	6	98	7
rect	98	6	99	7
rect	99	6	100	7
rect	100	6	101	7
rect	102	6	103	7
rect	103	6	104	7
rect	104	6	105	7
rect	105	6	106	7
rect	106	6	107	7
rect	107	6	108	7
rect	108	6	109	7
rect	109	6	110	7
rect	110	6	111	7
rect	111	6	112	7
rect	112	6	113	7
rect	113	6	114	7
rect	114	6	115	7
rect	115	6	116	7
rect	116	6	117	7
rect	117	6	118	7
rect	118	6	119	7
rect	119	6	120	7
rect	120	6	121	7
rect	121	6	122	7
rect	122	6	123	7
rect	123	6	124	7
rect	124	6	125	7
rect	125	6	126	7
rect	127	6	128	7
rect	128	6	129	7
rect	129	6	130	7
rect	130	6	131	7
rect	131	6	132	7
rect	132	6	133	7
rect	134	6	135	7
rect	135	6	136	7
rect	136	6	137	7
rect	137	6	138	7
rect	138	6	139	7
rect	139	6	140	7
rect	141	6	142	7
rect	142	6	143	7
rect	143	6	144	7
rect	144	6	145	7
rect	145	6	146	7
rect	146	6	147	7
rect	148	6	149	7
rect	149	6	150	7
rect	150	6	151	7
rect	151	6	152	7
rect	152	6	153	7
rect	153	6	154	7
rect	155	6	156	7
rect	156	6	157	7
rect	157	6	158	7
rect	158	6	159	7
rect	159	6	160	7
rect	160	6	161	7
rect	162	6	163	7
rect	163	6	164	7
rect	164	6	165	7
rect	165	6	166	7
rect	166	6	167	7
rect	167	6	168	7
rect	169	6	170	7
rect	170	6	171	7
rect	171	6	172	7
rect	172	6	173	7
rect	173	6	174	7
rect	174	6	175	7
rect	176	6	177	7
rect	177	6	178	7
rect	178	6	179	7
rect	179	6	180	7
rect	180	6	181	7
rect	181	6	182	7
rect	183	6	184	7
rect	184	6	185	7
rect	185	6	186	7
rect	186	6	187	7
rect	187	6	188	7
rect	188	6	189	7
rect	189	6	190	7
rect	190	6	191	7
rect	191	6	192	7
rect	192	6	193	7
rect	193	6	194	7
rect	194	6	195	7
rect	195	6	196	7
rect	196	6	197	7
rect	197	6	198	7
rect	199	6	200	7
rect	200	6	201	7
rect	201	6	202	7
rect	202	6	203	7
rect	203	6	204	7
rect	204	6	205	7
rect	206	6	207	7
rect	207	6	208	7
rect	208	6	209	7
rect	209	6	210	7
rect	210	6	211	7
rect	211	6	212	7
rect	213	6	214	7
rect	214	6	215	7
rect	215	6	216	7
rect	216	6	217	7
rect	217	6	218	7
rect	218	6	219	7
rect	219	6	220	7
rect	220	6	221	7
rect	221	6	222	7
rect	222	6	223	7
rect	223	6	224	7
rect	224	6	225	7
rect	225	6	226	7
rect	226	6	227	7
rect	227	6	228	7
rect	229	6	230	7
rect	230	6	231	7
rect	231	6	232	7
rect	232	6	233	7
rect	233	6	234	7
rect	234	6	235	7
rect	236	6	237	7
rect	237	6	238	7
rect	238	6	239	7
rect	239	6	240	7
rect	240	6	241	7
rect	241	6	242	7
rect	242	6	243	7
rect	243	6	244	7
rect	244	6	245	7
rect	245	6	246	7
rect	246	6	247	7
rect	247	6	248	7
rect	248	6	249	7
rect	249	6	250	7
rect	250	6	251	7
rect	251	6	252	7
rect	252	6	253	7
rect	253	6	254	7
rect	255	6	256	7
rect	256	6	257	7
rect	257	6	258	7
rect	258	6	259	7
rect	259	6	260	7
rect	260	6	261	7
rect	261	6	262	7
rect	262	6	263	7
rect	263	6	264	7
rect	264	6	265	7
rect	265	6	266	7
rect	266	6	267	7
rect	267	6	268	7
rect	268	6	269	7
rect	269	6	270	7
rect	0	7	1	8
rect	1	7	2	8
rect	2	7	3	8
rect	3	7	4	8
rect	4	7	5	8
rect	5	7	6	8
rect	7	7	8	8
rect	8	7	9	8
rect	9	7	10	8
rect	10	7	11	8
rect	11	7	12	8
rect	12	7	13	8
rect	14	7	15	8
rect	15	7	16	8
rect	16	7	17	8
rect	17	7	18	8
rect	18	7	19	8
rect	19	7	20	8
rect	21	7	22	8
rect	22	7	23	8
rect	23	7	24	8
rect	24	7	25	8
rect	25	7	26	8
rect	26	7	27	8
rect	28	7	29	8
rect	29	7	30	8
rect	30	7	31	8
rect	31	7	32	8
rect	32	7	33	8
rect	33	7	34	8
rect	35	7	36	8
rect	36	7	37	8
rect	37	7	38	8
rect	38	7	39	8
rect	39	7	40	8
rect	40	7	41	8
rect	42	7	43	8
rect	43	7	44	8
rect	44	7	45	8
rect	45	7	46	8
rect	46	7	47	8
rect	47	7	48	8
rect	49	7	50	8
rect	50	7	51	8
rect	51	7	52	8
rect	52	7	53	8
rect	53	7	54	8
rect	54	7	55	8
rect	55	7	56	8
rect	56	7	57	8
rect	57	7	58	8
rect	58	7	59	8
rect	59	7	60	8
rect	60	7	61	8
rect	61	7	62	8
rect	62	7	63	8
rect	63	7	64	8
rect	65	7	66	8
rect	66	7	67	8
rect	67	7	68	8
rect	68	7	69	8
rect	69	7	70	8
rect	70	7	71	8
rect	71	7	72	8
rect	72	7	73	8
rect	73	7	74	8
rect	74	7	75	8
rect	75	7	76	8
rect	76	7	77	8
rect	77	7	78	8
rect	78	7	79	8
rect	79	7	80	8
rect	81	7	82	8
rect	82	7	83	8
rect	83	7	84	8
rect	84	7	85	8
rect	85	7	86	8
rect	86	7	87	8
rect	88	7	89	8
rect	89	7	90	8
rect	90	7	91	8
rect	91	7	92	8
rect	92	7	93	8
rect	93	7	94	8
rect	95	7	96	8
rect	96	7	97	8
rect	97	7	98	8
rect	98	7	99	8
rect	99	7	100	8
rect	100	7	101	8
rect	102	7	103	8
rect	103	7	104	8
rect	104	7	105	8
rect	105	7	106	8
rect	106	7	107	8
rect	107	7	108	8
rect	108	7	109	8
rect	109	7	110	8
rect	110	7	111	8
rect	111	7	112	8
rect	112	7	113	8
rect	113	7	114	8
rect	114	7	115	8
rect	115	7	116	8
rect	116	7	117	8
rect	117	7	118	8
rect	118	7	119	8
rect	119	7	120	8
rect	120	7	121	8
rect	121	7	122	8
rect	122	7	123	8
rect	123	7	124	8
rect	124	7	125	8
rect	125	7	126	8
rect	127	7	128	8
rect	128	7	129	8
rect	129	7	130	8
rect	130	7	131	8
rect	131	7	132	8
rect	132	7	133	8
rect	134	7	135	8
rect	135	7	136	8
rect	136	7	137	8
rect	137	7	138	8
rect	138	7	139	8
rect	139	7	140	8
rect	141	7	142	8
rect	142	7	143	8
rect	143	7	144	8
rect	144	7	145	8
rect	145	7	146	8
rect	146	7	147	8
rect	148	7	149	8
rect	149	7	150	8
rect	150	7	151	8
rect	151	7	152	8
rect	152	7	153	8
rect	153	7	154	8
rect	155	7	156	8
rect	156	7	157	8
rect	157	7	158	8
rect	158	7	159	8
rect	159	7	160	8
rect	160	7	161	8
rect	162	7	163	8
rect	163	7	164	8
rect	164	7	165	8
rect	165	7	166	8
rect	166	7	167	8
rect	167	7	168	8
rect	169	7	170	8
rect	170	7	171	8
rect	171	7	172	8
rect	172	7	173	8
rect	173	7	174	8
rect	174	7	175	8
rect	176	7	177	8
rect	177	7	178	8
rect	178	7	179	8
rect	179	7	180	8
rect	180	7	181	8
rect	181	7	182	8
rect	183	7	184	8
rect	184	7	185	8
rect	185	7	186	8
rect	186	7	187	8
rect	187	7	188	8
rect	188	7	189	8
rect	189	7	190	8
rect	190	7	191	8
rect	191	7	192	8
rect	192	7	193	8
rect	193	7	194	8
rect	194	7	195	8
rect	195	7	196	8
rect	196	7	197	8
rect	197	7	198	8
rect	199	7	200	8
rect	200	7	201	8
rect	201	7	202	8
rect	202	7	203	8
rect	203	7	204	8
rect	204	7	205	8
rect	206	7	207	8
rect	207	7	208	8
rect	208	7	209	8
rect	209	7	210	8
rect	210	7	211	8
rect	211	7	212	8
rect	213	7	214	8
rect	214	7	215	8
rect	215	7	216	8
rect	216	7	217	8
rect	217	7	218	8
rect	218	7	219	8
rect	219	7	220	8
rect	220	7	221	8
rect	221	7	222	8
rect	222	7	223	8
rect	223	7	224	8
rect	224	7	225	8
rect	225	7	226	8
rect	226	7	227	8
rect	227	7	228	8
rect	229	7	230	8
rect	230	7	231	8
rect	231	7	232	8
rect	232	7	233	8
rect	233	7	234	8
rect	234	7	235	8
rect	236	7	237	8
rect	237	7	238	8
rect	238	7	239	8
rect	239	7	240	8
rect	240	7	241	8
rect	241	7	242	8
rect	242	7	243	8
rect	243	7	244	8
rect	244	7	245	8
rect	245	7	246	8
rect	246	7	247	8
rect	247	7	248	8
rect	248	7	249	8
rect	249	7	250	8
rect	250	7	251	8
rect	251	7	252	8
rect	252	7	253	8
rect	253	7	254	8
rect	255	7	256	8
rect	256	7	257	8
rect	257	7	258	8
rect	258	7	259	8
rect	259	7	260	8
rect	260	7	261	8
rect	261	7	262	8
rect	262	7	263	8
rect	263	7	264	8
rect	264	7	265	8
rect	265	7	266	8
rect	266	7	267	8
rect	267	7	268	8
rect	268	7	269	8
rect	269	7	270	8
rect	0	8	1	9
rect	1	8	2	9
rect	2	8	3	9
rect	3	8	4	9
rect	4	8	5	9
rect	5	8	6	9
rect	7	8	8	9
rect	8	8	9	9
rect	9	8	10	9
rect	10	8	11	9
rect	11	8	12	9
rect	12	8	13	9
rect	14	8	15	9
rect	15	8	16	9
rect	16	8	17	9
rect	17	8	18	9
rect	18	8	19	9
rect	19	8	20	9
rect	21	8	22	9
rect	22	8	23	9
rect	23	8	24	9
rect	24	8	25	9
rect	25	8	26	9
rect	26	8	27	9
rect	28	8	29	9
rect	29	8	30	9
rect	30	8	31	9
rect	31	8	32	9
rect	32	8	33	9
rect	33	8	34	9
rect	35	8	36	9
rect	36	8	37	9
rect	37	8	38	9
rect	38	8	39	9
rect	39	8	40	9
rect	40	8	41	9
rect	42	8	43	9
rect	43	8	44	9
rect	44	8	45	9
rect	45	8	46	9
rect	46	8	47	9
rect	47	8	48	9
rect	49	8	50	9
rect	50	8	51	9
rect	51	8	52	9
rect	52	8	53	9
rect	53	8	54	9
rect	54	8	55	9
rect	55	8	56	9
rect	56	8	57	9
rect	57	8	58	9
rect	58	8	59	9
rect	59	8	60	9
rect	60	8	61	9
rect	61	8	62	9
rect	62	8	63	9
rect	63	8	64	9
rect	65	8	66	9
rect	66	8	67	9
rect	67	8	68	9
rect	68	8	69	9
rect	69	8	70	9
rect	70	8	71	9
rect	71	8	72	9
rect	72	8	73	9
rect	73	8	74	9
rect	74	8	75	9
rect	75	8	76	9
rect	76	8	77	9
rect	77	8	78	9
rect	78	8	79	9
rect	79	8	80	9
rect	81	8	82	9
rect	82	8	83	9
rect	83	8	84	9
rect	84	8	85	9
rect	85	8	86	9
rect	86	8	87	9
rect	88	8	89	9
rect	89	8	90	9
rect	90	8	91	9
rect	91	8	92	9
rect	92	8	93	9
rect	93	8	94	9
rect	95	8	96	9
rect	96	8	97	9
rect	97	8	98	9
rect	98	8	99	9
rect	99	8	100	9
rect	100	8	101	9
rect	102	8	103	9
rect	103	8	104	9
rect	104	8	105	9
rect	105	8	106	9
rect	106	8	107	9
rect	107	8	108	9
rect	108	8	109	9
rect	109	8	110	9
rect	110	8	111	9
rect	111	8	112	9
rect	112	8	113	9
rect	113	8	114	9
rect	114	8	115	9
rect	115	8	116	9
rect	116	8	117	9
rect	117	8	118	9
rect	118	8	119	9
rect	119	8	120	9
rect	120	8	121	9
rect	121	8	122	9
rect	122	8	123	9
rect	123	8	124	9
rect	124	8	125	9
rect	125	8	126	9
rect	127	8	128	9
rect	128	8	129	9
rect	129	8	130	9
rect	130	8	131	9
rect	131	8	132	9
rect	132	8	133	9
rect	134	8	135	9
rect	135	8	136	9
rect	136	8	137	9
rect	137	8	138	9
rect	138	8	139	9
rect	139	8	140	9
rect	141	8	142	9
rect	142	8	143	9
rect	143	8	144	9
rect	144	8	145	9
rect	145	8	146	9
rect	146	8	147	9
rect	148	8	149	9
rect	149	8	150	9
rect	150	8	151	9
rect	151	8	152	9
rect	152	8	153	9
rect	153	8	154	9
rect	155	8	156	9
rect	156	8	157	9
rect	157	8	158	9
rect	158	8	159	9
rect	159	8	160	9
rect	160	8	161	9
rect	162	8	163	9
rect	163	8	164	9
rect	164	8	165	9
rect	165	8	166	9
rect	166	8	167	9
rect	167	8	168	9
rect	169	8	170	9
rect	170	8	171	9
rect	171	8	172	9
rect	172	8	173	9
rect	173	8	174	9
rect	174	8	175	9
rect	176	8	177	9
rect	177	8	178	9
rect	178	8	179	9
rect	179	8	180	9
rect	180	8	181	9
rect	181	8	182	9
rect	183	8	184	9
rect	184	8	185	9
rect	185	8	186	9
rect	186	8	187	9
rect	187	8	188	9
rect	188	8	189	9
rect	189	8	190	9
rect	190	8	191	9
rect	191	8	192	9
rect	192	8	193	9
rect	193	8	194	9
rect	194	8	195	9
rect	195	8	196	9
rect	196	8	197	9
rect	197	8	198	9
rect	199	8	200	9
rect	200	8	201	9
rect	201	8	202	9
rect	202	8	203	9
rect	203	8	204	9
rect	204	8	205	9
rect	206	8	207	9
rect	207	8	208	9
rect	208	8	209	9
rect	209	8	210	9
rect	210	8	211	9
rect	211	8	212	9
rect	213	8	214	9
rect	214	8	215	9
rect	215	8	216	9
rect	216	8	217	9
rect	217	8	218	9
rect	218	8	219	9
rect	219	8	220	9
rect	220	8	221	9
rect	221	8	222	9
rect	222	8	223	9
rect	223	8	224	9
rect	224	8	225	9
rect	225	8	226	9
rect	226	8	227	9
rect	227	8	228	9
rect	229	8	230	9
rect	230	8	231	9
rect	231	8	232	9
rect	232	8	233	9
rect	233	8	234	9
rect	234	8	235	9
rect	236	8	237	9
rect	237	8	238	9
rect	238	8	239	9
rect	239	8	240	9
rect	240	8	241	9
rect	241	8	242	9
rect	242	8	243	9
rect	243	8	244	9
rect	244	8	245	9
rect	245	8	246	9
rect	246	8	247	9
rect	247	8	248	9
rect	248	8	249	9
rect	249	8	250	9
rect	250	8	251	9
rect	251	8	252	9
rect	252	8	253	9
rect	253	8	254	9
rect	255	8	256	9
rect	256	8	257	9
rect	257	8	258	9
rect	258	8	259	9
rect	259	8	260	9
rect	260	8	261	9
rect	261	8	262	9
rect	262	8	263	9
rect	263	8	264	9
rect	264	8	265	9
rect	265	8	266	9
rect	266	8	267	9
rect	267	8	268	9
rect	268	8	269	9
rect	269	8	270	9
rect	0	9	1	10
rect	1	9	2	10
rect	2	9	3	10
rect	3	9	4	10
rect	4	9	5	10
rect	5	9	6	10
rect	7	9	8	10
rect	8	9	9	10
rect	9	9	10	10
rect	10	9	11	10
rect	11	9	12	10
rect	12	9	13	10
rect	14	9	15	10
rect	15	9	16	10
rect	16	9	17	10
rect	17	9	18	10
rect	18	9	19	10
rect	19	9	20	10
rect	21	9	22	10
rect	22	9	23	10
rect	23	9	24	10
rect	24	9	25	10
rect	25	9	26	10
rect	26	9	27	10
rect	28	9	29	10
rect	29	9	30	10
rect	30	9	31	10
rect	31	9	32	10
rect	32	9	33	10
rect	33	9	34	10
rect	35	9	36	10
rect	36	9	37	10
rect	37	9	38	10
rect	38	9	39	10
rect	39	9	40	10
rect	40	9	41	10
rect	42	9	43	10
rect	43	9	44	10
rect	44	9	45	10
rect	45	9	46	10
rect	46	9	47	10
rect	47	9	48	10
rect	49	9	50	10
rect	50	9	51	10
rect	51	9	52	10
rect	52	9	53	10
rect	53	9	54	10
rect	54	9	55	10
rect	55	9	56	10
rect	56	9	57	10
rect	57	9	58	10
rect	58	9	59	10
rect	59	9	60	10
rect	60	9	61	10
rect	61	9	62	10
rect	62	9	63	10
rect	63	9	64	10
rect	65	9	66	10
rect	66	9	67	10
rect	67	9	68	10
rect	68	9	69	10
rect	69	9	70	10
rect	70	9	71	10
rect	71	9	72	10
rect	72	9	73	10
rect	73	9	74	10
rect	74	9	75	10
rect	75	9	76	10
rect	76	9	77	10
rect	77	9	78	10
rect	78	9	79	10
rect	79	9	80	10
rect	81	9	82	10
rect	82	9	83	10
rect	83	9	84	10
rect	84	9	85	10
rect	85	9	86	10
rect	86	9	87	10
rect	88	9	89	10
rect	89	9	90	10
rect	90	9	91	10
rect	91	9	92	10
rect	92	9	93	10
rect	93	9	94	10
rect	95	9	96	10
rect	96	9	97	10
rect	97	9	98	10
rect	98	9	99	10
rect	99	9	100	10
rect	100	9	101	10
rect	102	9	103	10
rect	103	9	104	10
rect	104	9	105	10
rect	105	9	106	10
rect	106	9	107	10
rect	107	9	108	10
rect	108	9	109	10
rect	109	9	110	10
rect	110	9	111	10
rect	111	9	112	10
rect	112	9	113	10
rect	113	9	114	10
rect	114	9	115	10
rect	115	9	116	10
rect	116	9	117	10
rect	117	9	118	10
rect	118	9	119	10
rect	119	9	120	10
rect	120	9	121	10
rect	121	9	122	10
rect	122	9	123	10
rect	123	9	124	10
rect	124	9	125	10
rect	125	9	126	10
rect	127	9	128	10
rect	128	9	129	10
rect	129	9	130	10
rect	130	9	131	10
rect	131	9	132	10
rect	132	9	133	10
rect	134	9	135	10
rect	135	9	136	10
rect	136	9	137	10
rect	137	9	138	10
rect	138	9	139	10
rect	139	9	140	10
rect	141	9	142	10
rect	142	9	143	10
rect	143	9	144	10
rect	144	9	145	10
rect	145	9	146	10
rect	146	9	147	10
rect	148	9	149	10
rect	149	9	150	10
rect	150	9	151	10
rect	151	9	152	10
rect	152	9	153	10
rect	153	9	154	10
rect	155	9	156	10
rect	156	9	157	10
rect	157	9	158	10
rect	158	9	159	10
rect	159	9	160	10
rect	160	9	161	10
rect	162	9	163	10
rect	163	9	164	10
rect	164	9	165	10
rect	165	9	166	10
rect	166	9	167	10
rect	167	9	168	10
rect	169	9	170	10
rect	170	9	171	10
rect	171	9	172	10
rect	172	9	173	10
rect	173	9	174	10
rect	174	9	175	10
rect	176	9	177	10
rect	177	9	178	10
rect	178	9	179	10
rect	179	9	180	10
rect	180	9	181	10
rect	181	9	182	10
rect	183	9	184	10
rect	184	9	185	10
rect	185	9	186	10
rect	186	9	187	10
rect	187	9	188	10
rect	188	9	189	10
rect	189	9	190	10
rect	190	9	191	10
rect	191	9	192	10
rect	192	9	193	10
rect	193	9	194	10
rect	194	9	195	10
rect	195	9	196	10
rect	196	9	197	10
rect	197	9	198	10
rect	199	9	200	10
rect	200	9	201	10
rect	201	9	202	10
rect	202	9	203	10
rect	203	9	204	10
rect	204	9	205	10
rect	206	9	207	10
rect	207	9	208	10
rect	208	9	209	10
rect	209	9	210	10
rect	210	9	211	10
rect	211	9	212	10
rect	213	9	214	10
rect	214	9	215	10
rect	215	9	216	10
rect	216	9	217	10
rect	217	9	218	10
rect	218	9	219	10
rect	219	9	220	10
rect	220	9	221	10
rect	221	9	222	10
rect	222	9	223	10
rect	223	9	224	10
rect	224	9	225	10
rect	225	9	226	10
rect	226	9	227	10
rect	227	9	228	10
rect	229	9	230	10
rect	230	9	231	10
rect	231	9	232	10
rect	232	9	233	10
rect	233	9	234	10
rect	234	9	235	10
rect	236	9	237	10
rect	237	9	238	10
rect	238	9	239	10
rect	239	9	240	10
rect	240	9	241	10
rect	241	9	242	10
rect	242	9	243	10
rect	243	9	244	10
rect	244	9	245	10
rect	245	9	246	10
rect	246	9	247	10
rect	247	9	248	10
rect	248	9	249	10
rect	249	9	250	10
rect	250	9	251	10
rect	251	9	252	10
rect	252	9	253	10
rect	253	9	254	10
rect	255	9	256	10
rect	256	9	257	10
rect	257	9	258	10
rect	258	9	259	10
rect	259	9	260	10
rect	260	9	261	10
rect	261	9	262	10
rect	262	9	263	10
rect	263	9	264	10
rect	264	9	265	10
rect	265	9	266	10
rect	266	9	267	10
rect	267	9	268	10
rect	268	9	269	10
rect	269	9	270	10
rect	0	10	1	11
rect	1	10	2	11
rect	2	10	3	11
rect	3	10	4	11
rect	4	10	5	11
rect	5	10	6	11
rect	7	10	8	11
rect	8	10	9	11
rect	9	10	10	11
rect	10	10	11	11
rect	11	10	12	11
rect	12	10	13	11
rect	14	10	15	11
rect	15	10	16	11
rect	16	10	17	11
rect	17	10	18	11
rect	18	10	19	11
rect	19	10	20	11
rect	21	10	22	11
rect	22	10	23	11
rect	23	10	24	11
rect	24	10	25	11
rect	25	10	26	11
rect	26	10	27	11
rect	28	10	29	11
rect	29	10	30	11
rect	30	10	31	11
rect	31	10	32	11
rect	32	10	33	11
rect	33	10	34	11
rect	35	10	36	11
rect	36	10	37	11
rect	37	10	38	11
rect	38	10	39	11
rect	39	10	40	11
rect	40	10	41	11
rect	42	10	43	11
rect	43	10	44	11
rect	44	10	45	11
rect	45	10	46	11
rect	46	10	47	11
rect	47	10	48	11
rect	49	10	50	11
rect	50	10	51	11
rect	51	10	52	11
rect	52	10	53	11
rect	53	10	54	11
rect	54	10	55	11
rect	55	10	56	11
rect	56	10	57	11
rect	57	10	58	11
rect	58	10	59	11
rect	59	10	60	11
rect	60	10	61	11
rect	61	10	62	11
rect	62	10	63	11
rect	63	10	64	11
rect	65	10	66	11
rect	66	10	67	11
rect	67	10	68	11
rect	68	10	69	11
rect	69	10	70	11
rect	70	10	71	11
rect	71	10	72	11
rect	72	10	73	11
rect	73	10	74	11
rect	74	10	75	11
rect	75	10	76	11
rect	76	10	77	11
rect	77	10	78	11
rect	78	10	79	11
rect	79	10	80	11
rect	81	10	82	11
rect	82	10	83	11
rect	83	10	84	11
rect	84	10	85	11
rect	85	10	86	11
rect	86	10	87	11
rect	88	10	89	11
rect	89	10	90	11
rect	90	10	91	11
rect	91	10	92	11
rect	92	10	93	11
rect	93	10	94	11
rect	95	10	96	11
rect	96	10	97	11
rect	97	10	98	11
rect	98	10	99	11
rect	99	10	100	11
rect	100	10	101	11
rect	102	10	103	11
rect	103	10	104	11
rect	104	10	105	11
rect	105	10	106	11
rect	106	10	107	11
rect	107	10	108	11
rect	108	10	109	11
rect	109	10	110	11
rect	110	10	111	11
rect	111	10	112	11
rect	112	10	113	11
rect	113	10	114	11
rect	114	10	115	11
rect	115	10	116	11
rect	116	10	117	11
rect	117	10	118	11
rect	118	10	119	11
rect	119	10	120	11
rect	120	10	121	11
rect	121	10	122	11
rect	122	10	123	11
rect	123	10	124	11
rect	124	10	125	11
rect	125	10	126	11
rect	127	10	128	11
rect	128	10	129	11
rect	129	10	130	11
rect	130	10	131	11
rect	131	10	132	11
rect	132	10	133	11
rect	134	10	135	11
rect	135	10	136	11
rect	136	10	137	11
rect	137	10	138	11
rect	138	10	139	11
rect	139	10	140	11
rect	141	10	142	11
rect	142	10	143	11
rect	143	10	144	11
rect	144	10	145	11
rect	145	10	146	11
rect	146	10	147	11
rect	148	10	149	11
rect	149	10	150	11
rect	150	10	151	11
rect	151	10	152	11
rect	152	10	153	11
rect	153	10	154	11
rect	155	10	156	11
rect	156	10	157	11
rect	157	10	158	11
rect	158	10	159	11
rect	159	10	160	11
rect	160	10	161	11
rect	162	10	163	11
rect	163	10	164	11
rect	164	10	165	11
rect	165	10	166	11
rect	166	10	167	11
rect	167	10	168	11
rect	169	10	170	11
rect	170	10	171	11
rect	171	10	172	11
rect	172	10	173	11
rect	173	10	174	11
rect	174	10	175	11
rect	176	10	177	11
rect	177	10	178	11
rect	178	10	179	11
rect	179	10	180	11
rect	180	10	181	11
rect	181	10	182	11
rect	183	10	184	11
rect	184	10	185	11
rect	185	10	186	11
rect	186	10	187	11
rect	187	10	188	11
rect	188	10	189	11
rect	189	10	190	11
rect	190	10	191	11
rect	191	10	192	11
rect	192	10	193	11
rect	193	10	194	11
rect	194	10	195	11
rect	195	10	196	11
rect	196	10	197	11
rect	197	10	198	11
rect	199	10	200	11
rect	200	10	201	11
rect	201	10	202	11
rect	202	10	203	11
rect	203	10	204	11
rect	204	10	205	11
rect	206	10	207	11
rect	207	10	208	11
rect	208	10	209	11
rect	209	10	210	11
rect	210	10	211	11
rect	211	10	212	11
rect	213	10	214	11
rect	214	10	215	11
rect	215	10	216	11
rect	216	10	217	11
rect	217	10	218	11
rect	218	10	219	11
rect	219	10	220	11
rect	220	10	221	11
rect	221	10	222	11
rect	222	10	223	11
rect	223	10	224	11
rect	224	10	225	11
rect	225	10	226	11
rect	226	10	227	11
rect	227	10	228	11
rect	229	10	230	11
rect	230	10	231	11
rect	231	10	232	11
rect	232	10	233	11
rect	233	10	234	11
rect	234	10	235	11
rect	236	10	237	11
rect	237	10	238	11
rect	238	10	239	11
rect	239	10	240	11
rect	240	10	241	11
rect	241	10	242	11
rect	242	10	243	11
rect	243	10	244	11
rect	244	10	245	11
rect	245	10	246	11
rect	246	10	247	11
rect	247	10	248	11
rect	248	10	249	11
rect	249	10	250	11
rect	250	10	251	11
rect	251	10	252	11
rect	252	10	253	11
rect	253	10	254	11
rect	255	10	256	11
rect	256	10	257	11
rect	257	10	258	11
rect	258	10	259	11
rect	259	10	260	11
rect	260	10	261	11
rect	261	10	262	11
rect	262	10	263	11
rect	263	10	264	11
rect	264	10	265	11
rect	265	10	266	11
rect	266	10	267	11
rect	267	10	268	11
rect	268	10	269	11
rect	269	10	270	11
rect	0	11	1	12
rect	1	11	2	12
rect	2	11	3	12
rect	3	11	4	12
rect	4	11	5	12
rect	5	11	6	12
rect	7	11	8	12
rect	8	11	9	12
rect	9	11	10	12
rect	10	11	11	12
rect	11	11	12	12
rect	12	11	13	12
rect	14	11	15	12
rect	15	11	16	12
rect	16	11	17	12
rect	17	11	18	12
rect	18	11	19	12
rect	19	11	20	12
rect	21	11	22	12
rect	22	11	23	12
rect	23	11	24	12
rect	24	11	25	12
rect	25	11	26	12
rect	26	11	27	12
rect	28	11	29	12
rect	29	11	30	12
rect	30	11	31	12
rect	31	11	32	12
rect	32	11	33	12
rect	33	11	34	12
rect	35	11	36	12
rect	36	11	37	12
rect	37	11	38	12
rect	38	11	39	12
rect	39	11	40	12
rect	40	11	41	12
rect	42	11	43	12
rect	43	11	44	12
rect	44	11	45	12
rect	45	11	46	12
rect	46	11	47	12
rect	47	11	48	12
rect	49	11	50	12
rect	50	11	51	12
rect	51	11	52	12
rect	52	11	53	12
rect	53	11	54	12
rect	54	11	55	12
rect	55	11	56	12
rect	56	11	57	12
rect	57	11	58	12
rect	58	11	59	12
rect	59	11	60	12
rect	60	11	61	12
rect	61	11	62	12
rect	62	11	63	12
rect	63	11	64	12
rect	65	11	66	12
rect	66	11	67	12
rect	67	11	68	12
rect	68	11	69	12
rect	69	11	70	12
rect	70	11	71	12
rect	71	11	72	12
rect	72	11	73	12
rect	73	11	74	12
rect	74	11	75	12
rect	75	11	76	12
rect	76	11	77	12
rect	77	11	78	12
rect	78	11	79	12
rect	79	11	80	12
rect	81	11	82	12
rect	82	11	83	12
rect	83	11	84	12
rect	84	11	85	12
rect	85	11	86	12
rect	86	11	87	12
rect	88	11	89	12
rect	89	11	90	12
rect	90	11	91	12
rect	91	11	92	12
rect	92	11	93	12
rect	93	11	94	12
rect	95	11	96	12
rect	96	11	97	12
rect	97	11	98	12
rect	98	11	99	12
rect	99	11	100	12
rect	100	11	101	12
rect	102	11	103	12
rect	103	11	104	12
rect	104	11	105	12
rect	105	11	106	12
rect	106	11	107	12
rect	107	11	108	12
rect	108	11	109	12
rect	109	11	110	12
rect	110	11	111	12
rect	111	11	112	12
rect	112	11	113	12
rect	113	11	114	12
rect	114	11	115	12
rect	115	11	116	12
rect	116	11	117	12
rect	117	11	118	12
rect	118	11	119	12
rect	119	11	120	12
rect	120	11	121	12
rect	121	11	122	12
rect	122	11	123	12
rect	123	11	124	12
rect	124	11	125	12
rect	125	11	126	12
rect	127	11	128	12
rect	128	11	129	12
rect	129	11	130	12
rect	130	11	131	12
rect	131	11	132	12
rect	132	11	133	12
rect	134	11	135	12
rect	135	11	136	12
rect	136	11	137	12
rect	137	11	138	12
rect	138	11	139	12
rect	139	11	140	12
rect	141	11	142	12
rect	142	11	143	12
rect	143	11	144	12
rect	144	11	145	12
rect	145	11	146	12
rect	146	11	147	12
rect	148	11	149	12
rect	149	11	150	12
rect	150	11	151	12
rect	151	11	152	12
rect	152	11	153	12
rect	153	11	154	12
rect	155	11	156	12
rect	156	11	157	12
rect	157	11	158	12
rect	158	11	159	12
rect	159	11	160	12
rect	160	11	161	12
rect	162	11	163	12
rect	163	11	164	12
rect	164	11	165	12
rect	165	11	166	12
rect	166	11	167	12
rect	167	11	168	12
rect	169	11	170	12
rect	170	11	171	12
rect	171	11	172	12
rect	172	11	173	12
rect	173	11	174	12
rect	174	11	175	12
rect	176	11	177	12
rect	177	11	178	12
rect	178	11	179	12
rect	179	11	180	12
rect	180	11	181	12
rect	181	11	182	12
rect	183	11	184	12
rect	184	11	185	12
rect	185	11	186	12
rect	186	11	187	12
rect	187	11	188	12
rect	188	11	189	12
rect	189	11	190	12
rect	190	11	191	12
rect	191	11	192	12
rect	192	11	193	12
rect	193	11	194	12
rect	194	11	195	12
rect	195	11	196	12
rect	196	11	197	12
rect	197	11	198	12
rect	199	11	200	12
rect	200	11	201	12
rect	201	11	202	12
rect	202	11	203	12
rect	203	11	204	12
rect	204	11	205	12
rect	206	11	207	12
rect	207	11	208	12
rect	208	11	209	12
rect	209	11	210	12
rect	210	11	211	12
rect	211	11	212	12
rect	213	11	214	12
rect	214	11	215	12
rect	215	11	216	12
rect	216	11	217	12
rect	217	11	218	12
rect	218	11	219	12
rect	219	11	220	12
rect	220	11	221	12
rect	221	11	222	12
rect	222	11	223	12
rect	223	11	224	12
rect	224	11	225	12
rect	225	11	226	12
rect	226	11	227	12
rect	227	11	228	12
rect	229	11	230	12
rect	230	11	231	12
rect	231	11	232	12
rect	232	11	233	12
rect	233	11	234	12
rect	234	11	235	12
rect	236	11	237	12
rect	237	11	238	12
rect	238	11	239	12
rect	239	11	240	12
rect	240	11	241	12
rect	241	11	242	12
rect	242	11	243	12
rect	243	11	244	12
rect	244	11	245	12
rect	245	11	246	12
rect	246	11	247	12
rect	247	11	248	12
rect	248	11	249	12
rect	249	11	250	12
rect	250	11	251	12
rect	251	11	252	12
rect	252	11	253	12
rect	253	11	254	12
rect	255	11	256	12
rect	256	11	257	12
rect	257	11	258	12
rect	258	11	259	12
rect	259	11	260	12
rect	260	11	261	12
rect	261	11	262	12
rect	262	11	263	12
rect	263	11	264	12
rect	264	11	265	12
rect	265	11	266	12
rect	266	11	267	12
rect	267	11	268	12
rect	268	11	269	12
rect	269	11	270	12
rect	0	27	1	28
rect	1	27	2	28
rect	2	27	3	28
rect	3	27	4	28
rect	4	27	5	28
rect	5	27	6	28
rect	7	27	8	28
rect	8	27	9	28
rect	9	27	10	28
rect	10	27	11	28
rect	11	27	12	28
rect	12	27	13	28
rect	13	27	14	28
rect	14	27	15	28
rect	15	27	16	28
rect	16	27	17	28
rect	17	27	18	28
rect	18	27	19	28
rect	19	27	20	28
rect	20	27	21	28
rect	21	27	22	28
rect	23	27	24	28
rect	24	27	25	28
rect	25	27	26	28
rect	26	27	27	28
rect	27	27	28	28
rect	28	27	29	28
rect	29	27	30	28
rect	30	27	31	28
rect	31	27	32	28
rect	32	27	33	28
rect	33	27	34	28
rect	34	27	35	28
rect	35	27	36	28
rect	36	27	37	28
rect	37	27	38	28
rect	39	27	40	28
rect	40	27	41	28
rect	41	27	42	28
rect	42	27	43	28
rect	43	27	44	28
rect	44	27	45	28
rect	46	27	47	28
rect	47	27	48	28
rect	48	27	49	28
rect	49	27	50	28
rect	50	27	51	28
rect	51	27	52	28
rect	52	27	53	28
rect	53	27	54	28
rect	54	27	55	28
rect	55	27	56	28
rect	56	27	57	28
rect	57	27	58	28
rect	58	27	59	28
rect	59	27	60	28
rect	60	27	61	28
rect	61	27	62	28
rect	62	27	63	28
rect	63	27	64	28
rect	64	27	65	28
rect	65	27	66	28
rect	66	27	67	28
rect	67	27	68	28
rect	68	27	69	28
rect	69	27	70	28
rect	70	27	71	28
rect	71	27	72	28
rect	72	27	73	28
rect	73	27	74	28
rect	74	27	75	28
rect	75	27	76	28
rect	76	27	77	28
rect	77	27	78	28
rect	78	27	79	28
rect	80	27	81	28
rect	81	27	82	28
rect	82	27	83	28
rect	83	27	84	28
rect	84	27	85	28
rect	85	27	86	28
rect	87	27	88	28
rect	88	27	89	28
rect	89	27	90	28
rect	90	27	91	28
rect	91	27	92	28
rect	92	27	93	28
rect	94	27	95	28
rect	95	27	96	28
rect	96	27	97	28
rect	97	27	98	28
rect	98	27	99	28
rect	99	27	100	28
rect	101	27	102	28
rect	102	27	103	28
rect	103	27	104	28
rect	104	27	105	28
rect	105	27	106	28
rect	106	27	107	28
rect	107	27	108	28
rect	108	27	109	28
rect	109	27	110	28
rect	110	27	111	28
rect	111	27	112	28
rect	112	27	113	28
rect	113	27	114	28
rect	114	27	115	28
rect	115	27	116	28
rect	117	27	118	28
rect	118	27	119	28
rect	119	27	120	28
rect	120	27	121	28
rect	121	27	122	28
rect	122	27	123	28
rect	124	27	125	28
rect	125	27	126	28
rect	126	27	127	28
rect	127	27	128	28
rect	128	27	129	28
rect	129	27	130	28
rect	131	27	132	28
rect	132	27	133	28
rect	133	27	134	28
rect	134	27	135	28
rect	135	27	136	28
rect	136	27	137	28
rect	138	27	139	28
rect	139	27	140	28
rect	140	27	141	28
rect	141	27	142	28
rect	142	27	143	28
rect	143	27	144	28
rect	145	27	146	28
rect	146	27	147	28
rect	147	27	148	28
rect	148	27	149	28
rect	149	27	150	28
rect	150	27	151	28
rect	151	27	152	28
rect	152	27	153	28
rect	153	27	154	28
rect	154	27	155	28
rect	155	27	156	28
rect	156	27	157	28
rect	157	27	158	28
rect	158	27	159	28
rect	159	27	160	28
rect	160	27	161	28
rect	161	27	162	28
rect	162	27	163	28
rect	163	27	164	28
rect	164	27	165	28
rect	165	27	166	28
rect	166	27	167	28
rect	167	27	168	28
rect	168	27	169	28
rect	169	27	170	28
rect	170	27	171	28
rect	171	27	172	28
rect	172	27	173	28
rect	173	27	174	28
rect	174	27	175	28
rect	175	27	176	28
rect	176	27	177	28
rect	177	27	178	28
rect	178	27	179	28
rect	179	27	180	28
rect	180	27	181	28
rect	181	27	182	28
rect	182	27	183	28
rect	183	27	184	28
rect	184	27	185	28
rect	185	27	186	28
rect	186	27	187	28
rect	187	27	188	28
rect	188	27	189	28
rect	189	27	190	28
rect	190	27	191	28
rect	191	27	192	28
rect	192	27	193	28
rect	193	27	194	28
rect	194	27	195	28
rect	195	27	196	28
rect	196	27	197	28
rect	197	27	198	28
rect	198	27	199	28
rect	199	27	200	28
rect	200	27	201	28
rect	201	27	202	28
rect	202	27	203	28
rect	203	27	204	28
rect	204	27	205	28
rect	205	27	206	28
rect	206	27	207	28
rect	207	27	208	28
rect	208	27	209	28
rect	209	27	210	28
rect	210	27	211	28
rect	211	27	212	28
rect	212	27	213	28
rect	213	27	214	28
rect	214	27	215	28
rect	215	27	216	28
rect	216	27	217	28
rect	217	27	218	28
rect	218	27	219	28
rect	219	27	220	28
rect	220	27	221	28
rect	221	27	222	28
rect	222	27	223	28
rect	223	27	224	28
rect	224	27	225	28
rect	225	27	226	28
rect	226	27	227	28
rect	227	27	228	28
rect	228	27	229	28
rect	230	27	231	28
rect	231	27	232	28
rect	232	27	233	28
rect	233	27	234	28
rect	234	27	235	28
rect	235	27	236	28
rect	237	27	238	28
rect	238	27	239	28
rect	239	27	240	28
rect	240	27	241	28
rect	241	27	242	28
rect	242	27	243	28
rect	243	27	244	28
rect	244	27	245	28
rect	245	27	246	28
rect	246	27	247	28
rect	247	27	248	28
rect	248	27	249	28
rect	249	27	250	28
rect	250	27	251	28
rect	251	27	252	28
rect	252	27	253	28
rect	253	27	254	28
rect	254	27	255	28
rect	255	27	256	28
rect	256	27	257	28
rect	257	27	258	28
rect	258	27	259	28
rect	259	27	260	28
rect	260	27	261	28
rect	261	27	262	28
rect	262	27	263	28
rect	263	27	264	28
rect	264	27	265	28
rect	265	27	266	28
rect	266	27	267	28
rect	267	27	268	28
rect	268	27	269	28
rect	269	27	270	28
rect	270	27	271	28
rect	271	27	272	28
rect	272	27	273	28
rect	274	27	275	28
rect	275	27	276	28
rect	276	27	277	28
rect	277	27	278	28
rect	278	27	279	28
rect	279	27	280	28
rect	281	27	282	28
rect	282	27	283	28
rect	283	27	284	28
rect	284	27	285	28
rect	285	27	286	28
rect	286	27	287	28
rect	288	27	289	28
rect	289	27	290	28
rect	290	27	291	28
rect	291	27	292	28
rect	292	27	293	28
rect	293	27	294	28
rect	295	27	296	28
rect	296	27	297	28
rect	297	27	298	28
rect	298	27	299	28
rect	299	27	300	28
rect	300	27	301	28
rect	301	27	302	28
rect	302	27	303	28
rect	303	27	304	28
rect	304	27	305	28
rect	305	27	306	28
rect	306	27	307	28
rect	0	28	1	29
rect	1	28	2	29
rect	2	28	3	29
rect	3	28	4	29
rect	4	28	5	29
rect	5	28	6	29
rect	7	28	8	29
rect	8	28	9	29
rect	9	28	10	29
rect	10	28	11	29
rect	11	28	12	29
rect	12	28	13	29
rect	13	28	14	29
rect	14	28	15	29
rect	15	28	16	29
rect	16	28	17	29
rect	17	28	18	29
rect	18	28	19	29
rect	19	28	20	29
rect	20	28	21	29
rect	21	28	22	29
rect	23	28	24	29
rect	24	28	25	29
rect	25	28	26	29
rect	26	28	27	29
rect	27	28	28	29
rect	28	28	29	29
rect	29	28	30	29
rect	30	28	31	29
rect	31	28	32	29
rect	32	28	33	29
rect	33	28	34	29
rect	34	28	35	29
rect	35	28	36	29
rect	36	28	37	29
rect	37	28	38	29
rect	39	28	40	29
rect	40	28	41	29
rect	41	28	42	29
rect	42	28	43	29
rect	43	28	44	29
rect	44	28	45	29
rect	46	28	47	29
rect	47	28	48	29
rect	48	28	49	29
rect	49	28	50	29
rect	50	28	51	29
rect	51	28	52	29
rect	52	28	53	29
rect	53	28	54	29
rect	54	28	55	29
rect	55	28	56	29
rect	56	28	57	29
rect	57	28	58	29
rect	58	28	59	29
rect	59	28	60	29
rect	60	28	61	29
rect	61	28	62	29
rect	62	28	63	29
rect	63	28	64	29
rect	64	28	65	29
rect	65	28	66	29
rect	66	28	67	29
rect	67	28	68	29
rect	68	28	69	29
rect	69	28	70	29
rect	70	28	71	29
rect	71	28	72	29
rect	72	28	73	29
rect	73	28	74	29
rect	74	28	75	29
rect	75	28	76	29
rect	76	28	77	29
rect	77	28	78	29
rect	78	28	79	29
rect	80	28	81	29
rect	81	28	82	29
rect	82	28	83	29
rect	83	28	84	29
rect	84	28	85	29
rect	85	28	86	29
rect	87	28	88	29
rect	88	28	89	29
rect	89	28	90	29
rect	90	28	91	29
rect	91	28	92	29
rect	92	28	93	29
rect	94	28	95	29
rect	95	28	96	29
rect	96	28	97	29
rect	97	28	98	29
rect	98	28	99	29
rect	99	28	100	29
rect	101	28	102	29
rect	102	28	103	29
rect	103	28	104	29
rect	104	28	105	29
rect	105	28	106	29
rect	106	28	107	29
rect	107	28	108	29
rect	108	28	109	29
rect	109	28	110	29
rect	110	28	111	29
rect	111	28	112	29
rect	112	28	113	29
rect	113	28	114	29
rect	114	28	115	29
rect	115	28	116	29
rect	117	28	118	29
rect	118	28	119	29
rect	119	28	120	29
rect	120	28	121	29
rect	121	28	122	29
rect	122	28	123	29
rect	124	28	125	29
rect	125	28	126	29
rect	126	28	127	29
rect	127	28	128	29
rect	128	28	129	29
rect	129	28	130	29
rect	131	28	132	29
rect	132	28	133	29
rect	133	28	134	29
rect	134	28	135	29
rect	135	28	136	29
rect	136	28	137	29
rect	138	28	139	29
rect	139	28	140	29
rect	140	28	141	29
rect	141	28	142	29
rect	142	28	143	29
rect	143	28	144	29
rect	145	28	146	29
rect	146	28	147	29
rect	147	28	148	29
rect	148	28	149	29
rect	149	28	150	29
rect	150	28	151	29
rect	151	28	152	29
rect	152	28	153	29
rect	153	28	154	29
rect	154	28	155	29
rect	155	28	156	29
rect	156	28	157	29
rect	157	28	158	29
rect	158	28	159	29
rect	159	28	160	29
rect	160	28	161	29
rect	161	28	162	29
rect	162	28	163	29
rect	163	28	164	29
rect	164	28	165	29
rect	165	28	166	29
rect	166	28	167	29
rect	167	28	168	29
rect	168	28	169	29
rect	169	28	170	29
rect	170	28	171	29
rect	171	28	172	29
rect	172	28	173	29
rect	173	28	174	29
rect	174	28	175	29
rect	175	28	176	29
rect	176	28	177	29
rect	177	28	178	29
rect	178	28	179	29
rect	179	28	180	29
rect	180	28	181	29
rect	181	28	182	29
rect	182	28	183	29
rect	183	28	184	29
rect	184	28	185	29
rect	185	28	186	29
rect	186	28	187	29
rect	187	28	188	29
rect	188	28	189	29
rect	189	28	190	29
rect	190	28	191	29
rect	191	28	192	29
rect	192	28	193	29
rect	193	28	194	29
rect	194	28	195	29
rect	195	28	196	29
rect	196	28	197	29
rect	197	28	198	29
rect	198	28	199	29
rect	199	28	200	29
rect	200	28	201	29
rect	201	28	202	29
rect	202	28	203	29
rect	203	28	204	29
rect	204	28	205	29
rect	205	28	206	29
rect	206	28	207	29
rect	207	28	208	29
rect	208	28	209	29
rect	209	28	210	29
rect	210	28	211	29
rect	211	28	212	29
rect	212	28	213	29
rect	213	28	214	29
rect	214	28	215	29
rect	215	28	216	29
rect	216	28	217	29
rect	217	28	218	29
rect	218	28	219	29
rect	219	28	220	29
rect	220	28	221	29
rect	221	28	222	29
rect	222	28	223	29
rect	223	28	224	29
rect	224	28	225	29
rect	225	28	226	29
rect	226	28	227	29
rect	227	28	228	29
rect	228	28	229	29
rect	230	28	231	29
rect	231	28	232	29
rect	232	28	233	29
rect	233	28	234	29
rect	234	28	235	29
rect	235	28	236	29
rect	237	28	238	29
rect	238	28	239	29
rect	239	28	240	29
rect	240	28	241	29
rect	241	28	242	29
rect	242	28	243	29
rect	243	28	244	29
rect	244	28	245	29
rect	245	28	246	29
rect	246	28	247	29
rect	247	28	248	29
rect	248	28	249	29
rect	249	28	250	29
rect	250	28	251	29
rect	251	28	252	29
rect	252	28	253	29
rect	253	28	254	29
rect	254	28	255	29
rect	255	28	256	29
rect	256	28	257	29
rect	257	28	258	29
rect	258	28	259	29
rect	259	28	260	29
rect	260	28	261	29
rect	261	28	262	29
rect	262	28	263	29
rect	263	28	264	29
rect	264	28	265	29
rect	265	28	266	29
rect	266	28	267	29
rect	267	28	268	29
rect	268	28	269	29
rect	269	28	270	29
rect	270	28	271	29
rect	271	28	272	29
rect	272	28	273	29
rect	274	28	275	29
rect	275	28	276	29
rect	276	28	277	29
rect	277	28	278	29
rect	278	28	279	29
rect	279	28	280	29
rect	281	28	282	29
rect	282	28	283	29
rect	283	28	284	29
rect	284	28	285	29
rect	285	28	286	29
rect	286	28	287	29
rect	288	28	289	29
rect	289	28	290	29
rect	290	28	291	29
rect	291	28	292	29
rect	292	28	293	29
rect	293	28	294	29
rect	295	28	296	29
rect	296	28	297	29
rect	297	28	298	29
rect	298	28	299	29
rect	299	28	300	29
rect	300	28	301	29
rect	301	28	302	29
rect	302	28	303	29
rect	303	28	304	29
rect	304	28	305	29
rect	305	28	306	29
rect	306	28	307	29
rect	0	29	1	30
rect	1	29	2	30
rect	2	29	3	30
rect	3	29	4	30
rect	4	29	5	30
rect	5	29	6	30
rect	7	29	8	30
rect	8	29	9	30
rect	9	29	10	30
rect	10	29	11	30
rect	11	29	12	30
rect	12	29	13	30
rect	13	29	14	30
rect	14	29	15	30
rect	15	29	16	30
rect	16	29	17	30
rect	17	29	18	30
rect	18	29	19	30
rect	19	29	20	30
rect	20	29	21	30
rect	21	29	22	30
rect	23	29	24	30
rect	24	29	25	30
rect	25	29	26	30
rect	26	29	27	30
rect	27	29	28	30
rect	28	29	29	30
rect	29	29	30	30
rect	30	29	31	30
rect	31	29	32	30
rect	32	29	33	30
rect	33	29	34	30
rect	34	29	35	30
rect	35	29	36	30
rect	36	29	37	30
rect	37	29	38	30
rect	39	29	40	30
rect	40	29	41	30
rect	41	29	42	30
rect	42	29	43	30
rect	43	29	44	30
rect	44	29	45	30
rect	46	29	47	30
rect	47	29	48	30
rect	48	29	49	30
rect	49	29	50	30
rect	50	29	51	30
rect	51	29	52	30
rect	52	29	53	30
rect	53	29	54	30
rect	54	29	55	30
rect	55	29	56	30
rect	56	29	57	30
rect	57	29	58	30
rect	58	29	59	30
rect	59	29	60	30
rect	60	29	61	30
rect	61	29	62	30
rect	62	29	63	30
rect	63	29	64	30
rect	64	29	65	30
rect	65	29	66	30
rect	66	29	67	30
rect	67	29	68	30
rect	68	29	69	30
rect	69	29	70	30
rect	70	29	71	30
rect	71	29	72	30
rect	72	29	73	30
rect	73	29	74	30
rect	74	29	75	30
rect	75	29	76	30
rect	76	29	77	30
rect	77	29	78	30
rect	78	29	79	30
rect	80	29	81	30
rect	81	29	82	30
rect	82	29	83	30
rect	83	29	84	30
rect	84	29	85	30
rect	85	29	86	30
rect	87	29	88	30
rect	88	29	89	30
rect	89	29	90	30
rect	90	29	91	30
rect	91	29	92	30
rect	92	29	93	30
rect	94	29	95	30
rect	95	29	96	30
rect	96	29	97	30
rect	97	29	98	30
rect	98	29	99	30
rect	99	29	100	30
rect	101	29	102	30
rect	102	29	103	30
rect	103	29	104	30
rect	104	29	105	30
rect	105	29	106	30
rect	106	29	107	30
rect	107	29	108	30
rect	108	29	109	30
rect	109	29	110	30
rect	110	29	111	30
rect	111	29	112	30
rect	112	29	113	30
rect	113	29	114	30
rect	114	29	115	30
rect	115	29	116	30
rect	117	29	118	30
rect	118	29	119	30
rect	119	29	120	30
rect	120	29	121	30
rect	121	29	122	30
rect	122	29	123	30
rect	124	29	125	30
rect	125	29	126	30
rect	126	29	127	30
rect	127	29	128	30
rect	128	29	129	30
rect	129	29	130	30
rect	131	29	132	30
rect	132	29	133	30
rect	133	29	134	30
rect	134	29	135	30
rect	135	29	136	30
rect	136	29	137	30
rect	138	29	139	30
rect	139	29	140	30
rect	140	29	141	30
rect	141	29	142	30
rect	142	29	143	30
rect	143	29	144	30
rect	145	29	146	30
rect	146	29	147	30
rect	147	29	148	30
rect	148	29	149	30
rect	149	29	150	30
rect	150	29	151	30
rect	151	29	152	30
rect	152	29	153	30
rect	153	29	154	30
rect	154	29	155	30
rect	155	29	156	30
rect	156	29	157	30
rect	157	29	158	30
rect	158	29	159	30
rect	159	29	160	30
rect	160	29	161	30
rect	161	29	162	30
rect	162	29	163	30
rect	163	29	164	30
rect	164	29	165	30
rect	165	29	166	30
rect	166	29	167	30
rect	167	29	168	30
rect	168	29	169	30
rect	169	29	170	30
rect	170	29	171	30
rect	171	29	172	30
rect	172	29	173	30
rect	173	29	174	30
rect	174	29	175	30
rect	175	29	176	30
rect	176	29	177	30
rect	177	29	178	30
rect	178	29	179	30
rect	179	29	180	30
rect	180	29	181	30
rect	181	29	182	30
rect	182	29	183	30
rect	183	29	184	30
rect	184	29	185	30
rect	185	29	186	30
rect	186	29	187	30
rect	187	29	188	30
rect	188	29	189	30
rect	189	29	190	30
rect	190	29	191	30
rect	191	29	192	30
rect	192	29	193	30
rect	193	29	194	30
rect	194	29	195	30
rect	195	29	196	30
rect	196	29	197	30
rect	197	29	198	30
rect	198	29	199	30
rect	199	29	200	30
rect	200	29	201	30
rect	201	29	202	30
rect	202	29	203	30
rect	203	29	204	30
rect	204	29	205	30
rect	205	29	206	30
rect	206	29	207	30
rect	207	29	208	30
rect	208	29	209	30
rect	209	29	210	30
rect	210	29	211	30
rect	211	29	212	30
rect	212	29	213	30
rect	213	29	214	30
rect	214	29	215	30
rect	215	29	216	30
rect	216	29	217	30
rect	217	29	218	30
rect	218	29	219	30
rect	219	29	220	30
rect	220	29	221	30
rect	221	29	222	30
rect	222	29	223	30
rect	223	29	224	30
rect	224	29	225	30
rect	225	29	226	30
rect	226	29	227	30
rect	227	29	228	30
rect	228	29	229	30
rect	230	29	231	30
rect	231	29	232	30
rect	232	29	233	30
rect	233	29	234	30
rect	234	29	235	30
rect	235	29	236	30
rect	237	29	238	30
rect	238	29	239	30
rect	239	29	240	30
rect	240	29	241	30
rect	241	29	242	30
rect	242	29	243	30
rect	243	29	244	30
rect	244	29	245	30
rect	245	29	246	30
rect	246	29	247	30
rect	247	29	248	30
rect	248	29	249	30
rect	249	29	250	30
rect	250	29	251	30
rect	251	29	252	30
rect	252	29	253	30
rect	253	29	254	30
rect	254	29	255	30
rect	255	29	256	30
rect	256	29	257	30
rect	257	29	258	30
rect	258	29	259	30
rect	259	29	260	30
rect	260	29	261	30
rect	261	29	262	30
rect	262	29	263	30
rect	263	29	264	30
rect	264	29	265	30
rect	265	29	266	30
rect	266	29	267	30
rect	267	29	268	30
rect	268	29	269	30
rect	269	29	270	30
rect	270	29	271	30
rect	271	29	272	30
rect	272	29	273	30
rect	274	29	275	30
rect	275	29	276	30
rect	276	29	277	30
rect	277	29	278	30
rect	278	29	279	30
rect	279	29	280	30
rect	281	29	282	30
rect	282	29	283	30
rect	283	29	284	30
rect	284	29	285	30
rect	285	29	286	30
rect	286	29	287	30
rect	288	29	289	30
rect	289	29	290	30
rect	290	29	291	30
rect	291	29	292	30
rect	292	29	293	30
rect	293	29	294	30
rect	295	29	296	30
rect	296	29	297	30
rect	297	29	298	30
rect	298	29	299	30
rect	299	29	300	30
rect	300	29	301	30
rect	301	29	302	30
rect	302	29	303	30
rect	303	29	304	30
rect	304	29	305	30
rect	305	29	306	30
rect	306	29	307	30
rect	0	30	1	31
rect	1	30	2	31
rect	2	30	3	31
rect	3	30	4	31
rect	4	30	5	31
rect	5	30	6	31
rect	7	30	8	31
rect	8	30	9	31
rect	9	30	10	31
rect	10	30	11	31
rect	11	30	12	31
rect	12	30	13	31
rect	13	30	14	31
rect	14	30	15	31
rect	15	30	16	31
rect	16	30	17	31
rect	17	30	18	31
rect	18	30	19	31
rect	19	30	20	31
rect	20	30	21	31
rect	21	30	22	31
rect	23	30	24	31
rect	24	30	25	31
rect	25	30	26	31
rect	26	30	27	31
rect	27	30	28	31
rect	28	30	29	31
rect	29	30	30	31
rect	30	30	31	31
rect	31	30	32	31
rect	32	30	33	31
rect	33	30	34	31
rect	34	30	35	31
rect	35	30	36	31
rect	36	30	37	31
rect	37	30	38	31
rect	39	30	40	31
rect	40	30	41	31
rect	41	30	42	31
rect	42	30	43	31
rect	43	30	44	31
rect	44	30	45	31
rect	46	30	47	31
rect	47	30	48	31
rect	48	30	49	31
rect	49	30	50	31
rect	50	30	51	31
rect	51	30	52	31
rect	52	30	53	31
rect	53	30	54	31
rect	54	30	55	31
rect	55	30	56	31
rect	56	30	57	31
rect	57	30	58	31
rect	58	30	59	31
rect	59	30	60	31
rect	60	30	61	31
rect	61	30	62	31
rect	62	30	63	31
rect	63	30	64	31
rect	64	30	65	31
rect	65	30	66	31
rect	66	30	67	31
rect	67	30	68	31
rect	68	30	69	31
rect	69	30	70	31
rect	70	30	71	31
rect	71	30	72	31
rect	72	30	73	31
rect	73	30	74	31
rect	74	30	75	31
rect	75	30	76	31
rect	76	30	77	31
rect	77	30	78	31
rect	78	30	79	31
rect	80	30	81	31
rect	81	30	82	31
rect	82	30	83	31
rect	83	30	84	31
rect	84	30	85	31
rect	85	30	86	31
rect	87	30	88	31
rect	88	30	89	31
rect	89	30	90	31
rect	90	30	91	31
rect	91	30	92	31
rect	92	30	93	31
rect	94	30	95	31
rect	95	30	96	31
rect	96	30	97	31
rect	97	30	98	31
rect	98	30	99	31
rect	99	30	100	31
rect	101	30	102	31
rect	102	30	103	31
rect	103	30	104	31
rect	104	30	105	31
rect	105	30	106	31
rect	106	30	107	31
rect	107	30	108	31
rect	108	30	109	31
rect	109	30	110	31
rect	110	30	111	31
rect	111	30	112	31
rect	112	30	113	31
rect	113	30	114	31
rect	114	30	115	31
rect	115	30	116	31
rect	117	30	118	31
rect	118	30	119	31
rect	119	30	120	31
rect	120	30	121	31
rect	121	30	122	31
rect	122	30	123	31
rect	124	30	125	31
rect	125	30	126	31
rect	126	30	127	31
rect	127	30	128	31
rect	128	30	129	31
rect	129	30	130	31
rect	131	30	132	31
rect	132	30	133	31
rect	133	30	134	31
rect	134	30	135	31
rect	135	30	136	31
rect	136	30	137	31
rect	138	30	139	31
rect	139	30	140	31
rect	140	30	141	31
rect	141	30	142	31
rect	142	30	143	31
rect	143	30	144	31
rect	145	30	146	31
rect	146	30	147	31
rect	147	30	148	31
rect	148	30	149	31
rect	149	30	150	31
rect	150	30	151	31
rect	151	30	152	31
rect	152	30	153	31
rect	153	30	154	31
rect	154	30	155	31
rect	155	30	156	31
rect	156	30	157	31
rect	157	30	158	31
rect	158	30	159	31
rect	159	30	160	31
rect	160	30	161	31
rect	161	30	162	31
rect	162	30	163	31
rect	163	30	164	31
rect	164	30	165	31
rect	165	30	166	31
rect	166	30	167	31
rect	167	30	168	31
rect	168	30	169	31
rect	169	30	170	31
rect	170	30	171	31
rect	171	30	172	31
rect	172	30	173	31
rect	173	30	174	31
rect	174	30	175	31
rect	175	30	176	31
rect	176	30	177	31
rect	177	30	178	31
rect	178	30	179	31
rect	179	30	180	31
rect	180	30	181	31
rect	181	30	182	31
rect	182	30	183	31
rect	183	30	184	31
rect	184	30	185	31
rect	185	30	186	31
rect	186	30	187	31
rect	187	30	188	31
rect	188	30	189	31
rect	189	30	190	31
rect	190	30	191	31
rect	191	30	192	31
rect	192	30	193	31
rect	193	30	194	31
rect	194	30	195	31
rect	195	30	196	31
rect	196	30	197	31
rect	197	30	198	31
rect	198	30	199	31
rect	199	30	200	31
rect	200	30	201	31
rect	201	30	202	31
rect	202	30	203	31
rect	203	30	204	31
rect	204	30	205	31
rect	205	30	206	31
rect	206	30	207	31
rect	207	30	208	31
rect	208	30	209	31
rect	209	30	210	31
rect	210	30	211	31
rect	211	30	212	31
rect	212	30	213	31
rect	213	30	214	31
rect	214	30	215	31
rect	215	30	216	31
rect	216	30	217	31
rect	217	30	218	31
rect	218	30	219	31
rect	219	30	220	31
rect	220	30	221	31
rect	221	30	222	31
rect	222	30	223	31
rect	223	30	224	31
rect	224	30	225	31
rect	225	30	226	31
rect	226	30	227	31
rect	227	30	228	31
rect	228	30	229	31
rect	230	30	231	31
rect	231	30	232	31
rect	232	30	233	31
rect	233	30	234	31
rect	234	30	235	31
rect	235	30	236	31
rect	237	30	238	31
rect	238	30	239	31
rect	239	30	240	31
rect	240	30	241	31
rect	241	30	242	31
rect	242	30	243	31
rect	243	30	244	31
rect	244	30	245	31
rect	245	30	246	31
rect	246	30	247	31
rect	247	30	248	31
rect	248	30	249	31
rect	249	30	250	31
rect	250	30	251	31
rect	251	30	252	31
rect	252	30	253	31
rect	253	30	254	31
rect	254	30	255	31
rect	255	30	256	31
rect	256	30	257	31
rect	257	30	258	31
rect	258	30	259	31
rect	259	30	260	31
rect	260	30	261	31
rect	261	30	262	31
rect	262	30	263	31
rect	263	30	264	31
rect	264	30	265	31
rect	265	30	266	31
rect	266	30	267	31
rect	267	30	268	31
rect	268	30	269	31
rect	269	30	270	31
rect	270	30	271	31
rect	271	30	272	31
rect	272	30	273	31
rect	274	30	275	31
rect	275	30	276	31
rect	276	30	277	31
rect	277	30	278	31
rect	278	30	279	31
rect	279	30	280	31
rect	281	30	282	31
rect	282	30	283	31
rect	283	30	284	31
rect	284	30	285	31
rect	285	30	286	31
rect	286	30	287	31
rect	288	30	289	31
rect	289	30	290	31
rect	290	30	291	31
rect	291	30	292	31
rect	292	30	293	31
rect	293	30	294	31
rect	295	30	296	31
rect	296	30	297	31
rect	297	30	298	31
rect	298	30	299	31
rect	299	30	300	31
rect	300	30	301	31
rect	301	30	302	31
rect	302	30	303	31
rect	303	30	304	31
rect	304	30	305	31
rect	305	30	306	31
rect	306	30	307	31
rect	0	31	1	32
rect	1	31	2	32
rect	2	31	3	32
rect	3	31	4	32
rect	4	31	5	32
rect	5	31	6	32
rect	7	31	8	32
rect	8	31	9	32
rect	9	31	10	32
rect	10	31	11	32
rect	11	31	12	32
rect	12	31	13	32
rect	13	31	14	32
rect	14	31	15	32
rect	15	31	16	32
rect	16	31	17	32
rect	17	31	18	32
rect	18	31	19	32
rect	19	31	20	32
rect	20	31	21	32
rect	21	31	22	32
rect	23	31	24	32
rect	24	31	25	32
rect	25	31	26	32
rect	26	31	27	32
rect	27	31	28	32
rect	28	31	29	32
rect	29	31	30	32
rect	30	31	31	32
rect	31	31	32	32
rect	32	31	33	32
rect	33	31	34	32
rect	34	31	35	32
rect	35	31	36	32
rect	36	31	37	32
rect	37	31	38	32
rect	39	31	40	32
rect	40	31	41	32
rect	41	31	42	32
rect	42	31	43	32
rect	43	31	44	32
rect	44	31	45	32
rect	46	31	47	32
rect	47	31	48	32
rect	48	31	49	32
rect	49	31	50	32
rect	50	31	51	32
rect	51	31	52	32
rect	52	31	53	32
rect	53	31	54	32
rect	54	31	55	32
rect	55	31	56	32
rect	56	31	57	32
rect	57	31	58	32
rect	58	31	59	32
rect	59	31	60	32
rect	60	31	61	32
rect	61	31	62	32
rect	62	31	63	32
rect	63	31	64	32
rect	64	31	65	32
rect	65	31	66	32
rect	66	31	67	32
rect	67	31	68	32
rect	68	31	69	32
rect	69	31	70	32
rect	70	31	71	32
rect	71	31	72	32
rect	72	31	73	32
rect	73	31	74	32
rect	74	31	75	32
rect	75	31	76	32
rect	76	31	77	32
rect	77	31	78	32
rect	78	31	79	32
rect	80	31	81	32
rect	81	31	82	32
rect	82	31	83	32
rect	83	31	84	32
rect	84	31	85	32
rect	85	31	86	32
rect	87	31	88	32
rect	88	31	89	32
rect	89	31	90	32
rect	90	31	91	32
rect	91	31	92	32
rect	92	31	93	32
rect	94	31	95	32
rect	95	31	96	32
rect	96	31	97	32
rect	97	31	98	32
rect	98	31	99	32
rect	99	31	100	32
rect	101	31	102	32
rect	102	31	103	32
rect	103	31	104	32
rect	104	31	105	32
rect	105	31	106	32
rect	106	31	107	32
rect	107	31	108	32
rect	108	31	109	32
rect	109	31	110	32
rect	110	31	111	32
rect	111	31	112	32
rect	112	31	113	32
rect	113	31	114	32
rect	114	31	115	32
rect	115	31	116	32
rect	117	31	118	32
rect	118	31	119	32
rect	119	31	120	32
rect	120	31	121	32
rect	121	31	122	32
rect	122	31	123	32
rect	124	31	125	32
rect	125	31	126	32
rect	126	31	127	32
rect	127	31	128	32
rect	128	31	129	32
rect	129	31	130	32
rect	131	31	132	32
rect	132	31	133	32
rect	133	31	134	32
rect	134	31	135	32
rect	135	31	136	32
rect	136	31	137	32
rect	138	31	139	32
rect	139	31	140	32
rect	140	31	141	32
rect	141	31	142	32
rect	142	31	143	32
rect	143	31	144	32
rect	145	31	146	32
rect	146	31	147	32
rect	147	31	148	32
rect	148	31	149	32
rect	149	31	150	32
rect	150	31	151	32
rect	151	31	152	32
rect	152	31	153	32
rect	153	31	154	32
rect	154	31	155	32
rect	155	31	156	32
rect	156	31	157	32
rect	157	31	158	32
rect	158	31	159	32
rect	159	31	160	32
rect	160	31	161	32
rect	161	31	162	32
rect	162	31	163	32
rect	163	31	164	32
rect	164	31	165	32
rect	165	31	166	32
rect	166	31	167	32
rect	167	31	168	32
rect	168	31	169	32
rect	169	31	170	32
rect	170	31	171	32
rect	171	31	172	32
rect	172	31	173	32
rect	173	31	174	32
rect	174	31	175	32
rect	175	31	176	32
rect	176	31	177	32
rect	177	31	178	32
rect	178	31	179	32
rect	179	31	180	32
rect	180	31	181	32
rect	181	31	182	32
rect	182	31	183	32
rect	183	31	184	32
rect	184	31	185	32
rect	185	31	186	32
rect	186	31	187	32
rect	187	31	188	32
rect	188	31	189	32
rect	189	31	190	32
rect	190	31	191	32
rect	191	31	192	32
rect	192	31	193	32
rect	193	31	194	32
rect	194	31	195	32
rect	195	31	196	32
rect	196	31	197	32
rect	197	31	198	32
rect	198	31	199	32
rect	199	31	200	32
rect	200	31	201	32
rect	201	31	202	32
rect	202	31	203	32
rect	203	31	204	32
rect	204	31	205	32
rect	205	31	206	32
rect	206	31	207	32
rect	207	31	208	32
rect	208	31	209	32
rect	209	31	210	32
rect	210	31	211	32
rect	211	31	212	32
rect	212	31	213	32
rect	213	31	214	32
rect	214	31	215	32
rect	215	31	216	32
rect	216	31	217	32
rect	217	31	218	32
rect	218	31	219	32
rect	219	31	220	32
rect	220	31	221	32
rect	221	31	222	32
rect	222	31	223	32
rect	223	31	224	32
rect	224	31	225	32
rect	225	31	226	32
rect	226	31	227	32
rect	227	31	228	32
rect	228	31	229	32
rect	230	31	231	32
rect	231	31	232	32
rect	232	31	233	32
rect	233	31	234	32
rect	234	31	235	32
rect	235	31	236	32
rect	237	31	238	32
rect	238	31	239	32
rect	239	31	240	32
rect	240	31	241	32
rect	241	31	242	32
rect	242	31	243	32
rect	243	31	244	32
rect	244	31	245	32
rect	245	31	246	32
rect	246	31	247	32
rect	247	31	248	32
rect	248	31	249	32
rect	249	31	250	32
rect	250	31	251	32
rect	251	31	252	32
rect	252	31	253	32
rect	253	31	254	32
rect	254	31	255	32
rect	255	31	256	32
rect	256	31	257	32
rect	257	31	258	32
rect	258	31	259	32
rect	259	31	260	32
rect	260	31	261	32
rect	261	31	262	32
rect	262	31	263	32
rect	263	31	264	32
rect	264	31	265	32
rect	265	31	266	32
rect	266	31	267	32
rect	267	31	268	32
rect	268	31	269	32
rect	269	31	270	32
rect	270	31	271	32
rect	271	31	272	32
rect	272	31	273	32
rect	274	31	275	32
rect	275	31	276	32
rect	276	31	277	32
rect	277	31	278	32
rect	278	31	279	32
rect	279	31	280	32
rect	281	31	282	32
rect	282	31	283	32
rect	283	31	284	32
rect	284	31	285	32
rect	285	31	286	32
rect	286	31	287	32
rect	288	31	289	32
rect	289	31	290	32
rect	290	31	291	32
rect	291	31	292	32
rect	292	31	293	32
rect	293	31	294	32
rect	295	31	296	32
rect	296	31	297	32
rect	297	31	298	32
rect	298	31	299	32
rect	299	31	300	32
rect	300	31	301	32
rect	301	31	302	32
rect	302	31	303	32
rect	303	31	304	32
rect	304	31	305	32
rect	305	31	306	32
rect	306	31	307	32
rect	0	32	1	33
rect	1	32	2	33
rect	2	32	3	33
rect	3	32	4	33
rect	4	32	5	33
rect	5	32	6	33
rect	7	32	8	33
rect	8	32	9	33
rect	9	32	10	33
rect	10	32	11	33
rect	11	32	12	33
rect	12	32	13	33
rect	13	32	14	33
rect	14	32	15	33
rect	15	32	16	33
rect	16	32	17	33
rect	17	32	18	33
rect	18	32	19	33
rect	19	32	20	33
rect	20	32	21	33
rect	21	32	22	33
rect	23	32	24	33
rect	24	32	25	33
rect	25	32	26	33
rect	26	32	27	33
rect	27	32	28	33
rect	28	32	29	33
rect	29	32	30	33
rect	30	32	31	33
rect	31	32	32	33
rect	32	32	33	33
rect	33	32	34	33
rect	34	32	35	33
rect	35	32	36	33
rect	36	32	37	33
rect	37	32	38	33
rect	39	32	40	33
rect	40	32	41	33
rect	41	32	42	33
rect	42	32	43	33
rect	43	32	44	33
rect	44	32	45	33
rect	46	32	47	33
rect	47	32	48	33
rect	48	32	49	33
rect	49	32	50	33
rect	50	32	51	33
rect	51	32	52	33
rect	52	32	53	33
rect	53	32	54	33
rect	54	32	55	33
rect	55	32	56	33
rect	56	32	57	33
rect	57	32	58	33
rect	58	32	59	33
rect	59	32	60	33
rect	60	32	61	33
rect	61	32	62	33
rect	62	32	63	33
rect	63	32	64	33
rect	64	32	65	33
rect	65	32	66	33
rect	66	32	67	33
rect	67	32	68	33
rect	68	32	69	33
rect	69	32	70	33
rect	70	32	71	33
rect	71	32	72	33
rect	72	32	73	33
rect	73	32	74	33
rect	74	32	75	33
rect	75	32	76	33
rect	76	32	77	33
rect	77	32	78	33
rect	78	32	79	33
rect	80	32	81	33
rect	81	32	82	33
rect	82	32	83	33
rect	83	32	84	33
rect	84	32	85	33
rect	85	32	86	33
rect	87	32	88	33
rect	88	32	89	33
rect	89	32	90	33
rect	90	32	91	33
rect	91	32	92	33
rect	92	32	93	33
rect	94	32	95	33
rect	95	32	96	33
rect	96	32	97	33
rect	97	32	98	33
rect	98	32	99	33
rect	99	32	100	33
rect	101	32	102	33
rect	102	32	103	33
rect	103	32	104	33
rect	104	32	105	33
rect	105	32	106	33
rect	106	32	107	33
rect	107	32	108	33
rect	108	32	109	33
rect	109	32	110	33
rect	110	32	111	33
rect	111	32	112	33
rect	112	32	113	33
rect	113	32	114	33
rect	114	32	115	33
rect	115	32	116	33
rect	117	32	118	33
rect	118	32	119	33
rect	119	32	120	33
rect	120	32	121	33
rect	121	32	122	33
rect	122	32	123	33
rect	124	32	125	33
rect	125	32	126	33
rect	126	32	127	33
rect	127	32	128	33
rect	128	32	129	33
rect	129	32	130	33
rect	131	32	132	33
rect	132	32	133	33
rect	133	32	134	33
rect	134	32	135	33
rect	135	32	136	33
rect	136	32	137	33
rect	138	32	139	33
rect	139	32	140	33
rect	140	32	141	33
rect	141	32	142	33
rect	142	32	143	33
rect	143	32	144	33
rect	145	32	146	33
rect	146	32	147	33
rect	147	32	148	33
rect	148	32	149	33
rect	149	32	150	33
rect	150	32	151	33
rect	151	32	152	33
rect	152	32	153	33
rect	153	32	154	33
rect	154	32	155	33
rect	155	32	156	33
rect	156	32	157	33
rect	157	32	158	33
rect	158	32	159	33
rect	159	32	160	33
rect	160	32	161	33
rect	161	32	162	33
rect	162	32	163	33
rect	163	32	164	33
rect	164	32	165	33
rect	165	32	166	33
rect	166	32	167	33
rect	167	32	168	33
rect	168	32	169	33
rect	169	32	170	33
rect	170	32	171	33
rect	171	32	172	33
rect	172	32	173	33
rect	173	32	174	33
rect	174	32	175	33
rect	175	32	176	33
rect	176	32	177	33
rect	177	32	178	33
rect	178	32	179	33
rect	179	32	180	33
rect	180	32	181	33
rect	181	32	182	33
rect	182	32	183	33
rect	183	32	184	33
rect	184	32	185	33
rect	185	32	186	33
rect	186	32	187	33
rect	187	32	188	33
rect	188	32	189	33
rect	189	32	190	33
rect	190	32	191	33
rect	191	32	192	33
rect	192	32	193	33
rect	193	32	194	33
rect	194	32	195	33
rect	195	32	196	33
rect	196	32	197	33
rect	197	32	198	33
rect	198	32	199	33
rect	199	32	200	33
rect	200	32	201	33
rect	201	32	202	33
rect	202	32	203	33
rect	203	32	204	33
rect	204	32	205	33
rect	205	32	206	33
rect	206	32	207	33
rect	207	32	208	33
rect	208	32	209	33
rect	209	32	210	33
rect	210	32	211	33
rect	211	32	212	33
rect	212	32	213	33
rect	213	32	214	33
rect	214	32	215	33
rect	215	32	216	33
rect	216	32	217	33
rect	217	32	218	33
rect	218	32	219	33
rect	219	32	220	33
rect	220	32	221	33
rect	221	32	222	33
rect	222	32	223	33
rect	223	32	224	33
rect	224	32	225	33
rect	225	32	226	33
rect	226	32	227	33
rect	227	32	228	33
rect	228	32	229	33
rect	230	32	231	33
rect	231	32	232	33
rect	232	32	233	33
rect	233	32	234	33
rect	234	32	235	33
rect	235	32	236	33
rect	237	32	238	33
rect	238	32	239	33
rect	239	32	240	33
rect	240	32	241	33
rect	241	32	242	33
rect	242	32	243	33
rect	243	32	244	33
rect	244	32	245	33
rect	245	32	246	33
rect	246	32	247	33
rect	247	32	248	33
rect	248	32	249	33
rect	249	32	250	33
rect	250	32	251	33
rect	251	32	252	33
rect	252	32	253	33
rect	253	32	254	33
rect	254	32	255	33
rect	255	32	256	33
rect	256	32	257	33
rect	257	32	258	33
rect	258	32	259	33
rect	259	32	260	33
rect	260	32	261	33
rect	261	32	262	33
rect	262	32	263	33
rect	263	32	264	33
rect	264	32	265	33
rect	265	32	266	33
rect	266	32	267	33
rect	267	32	268	33
rect	268	32	269	33
rect	269	32	270	33
rect	270	32	271	33
rect	271	32	272	33
rect	272	32	273	33
rect	274	32	275	33
rect	275	32	276	33
rect	276	32	277	33
rect	277	32	278	33
rect	278	32	279	33
rect	279	32	280	33
rect	281	32	282	33
rect	282	32	283	33
rect	283	32	284	33
rect	284	32	285	33
rect	285	32	286	33
rect	286	32	287	33
rect	288	32	289	33
rect	289	32	290	33
rect	290	32	291	33
rect	291	32	292	33
rect	292	32	293	33
rect	293	32	294	33
rect	295	32	296	33
rect	296	32	297	33
rect	297	32	298	33
rect	298	32	299	33
rect	299	32	300	33
rect	300	32	301	33
rect	301	32	302	33
rect	302	32	303	33
rect	303	32	304	33
rect	304	32	305	33
rect	305	32	306	33
rect	306	32	307	33
rect	0	60	1	61
rect	1	60	2	61
rect	2	60	3	61
rect	3	60	4	61
rect	4	60	5	61
rect	5	60	6	61
rect	7	60	8	61
rect	8	60	9	61
rect	9	60	10	61
rect	10	60	11	61
rect	11	60	12	61
rect	12	60	13	61
rect	14	60	15	61
rect	15	60	16	61
rect	16	60	17	61
rect	17	60	18	61
rect	18	60	19	61
rect	19	60	20	61
rect	20	60	21	61
rect	21	60	22	61
rect	22	60	23	61
rect	23	60	24	61
rect	24	60	25	61
rect	25	60	26	61
rect	26	60	27	61
rect	27	60	28	61
rect	28	60	29	61
rect	30	60	31	61
rect	31	60	32	61
rect	32	60	33	61
rect	33	60	34	61
rect	34	60	35	61
rect	35	60	36	61
rect	36	60	37	61
rect	37	60	38	61
rect	38	60	39	61
rect	39	60	40	61
rect	40	60	41	61
rect	41	60	42	61
rect	42	60	43	61
rect	43	60	44	61
rect	44	60	45	61
rect	46	60	47	61
rect	47	60	48	61
rect	48	60	49	61
rect	49	60	50	61
rect	50	60	51	61
rect	51	60	52	61
rect	52	60	53	61
rect	53	60	54	61
rect	54	60	55	61
rect	55	60	56	61
rect	56	60	57	61
rect	57	60	58	61
rect	58	60	59	61
rect	59	60	60	61
rect	60	60	61	61
rect	61	60	62	61
rect	62	60	63	61
rect	63	60	64	61
rect	64	60	65	61
rect	65	60	66	61
rect	66	60	67	61
rect	67	60	68	61
rect	68	60	69	61
rect	69	60	70	61
rect	70	60	71	61
rect	71	60	72	61
rect	72	60	73	61
rect	73	60	74	61
rect	74	60	75	61
rect	75	60	76	61
rect	76	60	77	61
rect	77	60	78	61
rect	78	60	79	61
rect	79	60	80	61
rect	80	60	81	61
rect	81	60	82	61
rect	82	60	83	61
rect	83	60	84	61
rect	84	60	85	61
rect	85	60	86	61
rect	86	60	87	61
rect	87	60	88	61
rect	89	60	90	61
rect	90	60	91	61
rect	91	60	92	61
rect	92	60	93	61
rect	93	60	94	61
rect	94	60	95	61
rect	96	60	97	61
rect	97	60	98	61
rect	98	60	99	61
rect	99	60	100	61
rect	100	60	101	61
rect	101	60	102	61
rect	103	60	104	61
rect	104	60	105	61
rect	105	60	106	61
rect	106	60	107	61
rect	107	60	108	61
rect	108	60	109	61
rect	109	60	110	61
rect	110	60	111	61
rect	111	60	112	61
rect	112	60	113	61
rect	113	60	114	61
rect	114	60	115	61
rect	115	60	116	61
rect	116	60	117	61
rect	117	60	118	61
rect	118	60	119	61
rect	119	60	120	61
rect	120	60	121	61
rect	121	60	122	61
rect	122	60	123	61
rect	123	60	124	61
rect	124	60	125	61
rect	125	60	126	61
rect	126	60	127	61
rect	127	60	128	61
rect	128	60	129	61
rect	129	60	130	61
rect	130	60	131	61
rect	131	60	132	61
rect	132	60	133	61
rect	133	60	134	61
rect	134	60	135	61
rect	135	60	136	61
rect	137	60	138	61
rect	138	60	139	61
rect	139	60	140	61
rect	140	60	141	61
rect	141	60	142	61
rect	142	60	143	61
rect	144	60	145	61
rect	145	60	146	61
rect	146	60	147	61
rect	147	60	148	61
rect	148	60	149	61
rect	149	60	150	61
rect	151	60	152	61
rect	152	60	153	61
rect	153	60	154	61
rect	154	60	155	61
rect	155	60	156	61
rect	156	60	157	61
rect	157	60	158	61
rect	158	60	159	61
rect	159	60	160	61
rect	160	60	161	61
rect	161	60	162	61
rect	162	60	163	61
rect	163	60	164	61
rect	164	60	165	61
rect	165	60	166	61
rect	166	60	167	61
rect	167	60	168	61
rect	168	60	169	61
rect	169	60	170	61
rect	170	60	171	61
rect	171	60	172	61
rect	172	60	173	61
rect	173	60	174	61
rect	174	60	175	61
rect	175	60	176	61
rect	176	60	177	61
rect	177	60	178	61
rect	178	60	179	61
rect	179	60	180	61
rect	180	60	181	61
rect	181	60	182	61
rect	182	60	183	61
rect	183	60	184	61
rect	184	60	185	61
rect	185	60	186	61
rect	186	60	187	61
rect	187	60	188	61
rect	188	60	189	61
rect	189	60	190	61
rect	190	60	191	61
rect	191	60	192	61
rect	192	60	193	61
rect	193	60	194	61
rect	194	60	195	61
rect	195	60	196	61
rect	196	60	197	61
rect	197	60	198	61
rect	198	60	199	61
rect	199	60	200	61
rect	200	60	201	61
rect	201	60	202	61
rect	202	60	203	61
rect	203	60	204	61
rect	204	60	205	61
rect	205	60	206	61
rect	206	60	207	61
rect	207	60	208	61
rect	208	60	209	61
rect	209	60	210	61
rect	210	60	211	61
rect	211	60	212	61
rect	212	60	213	61
rect	213	60	214	61
rect	214	60	215	61
rect	215	60	216	61
rect	216	60	217	61
rect	217	60	218	61
rect	218	60	219	61
rect	219	60	220	61
rect	220	60	221	61
rect	221	60	222	61
rect	222	60	223	61
rect	223	60	224	61
rect	224	60	225	61
rect	225	60	226	61
rect	226	60	227	61
rect	227	60	228	61
rect	228	60	229	61
rect	229	60	230	61
rect	230	60	231	61
rect	231	60	232	61
rect	232	60	233	61
rect	233	60	234	61
rect	234	60	235	61
rect	235	60	236	61
rect	236	60	237	61
rect	237	60	238	61
rect	239	60	240	61
rect	240	60	241	61
rect	241	60	242	61
rect	242	60	243	61
rect	243	60	244	61
rect	244	60	245	61
rect	245	60	246	61
rect	246	60	247	61
rect	247	60	248	61
rect	248	60	249	61
rect	249	60	250	61
rect	250	60	251	61
rect	251	60	252	61
rect	252	60	253	61
rect	253	60	254	61
rect	254	60	255	61
rect	255	60	256	61
rect	256	60	257	61
rect	257	60	258	61
rect	258	60	259	61
rect	259	60	260	61
rect	260	60	261	61
rect	261	60	262	61
rect	262	60	263	61
rect	263	60	264	61
rect	264	60	265	61
rect	265	60	266	61
rect	266	60	267	61
rect	267	60	268	61
rect	268	60	269	61
rect	269	60	270	61
rect	270	60	271	61
rect	271	60	272	61
rect	272	60	273	61
rect	273	60	274	61
rect	274	60	275	61
rect	275	60	276	61
rect	276	60	277	61
rect	277	60	278	61
rect	278	60	279	61
rect	279	60	280	61
rect	280	60	281	61
rect	281	60	282	61
rect	282	60	283	61
rect	283	60	284	61
rect	284	60	285	61
rect	285	60	286	61
rect	286	60	287	61
rect	287	60	288	61
rect	288	60	289	61
rect	289	60	290	61
rect	290	60	291	61
rect	291	60	292	61
rect	292	60	293	61
rect	293	60	294	61
rect	294	60	295	61
rect	295	60	296	61
rect	296	60	297	61
rect	297	60	298	61
rect	298	60	299	61
rect	299	60	300	61
rect	300	60	301	61
rect	301	60	302	61
rect	302	60	303	61
rect	303	60	304	61
rect	304	60	305	61
rect	305	60	306	61
rect	306	60	307	61
rect	307	60	308	61
rect	308	60	309	61
rect	309	60	310	61
rect	310	60	311	61
rect	311	60	312	61
rect	312	60	313	61
rect	313	60	314	61
rect	314	60	315	61
rect	315	60	316	61
rect	316	60	317	61
rect	317	60	318	61
rect	318	60	319	61
rect	319	60	320	61
rect	320	60	321	61
rect	321	60	322	61
rect	322	60	323	61
rect	323	60	324	61
rect	324	60	325	61
rect	325	60	326	61
rect	326	60	327	61
rect	327	60	328	61
rect	328	60	329	61
rect	329	60	330	61
rect	330	60	331	61
rect	331	60	332	61
rect	332	60	333	61
rect	333	60	334	61
rect	334	60	335	61
rect	335	60	336	61
rect	336	60	337	61
rect	337	60	338	61
rect	338	60	339	61
rect	339	60	340	61
rect	340	60	341	61
rect	341	60	342	61
rect	342	60	343	61
rect	343	60	344	61
rect	344	60	345	61
rect	345	60	346	61
rect	346	60	347	61
rect	347	60	348	61
rect	348	60	349	61
rect	349	60	350	61
rect	350	60	351	61
rect	351	60	352	61
rect	352	60	353	61
rect	353	60	354	61
rect	354	60	355	61
rect	355	60	356	61
rect	356	60	357	61
rect	357	60	358	61
rect	358	60	359	61
rect	0	61	1	62
rect	1	61	2	62
rect	2	61	3	62
rect	3	61	4	62
rect	4	61	5	62
rect	5	61	6	62
rect	7	61	8	62
rect	8	61	9	62
rect	9	61	10	62
rect	10	61	11	62
rect	11	61	12	62
rect	12	61	13	62
rect	14	61	15	62
rect	15	61	16	62
rect	16	61	17	62
rect	17	61	18	62
rect	18	61	19	62
rect	19	61	20	62
rect	20	61	21	62
rect	21	61	22	62
rect	22	61	23	62
rect	23	61	24	62
rect	24	61	25	62
rect	25	61	26	62
rect	26	61	27	62
rect	27	61	28	62
rect	28	61	29	62
rect	30	61	31	62
rect	31	61	32	62
rect	32	61	33	62
rect	33	61	34	62
rect	34	61	35	62
rect	35	61	36	62
rect	36	61	37	62
rect	37	61	38	62
rect	38	61	39	62
rect	39	61	40	62
rect	40	61	41	62
rect	41	61	42	62
rect	42	61	43	62
rect	43	61	44	62
rect	44	61	45	62
rect	46	61	47	62
rect	47	61	48	62
rect	48	61	49	62
rect	49	61	50	62
rect	50	61	51	62
rect	51	61	52	62
rect	52	61	53	62
rect	53	61	54	62
rect	54	61	55	62
rect	55	61	56	62
rect	56	61	57	62
rect	57	61	58	62
rect	58	61	59	62
rect	59	61	60	62
rect	60	61	61	62
rect	61	61	62	62
rect	62	61	63	62
rect	63	61	64	62
rect	64	61	65	62
rect	65	61	66	62
rect	66	61	67	62
rect	67	61	68	62
rect	68	61	69	62
rect	69	61	70	62
rect	70	61	71	62
rect	71	61	72	62
rect	72	61	73	62
rect	73	61	74	62
rect	74	61	75	62
rect	75	61	76	62
rect	76	61	77	62
rect	77	61	78	62
rect	78	61	79	62
rect	79	61	80	62
rect	80	61	81	62
rect	81	61	82	62
rect	82	61	83	62
rect	83	61	84	62
rect	84	61	85	62
rect	85	61	86	62
rect	86	61	87	62
rect	87	61	88	62
rect	89	61	90	62
rect	90	61	91	62
rect	91	61	92	62
rect	92	61	93	62
rect	93	61	94	62
rect	94	61	95	62
rect	96	61	97	62
rect	97	61	98	62
rect	98	61	99	62
rect	99	61	100	62
rect	100	61	101	62
rect	101	61	102	62
rect	103	61	104	62
rect	104	61	105	62
rect	105	61	106	62
rect	106	61	107	62
rect	107	61	108	62
rect	108	61	109	62
rect	109	61	110	62
rect	110	61	111	62
rect	111	61	112	62
rect	112	61	113	62
rect	113	61	114	62
rect	114	61	115	62
rect	115	61	116	62
rect	116	61	117	62
rect	117	61	118	62
rect	118	61	119	62
rect	119	61	120	62
rect	120	61	121	62
rect	121	61	122	62
rect	122	61	123	62
rect	123	61	124	62
rect	124	61	125	62
rect	125	61	126	62
rect	126	61	127	62
rect	127	61	128	62
rect	128	61	129	62
rect	129	61	130	62
rect	130	61	131	62
rect	131	61	132	62
rect	132	61	133	62
rect	133	61	134	62
rect	134	61	135	62
rect	135	61	136	62
rect	137	61	138	62
rect	138	61	139	62
rect	139	61	140	62
rect	140	61	141	62
rect	141	61	142	62
rect	142	61	143	62
rect	144	61	145	62
rect	145	61	146	62
rect	146	61	147	62
rect	147	61	148	62
rect	148	61	149	62
rect	149	61	150	62
rect	151	61	152	62
rect	152	61	153	62
rect	153	61	154	62
rect	154	61	155	62
rect	155	61	156	62
rect	156	61	157	62
rect	157	61	158	62
rect	158	61	159	62
rect	159	61	160	62
rect	160	61	161	62
rect	161	61	162	62
rect	162	61	163	62
rect	163	61	164	62
rect	164	61	165	62
rect	165	61	166	62
rect	166	61	167	62
rect	167	61	168	62
rect	168	61	169	62
rect	169	61	170	62
rect	170	61	171	62
rect	171	61	172	62
rect	172	61	173	62
rect	173	61	174	62
rect	174	61	175	62
rect	175	61	176	62
rect	176	61	177	62
rect	177	61	178	62
rect	178	61	179	62
rect	179	61	180	62
rect	180	61	181	62
rect	181	61	182	62
rect	182	61	183	62
rect	183	61	184	62
rect	184	61	185	62
rect	185	61	186	62
rect	186	61	187	62
rect	187	61	188	62
rect	188	61	189	62
rect	189	61	190	62
rect	190	61	191	62
rect	191	61	192	62
rect	192	61	193	62
rect	193	61	194	62
rect	194	61	195	62
rect	195	61	196	62
rect	196	61	197	62
rect	197	61	198	62
rect	198	61	199	62
rect	199	61	200	62
rect	200	61	201	62
rect	201	61	202	62
rect	202	61	203	62
rect	203	61	204	62
rect	204	61	205	62
rect	205	61	206	62
rect	206	61	207	62
rect	207	61	208	62
rect	208	61	209	62
rect	209	61	210	62
rect	210	61	211	62
rect	211	61	212	62
rect	212	61	213	62
rect	213	61	214	62
rect	214	61	215	62
rect	215	61	216	62
rect	216	61	217	62
rect	217	61	218	62
rect	218	61	219	62
rect	219	61	220	62
rect	220	61	221	62
rect	221	61	222	62
rect	222	61	223	62
rect	223	61	224	62
rect	224	61	225	62
rect	225	61	226	62
rect	226	61	227	62
rect	227	61	228	62
rect	228	61	229	62
rect	229	61	230	62
rect	230	61	231	62
rect	231	61	232	62
rect	232	61	233	62
rect	233	61	234	62
rect	234	61	235	62
rect	235	61	236	62
rect	236	61	237	62
rect	237	61	238	62
rect	239	61	240	62
rect	240	61	241	62
rect	241	61	242	62
rect	242	61	243	62
rect	243	61	244	62
rect	244	61	245	62
rect	245	61	246	62
rect	246	61	247	62
rect	247	61	248	62
rect	248	61	249	62
rect	249	61	250	62
rect	250	61	251	62
rect	251	61	252	62
rect	252	61	253	62
rect	253	61	254	62
rect	254	61	255	62
rect	255	61	256	62
rect	256	61	257	62
rect	257	61	258	62
rect	258	61	259	62
rect	259	61	260	62
rect	260	61	261	62
rect	261	61	262	62
rect	262	61	263	62
rect	263	61	264	62
rect	264	61	265	62
rect	265	61	266	62
rect	266	61	267	62
rect	267	61	268	62
rect	268	61	269	62
rect	269	61	270	62
rect	270	61	271	62
rect	271	61	272	62
rect	272	61	273	62
rect	273	61	274	62
rect	274	61	275	62
rect	275	61	276	62
rect	276	61	277	62
rect	277	61	278	62
rect	278	61	279	62
rect	279	61	280	62
rect	280	61	281	62
rect	281	61	282	62
rect	282	61	283	62
rect	283	61	284	62
rect	284	61	285	62
rect	285	61	286	62
rect	286	61	287	62
rect	287	61	288	62
rect	288	61	289	62
rect	289	61	290	62
rect	290	61	291	62
rect	291	61	292	62
rect	292	61	293	62
rect	293	61	294	62
rect	294	61	295	62
rect	295	61	296	62
rect	296	61	297	62
rect	297	61	298	62
rect	298	61	299	62
rect	299	61	300	62
rect	300	61	301	62
rect	301	61	302	62
rect	302	61	303	62
rect	303	61	304	62
rect	304	61	305	62
rect	305	61	306	62
rect	306	61	307	62
rect	307	61	308	62
rect	308	61	309	62
rect	309	61	310	62
rect	310	61	311	62
rect	311	61	312	62
rect	312	61	313	62
rect	313	61	314	62
rect	314	61	315	62
rect	315	61	316	62
rect	316	61	317	62
rect	317	61	318	62
rect	318	61	319	62
rect	319	61	320	62
rect	320	61	321	62
rect	321	61	322	62
rect	322	61	323	62
rect	323	61	324	62
rect	324	61	325	62
rect	325	61	326	62
rect	326	61	327	62
rect	327	61	328	62
rect	328	61	329	62
rect	329	61	330	62
rect	330	61	331	62
rect	331	61	332	62
rect	332	61	333	62
rect	333	61	334	62
rect	334	61	335	62
rect	335	61	336	62
rect	336	61	337	62
rect	337	61	338	62
rect	338	61	339	62
rect	339	61	340	62
rect	340	61	341	62
rect	341	61	342	62
rect	342	61	343	62
rect	343	61	344	62
rect	344	61	345	62
rect	345	61	346	62
rect	346	61	347	62
rect	347	61	348	62
rect	348	61	349	62
rect	349	61	350	62
rect	350	61	351	62
rect	351	61	352	62
rect	352	61	353	62
rect	353	61	354	62
rect	354	61	355	62
rect	355	61	356	62
rect	356	61	357	62
rect	357	61	358	62
rect	358	61	359	62
rect	0	62	1	63
rect	1	62	2	63
rect	2	62	3	63
rect	3	62	4	63
rect	4	62	5	63
rect	5	62	6	63
rect	7	62	8	63
rect	8	62	9	63
rect	9	62	10	63
rect	10	62	11	63
rect	11	62	12	63
rect	12	62	13	63
rect	14	62	15	63
rect	15	62	16	63
rect	16	62	17	63
rect	17	62	18	63
rect	18	62	19	63
rect	19	62	20	63
rect	20	62	21	63
rect	21	62	22	63
rect	22	62	23	63
rect	23	62	24	63
rect	24	62	25	63
rect	25	62	26	63
rect	26	62	27	63
rect	27	62	28	63
rect	28	62	29	63
rect	30	62	31	63
rect	31	62	32	63
rect	32	62	33	63
rect	33	62	34	63
rect	34	62	35	63
rect	35	62	36	63
rect	36	62	37	63
rect	37	62	38	63
rect	38	62	39	63
rect	39	62	40	63
rect	40	62	41	63
rect	41	62	42	63
rect	42	62	43	63
rect	43	62	44	63
rect	44	62	45	63
rect	46	62	47	63
rect	47	62	48	63
rect	48	62	49	63
rect	49	62	50	63
rect	50	62	51	63
rect	51	62	52	63
rect	52	62	53	63
rect	53	62	54	63
rect	54	62	55	63
rect	55	62	56	63
rect	56	62	57	63
rect	57	62	58	63
rect	58	62	59	63
rect	59	62	60	63
rect	60	62	61	63
rect	61	62	62	63
rect	62	62	63	63
rect	63	62	64	63
rect	64	62	65	63
rect	65	62	66	63
rect	66	62	67	63
rect	67	62	68	63
rect	68	62	69	63
rect	69	62	70	63
rect	70	62	71	63
rect	71	62	72	63
rect	72	62	73	63
rect	73	62	74	63
rect	74	62	75	63
rect	75	62	76	63
rect	76	62	77	63
rect	77	62	78	63
rect	78	62	79	63
rect	79	62	80	63
rect	80	62	81	63
rect	81	62	82	63
rect	82	62	83	63
rect	83	62	84	63
rect	84	62	85	63
rect	85	62	86	63
rect	86	62	87	63
rect	87	62	88	63
rect	89	62	90	63
rect	90	62	91	63
rect	91	62	92	63
rect	92	62	93	63
rect	93	62	94	63
rect	94	62	95	63
rect	96	62	97	63
rect	97	62	98	63
rect	98	62	99	63
rect	99	62	100	63
rect	100	62	101	63
rect	101	62	102	63
rect	103	62	104	63
rect	104	62	105	63
rect	105	62	106	63
rect	106	62	107	63
rect	107	62	108	63
rect	108	62	109	63
rect	109	62	110	63
rect	110	62	111	63
rect	111	62	112	63
rect	112	62	113	63
rect	113	62	114	63
rect	114	62	115	63
rect	115	62	116	63
rect	116	62	117	63
rect	117	62	118	63
rect	118	62	119	63
rect	119	62	120	63
rect	120	62	121	63
rect	121	62	122	63
rect	122	62	123	63
rect	123	62	124	63
rect	124	62	125	63
rect	125	62	126	63
rect	126	62	127	63
rect	127	62	128	63
rect	128	62	129	63
rect	129	62	130	63
rect	130	62	131	63
rect	131	62	132	63
rect	132	62	133	63
rect	133	62	134	63
rect	134	62	135	63
rect	135	62	136	63
rect	137	62	138	63
rect	138	62	139	63
rect	139	62	140	63
rect	140	62	141	63
rect	141	62	142	63
rect	142	62	143	63
rect	144	62	145	63
rect	145	62	146	63
rect	146	62	147	63
rect	147	62	148	63
rect	148	62	149	63
rect	149	62	150	63
rect	151	62	152	63
rect	152	62	153	63
rect	153	62	154	63
rect	154	62	155	63
rect	155	62	156	63
rect	156	62	157	63
rect	157	62	158	63
rect	158	62	159	63
rect	159	62	160	63
rect	160	62	161	63
rect	161	62	162	63
rect	162	62	163	63
rect	163	62	164	63
rect	164	62	165	63
rect	165	62	166	63
rect	166	62	167	63
rect	167	62	168	63
rect	168	62	169	63
rect	169	62	170	63
rect	170	62	171	63
rect	171	62	172	63
rect	172	62	173	63
rect	173	62	174	63
rect	174	62	175	63
rect	175	62	176	63
rect	176	62	177	63
rect	177	62	178	63
rect	178	62	179	63
rect	179	62	180	63
rect	180	62	181	63
rect	181	62	182	63
rect	182	62	183	63
rect	183	62	184	63
rect	184	62	185	63
rect	185	62	186	63
rect	186	62	187	63
rect	187	62	188	63
rect	188	62	189	63
rect	189	62	190	63
rect	190	62	191	63
rect	191	62	192	63
rect	192	62	193	63
rect	193	62	194	63
rect	194	62	195	63
rect	195	62	196	63
rect	196	62	197	63
rect	197	62	198	63
rect	198	62	199	63
rect	199	62	200	63
rect	200	62	201	63
rect	201	62	202	63
rect	202	62	203	63
rect	203	62	204	63
rect	204	62	205	63
rect	205	62	206	63
rect	206	62	207	63
rect	207	62	208	63
rect	208	62	209	63
rect	209	62	210	63
rect	210	62	211	63
rect	211	62	212	63
rect	212	62	213	63
rect	213	62	214	63
rect	214	62	215	63
rect	215	62	216	63
rect	216	62	217	63
rect	217	62	218	63
rect	218	62	219	63
rect	219	62	220	63
rect	220	62	221	63
rect	221	62	222	63
rect	222	62	223	63
rect	223	62	224	63
rect	224	62	225	63
rect	225	62	226	63
rect	226	62	227	63
rect	227	62	228	63
rect	228	62	229	63
rect	229	62	230	63
rect	230	62	231	63
rect	231	62	232	63
rect	232	62	233	63
rect	233	62	234	63
rect	234	62	235	63
rect	235	62	236	63
rect	236	62	237	63
rect	237	62	238	63
rect	239	62	240	63
rect	240	62	241	63
rect	241	62	242	63
rect	242	62	243	63
rect	243	62	244	63
rect	244	62	245	63
rect	245	62	246	63
rect	246	62	247	63
rect	247	62	248	63
rect	248	62	249	63
rect	249	62	250	63
rect	250	62	251	63
rect	251	62	252	63
rect	252	62	253	63
rect	253	62	254	63
rect	254	62	255	63
rect	255	62	256	63
rect	256	62	257	63
rect	257	62	258	63
rect	258	62	259	63
rect	259	62	260	63
rect	260	62	261	63
rect	261	62	262	63
rect	262	62	263	63
rect	263	62	264	63
rect	264	62	265	63
rect	265	62	266	63
rect	266	62	267	63
rect	267	62	268	63
rect	268	62	269	63
rect	269	62	270	63
rect	270	62	271	63
rect	271	62	272	63
rect	272	62	273	63
rect	273	62	274	63
rect	274	62	275	63
rect	275	62	276	63
rect	276	62	277	63
rect	277	62	278	63
rect	278	62	279	63
rect	279	62	280	63
rect	280	62	281	63
rect	281	62	282	63
rect	282	62	283	63
rect	283	62	284	63
rect	284	62	285	63
rect	285	62	286	63
rect	286	62	287	63
rect	287	62	288	63
rect	288	62	289	63
rect	289	62	290	63
rect	290	62	291	63
rect	291	62	292	63
rect	292	62	293	63
rect	293	62	294	63
rect	294	62	295	63
rect	295	62	296	63
rect	296	62	297	63
rect	297	62	298	63
rect	298	62	299	63
rect	299	62	300	63
rect	300	62	301	63
rect	301	62	302	63
rect	302	62	303	63
rect	303	62	304	63
rect	304	62	305	63
rect	305	62	306	63
rect	306	62	307	63
rect	307	62	308	63
rect	308	62	309	63
rect	309	62	310	63
rect	310	62	311	63
rect	311	62	312	63
rect	312	62	313	63
rect	313	62	314	63
rect	314	62	315	63
rect	315	62	316	63
rect	316	62	317	63
rect	317	62	318	63
rect	318	62	319	63
rect	319	62	320	63
rect	320	62	321	63
rect	321	62	322	63
rect	322	62	323	63
rect	323	62	324	63
rect	324	62	325	63
rect	325	62	326	63
rect	326	62	327	63
rect	327	62	328	63
rect	328	62	329	63
rect	329	62	330	63
rect	330	62	331	63
rect	331	62	332	63
rect	332	62	333	63
rect	333	62	334	63
rect	334	62	335	63
rect	335	62	336	63
rect	336	62	337	63
rect	337	62	338	63
rect	338	62	339	63
rect	339	62	340	63
rect	340	62	341	63
rect	341	62	342	63
rect	342	62	343	63
rect	343	62	344	63
rect	344	62	345	63
rect	345	62	346	63
rect	346	62	347	63
rect	347	62	348	63
rect	348	62	349	63
rect	349	62	350	63
rect	350	62	351	63
rect	351	62	352	63
rect	352	62	353	63
rect	353	62	354	63
rect	354	62	355	63
rect	355	62	356	63
rect	356	62	357	63
rect	357	62	358	63
rect	358	62	359	63
rect	0	63	1	64
rect	1	63	2	64
rect	2	63	3	64
rect	3	63	4	64
rect	4	63	5	64
rect	5	63	6	64
rect	7	63	8	64
rect	8	63	9	64
rect	9	63	10	64
rect	10	63	11	64
rect	11	63	12	64
rect	12	63	13	64
rect	14	63	15	64
rect	15	63	16	64
rect	16	63	17	64
rect	17	63	18	64
rect	18	63	19	64
rect	19	63	20	64
rect	20	63	21	64
rect	21	63	22	64
rect	22	63	23	64
rect	23	63	24	64
rect	24	63	25	64
rect	25	63	26	64
rect	26	63	27	64
rect	27	63	28	64
rect	28	63	29	64
rect	30	63	31	64
rect	31	63	32	64
rect	32	63	33	64
rect	33	63	34	64
rect	34	63	35	64
rect	35	63	36	64
rect	36	63	37	64
rect	37	63	38	64
rect	38	63	39	64
rect	39	63	40	64
rect	40	63	41	64
rect	41	63	42	64
rect	42	63	43	64
rect	43	63	44	64
rect	44	63	45	64
rect	46	63	47	64
rect	47	63	48	64
rect	48	63	49	64
rect	49	63	50	64
rect	50	63	51	64
rect	51	63	52	64
rect	52	63	53	64
rect	53	63	54	64
rect	54	63	55	64
rect	55	63	56	64
rect	56	63	57	64
rect	57	63	58	64
rect	58	63	59	64
rect	59	63	60	64
rect	60	63	61	64
rect	61	63	62	64
rect	62	63	63	64
rect	63	63	64	64
rect	64	63	65	64
rect	65	63	66	64
rect	66	63	67	64
rect	67	63	68	64
rect	68	63	69	64
rect	69	63	70	64
rect	70	63	71	64
rect	71	63	72	64
rect	72	63	73	64
rect	73	63	74	64
rect	74	63	75	64
rect	75	63	76	64
rect	76	63	77	64
rect	77	63	78	64
rect	78	63	79	64
rect	79	63	80	64
rect	80	63	81	64
rect	81	63	82	64
rect	82	63	83	64
rect	83	63	84	64
rect	84	63	85	64
rect	85	63	86	64
rect	86	63	87	64
rect	87	63	88	64
rect	89	63	90	64
rect	90	63	91	64
rect	91	63	92	64
rect	92	63	93	64
rect	93	63	94	64
rect	94	63	95	64
rect	96	63	97	64
rect	97	63	98	64
rect	98	63	99	64
rect	99	63	100	64
rect	100	63	101	64
rect	101	63	102	64
rect	103	63	104	64
rect	104	63	105	64
rect	105	63	106	64
rect	106	63	107	64
rect	107	63	108	64
rect	108	63	109	64
rect	109	63	110	64
rect	110	63	111	64
rect	111	63	112	64
rect	112	63	113	64
rect	113	63	114	64
rect	114	63	115	64
rect	115	63	116	64
rect	116	63	117	64
rect	117	63	118	64
rect	118	63	119	64
rect	119	63	120	64
rect	120	63	121	64
rect	121	63	122	64
rect	122	63	123	64
rect	123	63	124	64
rect	124	63	125	64
rect	125	63	126	64
rect	126	63	127	64
rect	127	63	128	64
rect	128	63	129	64
rect	129	63	130	64
rect	130	63	131	64
rect	131	63	132	64
rect	132	63	133	64
rect	133	63	134	64
rect	134	63	135	64
rect	135	63	136	64
rect	137	63	138	64
rect	138	63	139	64
rect	139	63	140	64
rect	140	63	141	64
rect	141	63	142	64
rect	142	63	143	64
rect	144	63	145	64
rect	145	63	146	64
rect	146	63	147	64
rect	147	63	148	64
rect	148	63	149	64
rect	149	63	150	64
rect	151	63	152	64
rect	152	63	153	64
rect	153	63	154	64
rect	154	63	155	64
rect	155	63	156	64
rect	156	63	157	64
rect	157	63	158	64
rect	158	63	159	64
rect	159	63	160	64
rect	160	63	161	64
rect	161	63	162	64
rect	162	63	163	64
rect	163	63	164	64
rect	164	63	165	64
rect	165	63	166	64
rect	166	63	167	64
rect	167	63	168	64
rect	168	63	169	64
rect	169	63	170	64
rect	170	63	171	64
rect	171	63	172	64
rect	172	63	173	64
rect	173	63	174	64
rect	174	63	175	64
rect	175	63	176	64
rect	176	63	177	64
rect	177	63	178	64
rect	178	63	179	64
rect	179	63	180	64
rect	180	63	181	64
rect	181	63	182	64
rect	182	63	183	64
rect	183	63	184	64
rect	184	63	185	64
rect	185	63	186	64
rect	186	63	187	64
rect	187	63	188	64
rect	188	63	189	64
rect	189	63	190	64
rect	190	63	191	64
rect	191	63	192	64
rect	192	63	193	64
rect	193	63	194	64
rect	194	63	195	64
rect	195	63	196	64
rect	196	63	197	64
rect	197	63	198	64
rect	198	63	199	64
rect	199	63	200	64
rect	200	63	201	64
rect	201	63	202	64
rect	202	63	203	64
rect	203	63	204	64
rect	204	63	205	64
rect	205	63	206	64
rect	206	63	207	64
rect	207	63	208	64
rect	208	63	209	64
rect	209	63	210	64
rect	210	63	211	64
rect	211	63	212	64
rect	212	63	213	64
rect	213	63	214	64
rect	214	63	215	64
rect	215	63	216	64
rect	216	63	217	64
rect	217	63	218	64
rect	218	63	219	64
rect	219	63	220	64
rect	220	63	221	64
rect	221	63	222	64
rect	222	63	223	64
rect	223	63	224	64
rect	224	63	225	64
rect	225	63	226	64
rect	226	63	227	64
rect	227	63	228	64
rect	228	63	229	64
rect	229	63	230	64
rect	230	63	231	64
rect	231	63	232	64
rect	232	63	233	64
rect	233	63	234	64
rect	234	63	235	64
rect	235	63	236	64
rect	236	63	237	64
rect	237	63	238	64
rect	239	63	240	64
rect	240	63	241	64
rect	241	63	242	64
rect	242	63	243	64
rect	243	63	244	64
rect	244	63	245	64
rect	245	63	246	64
rect	246	63	247	64
rect	247	63	248	64
rect	248	63	249	64
rect	249	63	250	64
rect	250	63	251	64
rect	251	63	252	64
rect	252	63	253	64
rect	253	63	254	64
rect	254	63	255	64
rect	255	63	256	64
rect	256	63	257	64
rect	257	63	258	64
rect	258	63	259	64
rect	259	63	260	64
rect	260	63	261	64
rect	261	63	262	64
rect	262	63	263	64
rect	263	63	264	64
rect	264	63	265	64
rect	265	63	266	64
rect	266	63	267	64
rect	267	63	268	64
rect	268	63	269	64
rect	269	63	270	64
rect	270	63	271	64
rect	271	63	272	64
rect	272	63	273	64
rect	273	63	274	64
rect	274	63	275	64
rect	275	63	276	64
rect	276	63	277	64
rect	277	63	278	64
rect	278	63	279	64
rect	279	63	280	64
rect	280	63	281	64
rect	281	63	282	64
rect	282	63	283	64
rect	283	63	284	64
rect	284	63	285	64
rect	285	63	286	64
rect	286	63	287	64
rect	287	63	288	64
rect	288	63	289	64
rect	289	63	290	64
rect	290	63	291	64
rect	291	63	292	64
rect	292	63	293	64
rect	293	63	294	64
rect	294	63	295	64
rect	295	63	296	64
rect	296	63	297	64
rect	297	63	298	64
rect	298	63	299	64
rect	299	63	300	64
rect	300	63	301	64
rect	301	63	302	64
rect	302	63	303	64
rect	303	63	304	64
rect	304	63	305	64
rect	305	63	306	64
rect	306	63	307	64
rect	307	63	308	64
rect	308	63	309	64
rect	309	63	310	64
rect	310	63	311	64
rect	311	63	312	64
rect	312	63	313	64
rect	313	63	314	64
rect	314	63	315	64
rect	315	63	316	64
rect	316	63	317	64
rect	317	63	318	64
rect	318	63	319	64
rect	319	63	320	64
rect	320	63	321	64
rect	321	63	322	64
rect	322	63	323	64
rect	323	63	324	64
rect	324	63	325	64
rect	325	63	326	64
rect	326	63	327	64
rect	327	63	328	64
rect	328	63	329	64
rect	329	63	330	64
rect	330	63	331	64
rect	331	63	332	64
rect	332	63	333	64
rect	333	63	334	64
rect	334	63	335	64
rect	335	63	336	64
rect	336	63	337	64
rect	337	63	338	64
rect	338	63	339	64
rect	339	63	340	64
rect	340	63	341	64
rect	341	63	342	64
rect	342	63	343	64
rect	343	63	344	64
rect	344	63	345	64
rect	345	63	346	64
rect	346	63	347	64
rect	347	63	348	64
rect	348	63	349	64
rect	349	63	350	64
rect	350	63	351	64
rect	351	63	352	64
rect	352	63	353	64
rect	353	63	354	64
rect	354	63	355	64
rect	355	63	356	64
rect	356	63	357	64
rect	357	63	358	64
rect	358	63	359	64
rect	0	64	1	65
rect	1	64	2	65
rect	2	64	3	65
rect	3	64	4	65
rect	4	64	5	65
rect	5	64	6	65
rect	7	64	8	65
rect	8	64	9	65
rect	9	64	10	65
rect	10	64	11	65
rect	11	64	12	65
rect	12	64	13	65
rect	14	64	15	65
rect	15	64	16	65
rect	16	64	17	65
rect	17	64	18	65
rect	18	64	19	65
rect	19	64	20	65
rect	20	64	21	65
rect	21	64	22	65
rect	22	64	23	65
rect	23	64	24	65
rect	24	64	25	65
rect	25	64	26	65
rect	26	64	27	65
rect	27	64	28	65
rect	28	64	29	65
rect	30	64	31	65
rect	31	64	32	65
rect	32	64	33	65
rect	33	64	34	65
rect	34	64	35	65
rect	35	64	36	65
rect	36	64	37	65
rect	37	64	38	65
rect	38	64	39	65
rect	39	64	40	65
rect	40	64	41	65
rect	41	64	42	65
rect	42	64	43	65
rect	43	64	44	65
rect	44	64	45	65
rect	46	64	47	65
rect	47	64	48	65
rect	48	64	49	65
rect	49	64	50	65
rect	50	64	51	65
rect	51	64	52	65
rect	52	64	53	65
rect	53	64	54	65
rect	54	64	55	65
rect	55	64	56	65
rect	56	64	57	65
rect	57	64	58	65
rect	58	64	59	65
rect	59	64	60	65
rect	60	64	61	65
rect	61	64	62	65
rect	62	64	63	65
rect	63	64	64	65
rect	64	64	65	65
rect	65	64	66	65
rect	66	64	67	65
rect	67	64	68	65
rect	68	64	69	65
rect	69	64	70	65
rect	70	64	71	65
rect	71	64	72	65
rect	72	64	73	65
rect	73	64	74	65
rect	74	64	75	65
rect	75	64	76	65
rect	76	64	77	65
rect	77	64	78	65
rect	78	64	79	65
rect	79	64	80	65
rect	80	64	81	65
rect	81	64	82	65
rect	82	64	83	65
rect	83	64	84	65
rect	84	64	85	65
rect	85	64	86	65
rect	86	64	87	65
rect	87	64	88	65
rect	89	64	90	65
rect	90	64	91	65
rect	91	64	92	65
rect	92	64	93	65
rect	93	64	94	65
rect	94	64	95	65
rect	96	64	97	65
rect	97	64	98	65
rect	98	64	99	65
rect	99	64	100	65
rect	100	64	101	65
rect	101	64	102	65
rect	103	64	104	65
rect	104	64	105	65
rect	105	64	106	65
rect	106	64	107	65
rect	107	64	108	65
rect	108	64	109	65
rect	109	64	110	65
rect	110	64	111	65
rect	111	64	112	65
rect	112	64	113	65
rect	113	64	114	65
rect	114	64	115	65
rect	115	64	116	65
rect	116	64	117	65
rect	117	64	118	65
rect	118	64	119	65
rect	119	64	120	65
rect	120	64	121	65
rect	121	64	122	65
rect	122	64	123	65
rect	123	64	124	65
rect	124	64	125	65
rect	125	64	126	65
rect	126	64	127	65
rect	127	64	128	65
rect	128	64	129	65
rect	129	64	130	65
rect	130	64	131	65
rect	131	64	132	65
rect	132	64	133	65
rect	133	64	134	65
rect	134	64	135	65
rect	135	64	136	65
rect	137	64	138	65
rect	138	64	139	65
rect	139	64	140	65
rect	140	64	141	65
rect	141	64	142	65
rect	142	64	143	65
rect	144	64	145	65
rect	145	64	146	65
rect	146	64	147	65
rect	147	64	148	65
rect	148	64	149	65
rect	149	64	150	65
rect	151	64	152	65
rect	152	64	153	65
rect	153	64	154	65
rect	154	64	155	65
rect	155	64	156	65
rect	156	64	157	65
rect	157	64	158	65
rect	158	64	159	65
rect	159	64	160	65
rect	160	64	161	65
rect	161	64	162	65
rect	162	64	163	65
rect	163	64	164	65
rect	164	64	165	65
rect	165	64	166	65
rect	166	64	167	65
rect	167	64	168	65
rect	168	64	169	65
rect	169	64	170	65
rect	170	64	171	65
rect	171	64	172	65
rect	172	64	173	65
rect	173	64	174	65
rect	174	64	175	65
rect	175	64	176	65
rect	176	64	177	65
rect	177	64	178	65
rect	178	64	179	65
rect	179	64	180	65
rect	180	64	181	65
rect	181	64	182	65
rect	182	64	183	65
rect	183	64	184	65
rect	184	64	185	65
rect	185	64	186	65
rect	186	64	187	65
rect	187	64	188	65
rect	188	64	189	65
rect	189	64	190	65
rect	190	64	191	65
rect	191	64	192	65
rect	192	64	193	65
rect	193	64	194	65
rect	194	64	195	65
rect	195	64	196	65
rect	196	64	197	65
rect	197	64	198	65
rect	198	64	199	65
rect	199	64	200	65
rect	200	64	201	65
rect	201	64	202	65
rect	202	64	203	65
rect	203	64	204	65
rect	204	64	205	65
rect	205	64	206	65
rect	206	64	207	65
rect	207	64	208	65
rect	208	64	209	65
rect	209	64	210	65
rect	210	64	211	65
rect	211	64	212	65
rect	212	64	213	65
rect	213	64	214	65
rect	214	64	215	65
rect	215	64	216	65
rect	216	64	217	65
rect	217	64	218	65
rect	218	64	219	65
rect	219	64	220	65
rect	220	64	221	65
rect	221	64	222	65
rect	222	64	223	65
rect	223	64	224	65
rect	224	64	225	65
rect	225	64	226	65
rect	226	64	227	65
rect	227	64	228	65
rect	228	64	229	65
rect	229	64	230	65
rect	230	64	231	65
rect	231	64	232	65
rect	232	64	233	65
rect	233	64	234	65
rect	234	64	235	65
rect	235	64	236	65
rect	236	64	237	65
rect	237	64	238	65
rect	239	64	240	65
rect	240	64	241	65
rect	241	64	242	65
rect	242	64	243	65
rect	243	64	244	65
rect	244	64	245	65
rect	245	64	246	65
rect	246	64	247	65
rect	247	64	248	65
rect	248	64	249	65
rect	249	64	250	65
rect	250	64	251	65
rect	251	64	252	65
rect	252	64	253	65
rect	253	64	254	65
rect	254	64	255	65
rect	255	64	256	65
rect	256	64	257	65
rect	257	64	258	65
rect	258	64	259	65
rect	259	64	260	65
rect	260	64	261	65
rect	261	64	262	65
rect	262	64	263	65
rect	263	64	264	65
rect	264	64	265	65
rect	265	64	266	65
rect	266	64	267	65
rect	267	64	268	65
rect	268	64	269	65
rect	269	64	270	65
rect	270	64	271	65
rect	271	64	272	65
rect	272	64	273	65
rect	273	64	274	65
rect	274	64	275	65
rect	275	64	276	65
rect	276	64	277	65
rect	277	64	278	65
rect	278	64	279	65
rect	279	64	280	65
rect	280	64	281	65
rect	281	64	282	65
rect	282	64	283	65
rect	283	64	284	65
rect	284	64	285	65
rect	285	64	286	65
rect	286	64	287	65
rect	287	64	288	65
rect	288	64	289	65
rect	289	64	290	65
rect	290	64	291	65
rect	291	64	292	65
rect	292	64	293	65
rect	293	64	294	65
rect	294	64	295	65
rect	295	64	296	65
rect	296	64	297	65
rect	297	64	298	65
rect	298	64	299	65
rect	299	64	300	65
rect	300	64	301	65
rect	301	64	302	65
rect	302	64	303	65
rect	303	64	304	65
rect	304	64	305	65
rect	305	64	306	65
rect	306	64	307	65
rect	307	64	308	65
rect	308	64	309	65
rect	309	64	310	65
rect	310	64	311	65
rect	311	64	312	65
rect	312	64	313	65
rect	313	64	314	65
rect	314	64	315	65
rect	315	64	316	65
rect	316	64	317	65
rect	317	64	318	65
rect	318	64	319	65
rect	319	64	320	65
rect	320	64	321	65
rect	321	64	322	65
rect	322	64	323	65
rect	323	64	324	65
rect	324	64	325	65
rect	325	64	326	65
rect	326	64	327	65
rect	327	64	328	65
rect	328	64	329	65
rect	329	64	330	65
rect	330	64	331	65
rect	331	64	332	65
rect	332	64	333	65
rect	333	64	334	65
rect	334	64	335	65
rect	335	64	336	65
rect	336	64	337	65
rect	337	64	338	65
rect	338	64	339	65
rect	339	64	340	65
rect	340	64	341	65
rect	341	64	342	65
rect	342	64	343	65
rect	343	64	344	65
rect	344	64	345	65
rect	345	64	346	65
rect	346	64	347	65
rect	347	64	348	65
rect	348	64	349	65
rect	349	64	350	65
rect	350	64	351	65
rect	351	64	352	65
rect	352	64	353	65
rect	353	64	354	65
rect	354	64	355	65
rect	355	64	356	65
rect	356	64	357	65
rect	357	64	358	65
rect	358	64	359	65
rect	0	65	1	66
rect	1	65	2	66
rect	2	65	3	66
rect	3	65	4	66
rect	4	65	5	66
rect	5	65	6	66
rect	7	65	8	66
rect	8	65	9	66
rect	9	65	10	66
rect	10	65	11	66
rect	11	65	12	66
rect	12	65	13	66
rect	14	65	15	66
rect	15	65	16	66
rect	16	65	17	66
rect	17	65	18	66
rect	18	65	19	66
rect	19	65	20	66
rect	20	65	21	66
rect	21	65	22	66
rect	22	65	23	66
rect	23	65	24	66
rect	24	65	25	66
rect	25	65	26	66
rect	26	65	27	66
rect	27	65	28	66
rect	28	65	29	66
rect	30	65	31	66
rect	31	65	32	66
rect	32	65	33	66
rect	33	65	34	66
rect	34	65	35	66
rect	35	65	36	66
rect	36	65	37	66
rect	37	65	38	66
rect	38	65	39	66
rect	39	65	40	66
rect	40	65	41	66
rect	41	65	42	66
rect	42	65	43	66
rect	43	65	44	66
rect	44	65	45	66
rect	46	65	47	66
rect	47	65	48	66
rect	48	65	49	66
rect	49	65	50	66
rect	50	65	51	66
rect	51	65	52	66
rect	52	65	53	66
rect	53	65	54	66
rect	54	65	55	66
rect	55	65	56	66
rect	56	65	57	66
rect	57	65	58	66
rect	58	65	59	66
rect	59	65	60	66
rect	60	65	61	66
rect	61	65	62	66
rect	62	65	63	66
rect	63	65	64	66
rect	64	65	65	66
rect	65	65	66	66
rect	66	65	67	66
rect	67	65	68	66
rect	68	65	69	66
rect	69	65	70	66
rect	70	65	71	66
rect	71	65	72	66
rect	72	65	73	66
rect	73	65	74	66
rect	74	65	75	66
rect	75	65	76	66
rect	76	65	77	66
rect	77	65	78	66
rect	78	65	79	66
rect	79	65	80	66
rect	80	65	81	66
rect	81	65	82	66
rect	82	65	83	66
rect	83	65	84	66
rect	84	65	85	66
rect	85	65	86	66
rect	86	65	87	66
rect	87	65	88	66
rect	89	65	90	66
rect	90	65	91	66
rect	91	65	92	66
rect	92	65	93	66
rect	93	65	94	66
rect	94	65	95	66
rect	96	65	97	66
rect	97	65	98	66
rect	98	65	99	66
rect	99	65	100	66
rect	100	65	101	66
rect	101	65	102	66
rect	103	65	104	66
rect	104	65	105	66
rect	105	65	106	66
rect	106	65	107	66
rect	107	65	108	66
rect	108	65	109	66
rect	109	65	110	66
rect	110	65	111	66
rect	111	65	112	66
rect	112	65	113	66
rect	113	65	114	66
rect	114	65	115	66
rect	115	65	116	66
rect	116	65	117	66
rect	117	65	118	66
rect	118	65	119	66
rect	119	65	120	66
rect	120	65	121	66
rect	121	65	122	66
rect	122	65	123	66
rect	123	65	124	66
rect	124	65	125	66
rect	125	65	126	66
rect	126	65	127	66
rect	127	65	128	66
rect	128	65	129	66
rect	129	65	130	66
rect	130	65	131	66
rect	131	65	132	66
rect	132	65	133	66
rect	133	65	134	66
rect	134	65	135	66
rect	135	65	136	66
rect	137	65	138	66
rect	138	65	139	66
rect	139	65	140	66
rect	140	65	141	66
rect	141	65	142	66
rect	142	65	143	66
rect	144	65	145	66
rect	145	65	146	66
rect	146	65	147	66
rect	147	65	148	66
rect	148	65	149	66
rect	149	65	150	66
rect	151	65	152	66
rect	152	65	153	66
rect	153	65	154	66
rect	154	65	155	66
rect	155	65	156	66
rect	156	65	157	66
rect	157	65	158	66
rect	158	65	159	66
rect	159	65	160	66
rect	160	65	161	66
rect	161	65	162	66
rect	162	65	163	66
rect	163	65	164	66
rect	164	65	165	66
rect	165	65	166	66
rect	166	65	167	66
rect	167	65	168	66
rect	168	65	169	66
rect	169	65	170	66
rect	170	65	171	66
rect	171	65	172	66
rect	172	65	173	66
rect	173	65	174	66
rect	174	65	175	66
rect	175	65	176	66
rect	176	65	177	66
rect	177	65	178	66
rect	178	65	179	66
rect	179	65	180	66
rect	180	65	181	66
rect	181	65	182	66
rect	182	65	183	66
rect	183	65	184	66
rect	184	65	185	66
rect	185	65	186	66
rect	186	65	187	66
rect	187	65	188	66
rect	188	65	189	66
rect	189	65	190	66
rect	190	65	191	66
rect	191	65	192	66
rect	192	65	193	66
rect	193	65	194	66
rect	194	65	195	66
rect	195	65	196	66
rect	196	65	197	66
rect	197	65	198	66
rect	198	65	199	66
rect	199	65	200	66
rect	200	65	201	66
rect	201	65	202	66
rect	202	65	203	66
rect	203	65	204	66
rect	204	65	205	66
rect	205	65	206	66
rect	206	65	207	66
rect	207	65	208	66
rect	208	65	209	66
rect	209	65	210	66
rect	210	65	211	66
rect	211	65	212	66
rect	212	65	213	66
rect	213	65	214	66
rect	214	65	215	66
rect	215	65	216	66
rect	216	65	217	66
rect	217	65	218	66
rect	218	65	219	66
rect	219	65	220	66
rect	220	65	221	66
rect	221	65	222	66
rect	222	65	223	66
rect	223	65	224	66
rect	224	65	225	66
rect	225	65	226	66
rect	226	65	227	66
rect	227	65	228	66
rect	228	65	229	66
rect	229	65	230	66
rect	230	65	231	66
rect	231	65	232	66
rect	232	65	233	66
rect	233	65	234	66
rect	234	65	235	66
rect	235	65	236	66
rect	236	65	237	66
rect	237	65	238	66
rect	239	65	240	66
rect	240	65	241	66
rect	241	65	242	66
rect	242	65	243	66
rect	243	65	244	66
rect	244	65	245	66
rect	245	65	246	66
rect	246	65	247	66
rect	247	65	248	66
rect	248	65	249	66
rect	249	65	250	66
rect	250	65	251	66
rect	251	65	252	66
rect	252	65	253	66
rect	253	65	254	66
rect	254	65	255	66
rect	255	65	256	66
rect	256	65	257	66
rect	257	65	258	66
rect	258	65	259	66
rect	259	65	260	66
rect	260	65	261	66
rect	261	65	262	66
rect	262	65	263	66
rect	263	65	264	66
rect	264	65	265	66
rect	265	65	266	66
rect	266	65	267	66
rect	267	65	268	66
rect	268	65	269	66
rect	269	65	270	66
rect	270	65	271	66
rect	271	65	272	66
rect	272	65	273	66
rect	273	65	274	66
rect	274	65	275	66
rect	275	65	276	66
rect	276	65	277	66
rect	277	65	278	66
rect	278	65	279	66
rect	279	65	280	66
rect	280	65	281	66
rect	281	65	282	66
rect	282	65	283	66
rect	283	65	284	66
rect	284	65	285	66
rect	285	65	286	66
rect	286	65	287	66
rect	287	65	288	66
rect	288	65	289	66
rect	289	65	290	66
rect	290	65	291	66
rect	291	65	292	66
rect	292	65	293	66
rect	293	65	294	66
rect	294	65	295	66
rect	295	65	296	66
rect	296	65	297	66
rect	297	65	298	66
rect	298	65	299	66
rect	299	65	300	66
rect	300	65	301	66
rect	301	65	302	66
rect	302	65	303	66
rect	303	65	304	66
rect	304	65	305	66
rect	305	65	306	66
rect	306	65	307	66
rect	307	65	308	66
rect	308	65	309	66
rect	309	65	310	66
rect	310	65	311	66
rect	311	65	312	66
rect	312	65	313	66
rect	313	65	314	66
rect	314	65	315	66
rect	315	65	316	66
rect	316	65	317	66
rect	317	65	318	66
rect	318	65	319	66
rect	319	65	320	66
rect	320	65	321	66
rect	321	65	322	66
rect	322	65	323	66
rect	323	65	324	66
rect	324	65	325	66
rect	325	65	326	66
rect	326	65	327	66
rect	327	65	328	66
rect	328	65	329	66
rect	329	65	330	66
rect	330	65	331	66
rect	331	65	332	66
rect	332	65	333	66
rect	333	65	334	66
rect	334	65	335	66
rect	335	65	336	66
rect	336	65	337	66
rect	337	65	338	66
rect	338	65	339	66
rect	339	65	340	66
rect	340	65	341	66
rect	341	65	342	66
rect	342	65	343	66
rect	343	65	344	66
rect	344	65	345	66
rect	345	65	346	66
rect	346	65	347	66
rect	347	65	348	66
rect	348	65	349	66
rect	349	65	350	66
rect	350	65	351	66
rect	351	65	352	66
rect	352	65	353	66
rect	353	65	354	66
rect	354	65	355	66
rect	355	65	356	66
rect	356	65	357	66
rect	357	65	358	66
rect	358	65	359	66
rect	0	97	1	98
rect	1	97	2	98
rect	2	97	3	98
rect	3	97	4	98
rect	4	97	5	98
rect	5	97	6	98
rect	7	97	8	98
rect	8	97	9	98
rect	9	97	10	98
rect	10	97	11	98
rect	11	97	12	98
rect	12	97	13	98
rect	14	97	15	98
rect	15	97	16	98
rect	16	97	17	98
rect	17	97	18	98
rect	18	97	19	98
rect	19	97	20	98
rect	21	97	22	98
rect	22	97	23	98
rect	23	97	24	98
rect	24	97	25	98
rect	25	97	26	98
rect	26	97	27	98
rect	27	97	28	98
rect	28	97	29	98
rect	29	97	30	98
rect	30	97	31	98
rect	31	97	32	98
rect	32	97	33	98
rect	33	97	34	98
rect	34	97	35	98
rect	35	97	36	98
rect	36	97	37	98
rect	37	97	38	98
rect	38	97	39	98
rect	39	97	40	98
rect	40	97	41	98
rect	41	97	42	98
rect	42	97	43	98
rect	43	97	44	98
rect	44	97	45	98
rect	45	97	46	98
rect	46	97	47	98
rect	47	97	48	98
rect	49	97	50	98
rect	50	97	51	98
rect	51	97	52	98
rect	52	97	53	98
rect	53	97	54	98
rect	54	97	55	98
rect	55	97	56	98
rect	56	97	57	98
rect	57	97	58	98
rect	58	97	59	98
rect	59	97	60	98
rect	60	97	61	98
rect	61	97	62	98
rect	62	97	63	98
rect	63	97	64	98
rect	64	97	65	98
rect	65	97	66	98
rect	66	97	67	98
rect	67	97	68	98
rect	68	97	69	98
rect	69	97	70	98
rect	70	97	71	98
rect	71	97	72	98
rect	72	97	73	98
rect	73	97	74	98
rect	74	97	75	98
rect	75	97	76	98
rect	76	97	77	98
rect	77	97	78	98
rect	78	97	79	98
rect	79	97	80	98
rect	80	97	81	98
rect	81	97	82	98
rect	82	97	83	98
rect	83	97	84	98
rect	84	97	85	98
rect	85	97	86	98
rect	86	97	87	98
rect	87	97	88	98
rect	88	97	89	98
rect	89	97	90	98
rect	90	97	91	98
rect	91	97	92	98
rect	92	97	93	98
rect	93	97	94	98
rect	94	97	95	98
rect	95	97	96	98
rect	96	97	97	98
rect	98	97	99	98
rect	99	97	100	98
rect	100	97	101	98
rect	101	97	102	98
rect	102	97	103	98
rect	103	97	104	98
rect	105	97	106	98
rect	106	97	107	98
rect	107	97	108	98
rect	108	97	109	98
rect	109	97	110	98
rect	110	97	111	98
rect	111	97	112	98
rect	112	97	113	98
rect	113	97	114	98
rect	114	97	115	98
rect	115	97	116	98
rect	116	97	117	98
rect	117	97	118	98
rect	118	97	119	98
rect	119	97	120	98
rect	120	97	121	98
rect	121	97	122	98
rect	122	97	123	98
rect	123	97	124	98
rect	124	97	125	98
rect	125	97	126	98
rect	126	97	127	98
rect	127	97	128	98
rect	128	97	129	98
rect	129	97	130	98
rect	130	97	131	98
rect	131	97	132	98
rect	132	97	133	98
rect	133	97	134	98
rect	134	97	135	98
rect	135	97	136	98
rect	136	97	137	98
rect	137	97	138	98
rect	138	97	139	98
rect	139	97	140	98
rect	140	97	141	98
rect	141	97	142	98
rect	142	97	143	98
rect	143	97	144	98
rect	144	97	145	98
rect	145	97	146	98
rect	146	97	147	98
rect	147	97	148	98
rect	148	97	149	98
rect	149	97	150	98
rect	150	97	151	98
rect	151	97	152	98
rect	152	97	153	98
rect	153	97	154	98
rect	154	97	155	98
rect	155	97	156	98
rect	156	97	157	98
rect	157	97	158	98
rect	158	97	159	98
rect	160	97	161	98
rect	161	97	162	98
rect	162	97	163	98
rect	163	97	164	98
rect	164	97	165	98
rect	165	97	166	98
rect	166	97	167	98
rect	167	97	168	98
rect	168	97	169	98
rect	169	97	170	98
rect	170	97	171	98
rect	171	97	172	98
rect	172	97	173	98
rect	173	97	174	98
rect	174	97	175	98
rect	175	97	176	98
rect	176	97	177	98
rect	177	97	178	98
rect	178	97	179	98
rect	179	97	180	98
rect	180	97	181	98
rect	181	97	182	98
rect	182	97	183	98
rect	183	97	184	98
rect	184	97	185	98
rect	185	97	186	98
rect	186	97	187	98
rect	187	97	188	98
rect	188	97	189	98
rect	189	97	190	98
rect	190	97	191	98
rect	191	97	192	98
rect	192	97	193	98
rect	193	97	194	98
rect	194	97	195	98
rect	195	97	196	98
rect	196	97	197	98
rect	197	97	198	98
rect	198	97	199	98
rect	199	97	200	98
rect	200	97	201	98
rect	201	97	202	98
rect	202	97	203	98
rect	203	97	204	98
rect	204	97	205	98
rect	205	97	206	98
rect	206	97	207	98
rect	207	97	208	98
rect	208	97	209	98
rect	209	97	210	98
rect	210	97	211	98
rect	212	97	213	98
rect	213	97	214	98
rect	214	97	215	98
rect	215	97	216	98
rect	216	97	217	98
rect	217	97	218	98
rect	218	97	219	98
rect	219	97	220	98
rect	220	97	221	98
rect	221	97	222	98
rect	222	97	223	98
rect	223	97	224	98
rect	224	97	225	98
rect	225	97	226	98
rect	226	97	227	98
rect	227	97	228	98
rect	228	97	229	98
rect	229	97	230	98
rect	230	97	231	98
rect	231	97	232	98
rect	232	97	233	98
rect	233	97	234	98
rect	234	97	235	98
rect	235	97	236	98
rect	236	97	237	98
rect	237	97	238	98
rect	238	97	239	98
rect	239	97	240	98
rect	240	97	241	98
rect	241	97	242	98
rect	242	97	243	98
rect	243	97	244	98
rect	244	97	245	98
rect	245	97	246	98
rect	246	97	247	98
rect	247	97	248	98
rect	248	97	249	98
rect	249	97	250	98
rect	250	97	251	98
rect	251	97	252	98
rect	252	97	253	98
rect	253	97	254	98
rect	254	97	255	98
rect	255	97	256	98
rect	256	97	257	98
rect	257	97	258	98
rect	258	97	259	98
rect	259	97	260	98
rect	260	97	261	98
rect	261	97	262	98
rect	262	97	263	98
rect	263	97	264	98
rect	264	97	265	98
rect	265	97	266	98
rect	266	97	267	98
rect	267	97	268	98
rect	268	97	269	98
rect	269	97	270	98
rect	270	97	271	98
rect	271	97	272	98
rect	272	97	273	98
rect	273	97	274	98
rect	274	97	275	98
rect	275	97	276	98
rect	276	97	277	98
rect	277	97	278	98
rect	278	97	279	98
rect	279	97	280	98
rect	280	97	281	98
rect	281	97	282	98
rect	282	97	283	98
rect	283	97	284	98
rect	284	97	285	98
rect	285	97	286	98
rect	286	97	287	98
rect	287	97	288	98
rect	288	97	289	98
rect	289	97	290	98
rect	290	97	291	98
rect	291	97	292	98
rect	292	97	293	98
rect	293	97	294	98
rect	294	97	295	98
rect	295	97	296	98
rect	296	97	297	98
rect	297	97	298	98
rect	298	97	299	98
rect	299	97	300	98
rect	300	97	301	98
rect	301	97	302	98
rect	302	97	303	98
rect	303	97	304	98
rect	304	97	305	98
rect	305	97	306	98
rect	306	97	307	98
rect	307	97	308	98
rect	308	97	309	98
rect	309	97	310	98
rect	310	97	311	98
rect	311	97	312	98
rect	312	97	313	98
rect	313	97	314	98
rect	314	97	315	98
rect	315	97	316	98
rect	316	97	317	98
rect	317	97	318	98
rect	318	97	319	98
rect	319	97	320	98
rect	320	97	321	98
rect	321	97	322	98
rect	322	97	323	98
rect	323	97	324	98
rect	324	97	325	98
rect	325	97	326	98
rect	326	97	327	98
rect	327	97	328	98
rect	328	97	329	98
rect	329	97	330	98
rect	330	97	331	98
rect	331	97	332	98
rect	332	97	333	98
rect	333	97	334	98
rect	334	97	335	98
rect	335	97	336	98
rect	336	97	337	98
rect	337	97	338	98
rect	338	97	339	98
rect	339	97	340	98
rect	340	97	341	98
rect	341	97	342	98
rect	342	97	343	98
rect	343	97	344	98
rect	344	97	345	98
rect	345	97	346	98
rect	346	97	347	98
rect	347	97	348	98
rect	348	97	349	98
rect	349	97	350	98
rect	350	97	351	98
rect	351	97	352	98
rect	352	97	353	98
rect	353	97	354	98
rect	354	97	355	98
rect	355	97	356	98
rect	356	97	357	98
rect	357	97	358	98
rect	358	97	359	98
rect	359	97	360	98
rect	360	97	361	98
rect	361	97	362	98
rect	362	97	363	98
rect	363	97	364	98
rect	364	97	365	98
rect	365	97	366	98
rect	366	97	367	98
rect	367	97	368	98
rect	368	97	369	98
rect	369	97	370	98
rect	370	97	371	98
rect	371	97	372	98
rect	372	97	373	98
rect	373	97	374	98
rect	374	97	375	98
rect	375	97	376	98
rect	376	97	377	98
rect	377	97	378	98
rect	378	97	379	98
rect	379	97	380	98
rect	380	97	381	98
rect	381	97	382	98
rect	382	97	383	98
rect	383	97	384	98
rect	384	97	385	98
rect	385	97	386	98
rect	386	97	387	98
rect	387	97	388	98
rect	388	97	389	98
rect	389	97	390	98
rect	390	97	391	98
rect	391	97	392	98
rect	392	97	393	98
rect	393	97	394	98
rect	394	97	395	98
rect	395	97	396	98
rect	396	97	397	98
rect	397	97	398	98
rect	398	97	399	98
rect	399	97	400	98
rect	400	97	401	98
rect	401	97	402	98
rect	402	97	403	98
rect	403	97	404	98
rect	0	98	1	99
rect	1	98	2	99
rect	2	98	3	99
rect	3	98	4	99
rect	4	98	5	99
rect	5	98	6	99
rect	7	98	8	99
rect	8	98	9	99
rect	9	98	10	99
rect	10	98	11	99
rect	11	98	12	99
rect	12	98	13	99
rect	14	98	15	99
rect	15	98	16	99
rect	16	98	17	99
rect	17	98	18	99
rect	18	98	19	99
rect	19	98	20	99
rect	21	98	22	99
rect	22	98	23	99
rect	23	98	24	99
rect	24	98	25	99
rect	25	98	26	99
rect	26	98	27	99
rect	27	98	28	99
rect	28	98	29	99
rect	29	98	30	99
rect	30	98	31	99
rect	31	98	32	99
rect	32	98	33	99
rect	33	98	34	99
rect	34	98	35	99
rect	35	98	36	99
rect	36	98	37	99
rect	37	98	38	99
rect	38	98	39	99
rect	39	98	40	99
rect	40	98	41	99
rect	41	98	42	99
rect	42	98	43	99
rect	43	98	44	99
rect	44	98	45	99
rect	45	98	46	99
rect	46	98	47	99
rect	47	98	48	99
rect	49	98	50	99
rect	50	98	51	99
rect	51	98	52	99
rect	52	98	53	99
rect	53	98	54	99
rect	54	98	55	99
rect	55	98	56	99
rect	56	98	57	99
rect	57	98	58	99
rect	58	98	59	99
rect	59	98	60	99
rect	60	98	61	99
rect	61	98	62	99
rect	62	98	63	99
rect	63	98	64	99
rect	64	98	65	99
rect	65	98	66	99
rect	66	98	67	99
rect	67	98	68	99
rect	68	98	69	99
rect	69	98	70	99
rect	70	98	71	99
rect	71	98	72	99
rect	72	98	73	99
rect	73	98	74	99
rect	74	98	75	99
rect	75	98	76	99
rect	76	98	77	99
rect	77	98	78	99
rect	78	98	79	99
rect	79	98	80	99
rect	80	98	81	99
rect	81	98	82	99
rect	82	98	83	99
rect	83	98	84	99
rect	84	98	85	99
rect	85	98	86	99
rect	86	98	87	99
rect	87	98	88	99
rect	88	98	89	99
rect	89	98	90	99
rect	90	98	91	99
rect	91	98	92	99
rect	92	98	93	99
rect	93	98	94	99
rect	94	98	95	99
rect	95	98	96	99
rect	96	98	97	99
rect	98	98	99	99
rect	99	98	100	99
rect	100	98	101	99
rect	101	98	102	99
rect	102	98	103	99
rect	103	98	104	99
rect	105	98	106	99
rect	106	98	107	99
rect	107	98	108	99
rect	108	98	109	99
rect	109	98	110	99
rect	110	98	111	99
rect	111	98	112	99
rect	112	98	113	99
rect	113	98	114	99
rect	114	98	115	99
rect	115	98	116	99
rect	116	98	117	99
rect	117	98	118	99
rect	118	98	119	99
rect	119	98	120	99
rect	120	98	121	99
rect	121	98	122	99
rect	122	98	123	99
rect	123	98	124	99
rect	124	98	125	99
rect	125	98	126	99
rect	126	98	127	99
rect	127	98	128	99
rect	128	98	129	99
rect	129	98	130	99
rect	130	98	131	99
rect	131	98	132	99
rect	132	98	133	99
rect	133	98	134	99
rect	134	98	135	99
rect	135	98	136	99
rect	136	98	137	99
rect	137	98	138	99
rect	138	98	139	99
rect	139	98	140	99
rect	140	98	141	99
rect	141	98	142	99
rect	142	98	143	99
rect	143	98	144	99
rect	144	98	145	99
rect	145	98	146	99
rect	146	98	147	99
rect	147	98	148	99
rect	148	98	149	99
rect	149	98	150	99
rect	150	98	151	99
rect	151	98	152	99
rect	152	98	153	99
rect	153	98	154	99
rect	154	98	155	99
rect	155	98	156	99
rect	156	98	157	99
rect	157	98	158	99
rect	158	98	159	99
rect	160	98	161	99
rect	161	98	162	99
rect	162	98	163	99
rect	163	98	164	99
rect	164	98	165	99
rect	165	98	166	99
rect	166	98	167	99
rect	167	98	168	99
rect	168	98	169	99
rect	169	98	170	99
rect	170	98	171	99
rect	171	98	172	99
rect	172	98	173	99
rect	173	98	174	99
rect	174	98	175	99
rect	175	98	176	99
rect	176	98	177	99
rect	177	98	178	99
rect	178	98	179	99
rect	179	98	180	99
rect	180	98	181	99
rect	181	98	182	99
rect	182	98	183	99
rect	183	98	184	99
rect	184	98	185	99
rect	185	98	186	99
rect	186	98	187	99
rect	187	98	188	99
rect	188	98	189	99
rect	189	98	190	99
rect	190	98	191	99
rect	191	98	192	99
rect	192	98	193	99
rect	193	98	194	99
rect	194	98	195	99
rect	195	98	196	99
rect	196	98	197	99
rect	197	98	198	99
rect	198	98	199	99
rect	199	98	200	99
rect	200	98	201	99
rect	201	98	202	99
rect	202	98	203	99
rect	203	98	204	99
rect	204	98	205	99
rect	205	98	206	99
rect	206	98	207	99
rect	207	98	208	99
rect	208	98	209	99
rect	209	98	210	99
rect	210	98	211	99
rect	212	98	213	99
rect	213	98	214	99
rect	214	98	215	99
rect	215	98	216	99
rect	216	98	217	99
rect	217	98	218	99
rect	218	98	219	99
rect	219	98	220	99
rect	220	98	221	99
rect	221	98	222	99
rect	222	98	223	99
rect	223	98	224	99
rect	224	98	225	99
rect	225	98	226	99
rect	226	98	227	99
rect	227	98	228	99
rect	228	98	229	99
rect	229	98	230	99
rect	230	98	231	99
rect	231	98	232	99
rect	232	98	233	99
rect	233	98	234	99
rect	234	98	235	99
rect	235	98	236	99
rect	236	98	237	99
rect	237	98	238	99
rect	238	98	239	99
rect	239	98	240	99
rect	240	98	241	99
rect	241	98	242	99
rect	242	98	243	99
rect	243	98	244	99
rect	244	98	245	99
rect	245	98	246	99
rect	246	98	247	99
rect	247	98	248	99
rect	248	98	249	99
rect	249	98	250	99
rect	250	98	251	99
rect	251	98	252	99
rect	252	98	253	99
rect	253	98	254	99
rect	254	98	255	99
rect	255	98	256	99
rect	256	98	257	99
rect	257	98	258	99
rect	258	98	259	99
rect	259	98	260	99
rect	260	98	261	99
rect	261	98	262	99
rect	262	98	263	99
rect	263	98	264	99
rect	264	98	265	99
rect	265	98	266	99
rect	266	98	267	99
rect	267	98	268	99
rect	268	98	269	99
rect	269	98	270	99
rect	270	98	271	99
rect	271	98	272	99
rect	272	98	273	99
rect	273	98	274	99
rect	274	98	275	99
rect	275	98	276	99
rect	276	98	277	99
rect	277	98	278	99
rect	278	98	279	99
rect	279	98	280	99
rect	280	98	281	99
rect	281	98	282	99
rect	282	98	283	99
rect	283	98	284	99
rect	284	98	285	99
rect	285	98	286	99
rect	286	98	287	99
rect	287	98	288	99
rect	288	98	289	99
rect	289	98	290	99
rect	290	98	291	99
rect	291	98	292	99
rect	292	98	293	99
rect	293	98	294	99
rect	294	98	295	99
rect	295	98	296	99
rect	296	98	297	99
rect	297	98	298	99
rect	298	98	299	99
rect	299	98	300	99
rect	300	98	301	99
rect	301	98	302	99
rect	302	98	303	99
rect	303	98	304	99
rect	304	98	305	99
rect	305	98	306	99
rect	306	98	307	99
rect	307	98	308	99
rect	308	98	309	99
rect	309	98	310	99
rect	310	98	311	99
rect	311	98	312	99
rect	312	98	313	99
rect	313	98	314	99
rect	314	98	315	99
rect	315	98	316	99
rect	316	98	317	99
rect	317	98	318	99
rect	318	98	319	99
rect	319	98	320	99
rect	320	98	321	99
rect	321	98	322	99
rect	322	98	323	99
rect	323	98	324	99
rect	324	98	325	99
rect	325	98	326	99
rect	326	98	327	99
rect	327	98	328	99
rect	328	98	329	99
rect	329	98	330	99
rect	330	98	331	99
rect	331	98	332	99
rect	332	98	333	99
rect	333	98	334	99
rect	334	98	335	99
rect	335	98	336	99
rect	336	98	337	99
rect	337	98	338	99
rect	338	98	339	99
rect	339	98	340	99
rect	340	98	341	99
rect	341	98	342	99
rect	342	98	343	99
rect	343	98	344	99
rect	344	98	345	99
rect	345	98	346	99
rect	346	98	347	99
rect	347	98	348	99
rect	348	98	349	99
rect	349	98	350	99
rect	350	98	351	99
rect	351	98	352	99
rect	352	98	353	99
rect	353	98	354	99
rect	354	98	355	99
rect	355	98	356	99
rect	356	98	357	99
rect	357	98	358	99
rect	358	98	359	99
rect	359	98	360	99
rect	360	98	361	99
rect	361	98	362	99
rect	362	98	363	99
rect	363	98	364	99
rect	364	98	365	99
rect	365	98	366	99
rect	366	98	367	99
rect	367	98	368	99
rect	368	98	369	99
rect	369	98	370	99
rect	370	98	371	99
rect	371	98	372	99
rect	372	98	373	99
rect	373	98	374	99
rect	374	98	375	99
rect	375	98	376	99
rect	376	98	377	99
rect	377	98	378	99
rect	378	98	379	99
rect	379	98	380	99
rect	380	98	381	99
rect	381	98	382	99
rect	382	98	383	99
rect	383	98	384	99
rect	384	98	385	99
rect	385	98	386	99
rect	386	98	387	99
rect	387	98	388	99
rect	388	98	389	99
rect	389	98	390	99
rect	390	98	391	99
rect	391	98	392	99
rect	392	98	393	99
rect	393	98	394	99
rect	394	98	395	99
rect	395	98	396	99
rect	396	98	397	99
rect	397	98	398	99
rect	398	98	399	99
rect	399	98	400	99
rect	400	98	401	99
rect	401	98	402	99
rect	402	98	403	99
rect	403	98	404	99
rect	0	99	1	100
rect	1	99	2	100
rect	2	99	3	100
rect	3	99	4	100
rect	4	99	5	100
rect	5	99	6	100
rect	7	99	8	100
rect	8	99	9	100
rect	9	99	10	100
rect	10	99	11	100
rect	11	99	12	100
rect	12	99	13	100
rect	14	99	15	100
rect	15	99	16	100
rect	16	99	17	100
rect	17	99	18	100
rect	18	99	19	100
rect	19	99	20	100
rect	21	99	22	100
rect	22	99	23	100
rect	23	99	24	100
rect	24	99	25	100
rect	25	99	26	100
rect	26	99	27	100
rect	27	99	28	100
rect	28	99	29	100
rect	29	99	30	100
rect	30	99	31	100
rect	31	99	32	100
rect	32	99	33	100
rect	33	99	34	100
rect	34	99	35	100
rect	35	99	36	100
rect	36	99	37	100
rect	37	99	38	100
rect	38	99	39	100
rect	39	99	40	100
rect	40	99	41	100
rect	41	99	42	100
rect	42	99	43	100
rect	43	99	44	100
rect	44	99	45	100
rect	45	99	46	100
rect	46	99	47	100
rect	47	99	48	100
rect	49	99	50	100
rect	50	99	51	100
rect	51	99	52	100
rect	52	99	53	100
rect	53	99	54	100
rect	54	99	55	100
rect	55	99	56	100
rect	56	99	57	100
rect	57	99	58	100
rect	58	99	59	100
rect	59	99	60	100
rect	60	99	61	100
rect	61	99	62	100
rect	62	99	63	100
rect	63	99	64	100
rect	64	99	65	100
rect	65	99	66	100
rect	66	99	67	100
rect	67	99	68	100
rect	68	99	69	100
rect	69	99	70	100
rect	70	99	71	100
rect	71	99	72	100
rect	72	99	73	100
rect	73	99	74	100
rect	74	99	75	100
rect	75	99	76	100
rect	76	99	77	100
rect	77	99	78	100
rect	78	99	79	100
rect	79	99	80	100
rect	80	99	81	100
rect	81	99	82	100
rect	82	99	83	100
rect	83	99	84	100
rect	84	99	85	100
rect	85	99	86	100
rect	86	99	87	100
rect	87	99	88	100
rect	88	99	89	100
rect	89	99	90	100
rect	90	99	91	100
rect	91	99	92	100
rect	92	99	93	100
rect	93	99	94	100
rect	94	99	95	100
rect	95	99	96	100
rect	96	99	97	100
rect	98	99	99	100
rect	99	99	100	100
rect	100	99	101	100
rect	101	99	102	100
rect	102	99	103	100
rect	103	99	104	100
rect	105	99	106	100
rect	106	99	107	100
rect	107	99	108	100
rect	108	99	109	100
rect	109	99	110	100
rect	110	99	111	100
rect	111	99	112	100
rect	112	99	113	100
rect	113	99	114	100
rect	114	99	115	100
rect	115	99	116	100
rect	116	99	117	100
rect	117	99	118	100
rect	118	99	119	100
rect	119	99	120	100
rect	120	99	121	100
rect	121	99	122	100
rect	122	99	123	100
rect	123	99	124	100
rect	124	99	125	100
rect	125	99	126	100
rect	126	99	127	100
rect	127	99	128	100
rect	128	99	129	100
rect	129	99	130	100
rect	130	99	131	100
rect	131	99	132	100
rect	132	99	133	100
rect	133	99	134	100
rect	134	99	135	100
rect	135	99	136	100
rect	136	99	137	100
rect	137	99	138	100
rect	138	99	139	100
rect	139	99	140	100
rect	140	99	141	100
rect	141	99	142	100
rect	142	99	143	100
rect	143	99	144	100
rect	144	99	145	100
rect	145	99	146	100
rect	146	99	147	100
rect	147	99	148	100
rect	148	99	149	100
rect	149	99	150	100
rect	150	99	151	100
rect	151	99	152	100
rect	152	99	153	100
rect	153	99	154	100
rect	154	99	155	100
rect	155	99	156	100
rect	156	99	157	100
rect	157	99	158	100
rect	158	99	159	100
rect	160	99	161	100
rect	161	99	162	100
rect	162	99	163	100
rect	163	99	164	100
rect	164	99	165	100
rect	165	99	166	100
rect	166	99	167	100
rect	167	99	168	100
rect	168	99	169	100
rect	169	99	170	100
rect	170	99	171	100
rect	171	99	172	100
rect	172	99	173	100
rect	173	99	174	100
rect	174	99	175	100
rect	175	99	176	100
rect	176	99	177	100
rect	177	99	178	100
rect	178	99	179	100
rect	179	99	180	100
rect	180	99	181	100
rect	181	99	182	100
rect	182	99	183	100
rect	183	99	184	100
rect	184	99	185	100
rect	185	99	186	100
rect	186	99	187	100
rect	187	99	188	100
rect	188	99	189	100
rect	189	99	190	100
rect	190	99	191	100
rect	191	99	192	100
rect	192	99	193	100
rect	193	99	194	100
rect	194	99	195	100
rect	195	99	196	100
rect	196	99	197	100
rect	197	99	198	100
rect	198	99	199	100
rect	199	99	200	100
rect	200	99	201	100
rect	201	99	202	100
rect	202	99	203	100
rect	203	99	204	100
rect	204	99	205	100
rect	205	99	206	100
rect	206	99	207	100
rect	207	99	208	100
rect	208	99	209	100
rect	209	99	210	100
rect	210	99	211	100
rect	212	99	213	100
rect	213	99	214	100
rect	214	99	215	100
rect	215	99	216	100
rect	216	99	217	100
rect	217	99	218	100
rect	218	99	219	100
rect	219	99	220	100
rect	220	99	221	100
rect	221	99	222	100
rect	222	99	223	100
rect	223	99	224	100
rect	224	99	225	100
rect	225	99	226	100
rect	226	99	227	100
rect	227	99	228	100
rect	228	99	229	100
rect	229	99	230	100
rect	230	99	231	100
rect	231	99	232	100
rect	232	99	233	100
rect	233	99	234	100
rect	234	99	235	100
rect	235	99	236	100
rect	236	99	237	100
rect	237	99	238	100
rect	238	99	239	100
rect	239	99	240	100
rect	240	99	241	100
rect	241	99	242	100
rect	242	99	243	100
rect	243	99	244	100
rect	244	99	245	100
rect	245	99	246	100
rect	246	99	247	100
rect	247	99	248	100
rect	248	99	249	100
rect	249	99	250	100
rect	250	99	251	100
rect	251	99	252	100
rect	252	99	253	100
rect	253	99	254	100
rect	254	99	255	100
rect	255	99	256	100
rect	256	99	257	100
rect	257	99	258	100
rect	258	99	259	100
rect	259	99	260	100
rect	260	99	261	100
rect	261	99	262	100
rect	262	99	263	100
rect	263	99	264	100
rect	264	99	265	100
rect	265	99	266	100
rect	266	99	267	100
rect	267	99	268	100
rect	268	99	269	100
rect	269	99	270	100
rect	270	99	271	100
rect	271	99	272	100
rect	272	99	273	100
rect	273	99	274	100
rect	274	99	275	100
rect	275	99	276	100
rect	276	99	277	100
rect	277	99	278	100
rect	278	99	279	100
rect	279	99	280	100
rect	280	99	281	100
rect	281	99	282	100
rect	282	99	283	100
rect	283	99	284	100
rect	284	99	285	100
rect	285	99	286	100
rect	286	99	287	100
rect	287	99	288	100
rect	288	99	289	100
rect	289	99	290	100
rect	290	99	291	100
rect	291	99	292	100
rect	292	99	293	100
rect	293	99	294	100
rect	294	99	295	100
rect	295	99	296	100
rect	296	99	297	100
rect	297	99	298	100
rect	298	99	299	100
rect	299	99	300	100
rect	300	99	301	100
rect	301	99	302	100
rect	302	99	303	100
rect	303	99	304	100
rect	304	99	305	100
rect	305	99	306	100
rect	306	99	307	100
rect	307	99	308	100
rect	308	99	309	100
rect	309	99	310	100
rect	310	99	311	100
rect	311	99	312	100
rect	312	99	313	100
rect	313	99	314	100
rect	314	99	315	100
rect	315	99	316	100
rect	316	99	317	100
rect	317	99	318	100
rect	318	99	319	100
rect	319	99	320	100
rect	320	99	321	100
rect	321	99	322	100
rect	322	99	323	100
rect	323	99	324	100
rect	324	99	325	100
rect	325	99	326	100
rect	326	99	327	100
rect	327	99	328	100
rect	328	99	329	100
rect	329	99	330	100
rect	330	99	331	100
rect	331	99	332	100
rect	332	99	333	100
rect	333	99	334	100
rect	334	99	335	100
rect	335	99	336	100
rect	336	99	337	100
rect	337	99	338	100
rect	338	99	339	100
rect	339	99	340	100
rect	340	99	341	100
rect	341	99	342	100
rect	342	99	343	100
rect	343	99	344	100
rect	344	99	345	100
rect	345	99	346	100
rect	346	99	347	100
rect	347	99	348	100
rect	348	99	349	100
rect	349	99	350	100
rect	350	99	351	100
rect	351	99	352	100
rect	352	99	353	100
rect	353	99	354	100
rect	354	99	355	100
rect	355	99	356	100
rect	356	99	357	100
rect	357	99	358	100
rect	358	99	359	100
rect	359	99	360	100
rect	360	99	361	100
rect	361	99	362	100
rect	362	99	363	100
rect	363	99	364	100
rect	364	99	365	100
rect	365	99	366	100
rect	366	99	367	100
rect	367	99	368	100
rect	368	99	369	100
rect	369	99	370	100
rect	370	99	371	100
rect	371	99	372	100
rect	372	99	373	100
rect	373	99	374	100
rect	374	99	375	100
rect	375	99	376	100
rect	376	99	377	100
rect	377	99	378	100
rect	378	99	379	100
rect	379	99	380	100
rect	380	99	381	100
rect	381	99	382	100
rect	382	99	383	100
rect	383	99	384	100
rect	384	99	385	100
rect	385	99	386	100
rect	386	99	387	100
rect	387	99	388	100
rect	388	99	389	100
rect	389	99	390	100
rect	390	99	391	100
rect	391	99	392	100
rect	392	99	393	100
rect	393	99	394	100
rect	394	99	395	100
rect	395	99	396	100
rect	396	99	397	100
rect	397	99	398	100
rect	398	99	399	100
rect	399	99	400	100
rect	400	99	401	100
rect	401	99	402	100
rect	402	99	403	100
rect	403	99	404	100
rect	0	100	1	101
rect	1	100	2	101
rect	2	100	3	101
rect	3	100	4	101
rect	4	100	5	101
rect	5	100	6	101
rect	7	100	8	101
rect	8	100	9	101
rect	9	100	10	101
rect	10	100	11	101
rect	11	100	12	101
rect	12	100	13	101
rect	14	100	15	101
rect	15	100	16	101
rect	16	100	17	101
rect	17	100	18	101
rect	18	100	19	101
rect	19	100	20	101
rect	21	100	22	101
rect	22	100	23	101
rect	23	100	24	101
rect	24	100	25	101
rect	25	100	26	101
rect	26	100	27	101
rect	27	100	28	101
rect	28	100	29	101
rect	29	100	30	101
rect	30	100	31	101
rect	31	100	32	101
rect	32	100	33	101
rect	33	100	34	101
rect	34	100	35	101
rect	35	100	36	101
rect	36	100	37	101
rect	37	100	38	101
rect	38	100	39	101
rect	39	100	40	101
rect	40	100	41	101
rect	41	100	42	101
rect	42	100	43	101
rect	43	100	44	101
rect	44	100	45	101
rect	45	100	46	101
rect	46	100	47	101
rect	47	100	48	101
rect	49	100	50	101
rect	50	100	51	101
rect	51	100	52	101
rect	52	100	53	101
rect	53	100	54	101
rect	54	100	55	101
rect	55	100	56	101
rect	56	100	57	101
rect	57	100	58	101
rect	58	100	59	101
rect	59	100	60	101
rect	60	100	61	101
rect	61	100	62	101
rect	62	100	63	101
rect	63	100	64	101
rect	64	100	65	101
rect	65	100	66	101
rect	66	100	67	101
rect	67	100	68	101
rect	68	100	69	101
rect	69	100	70	101
rect	70	100	71	101
rect	71	100	72	101
rect	72	100	73	101
rect	73	100	74	101
rect	74	100	75	101
rect	75	100	76	101
rect	76	100	77	101
rect	77	100	78	101
rect	78	100	79	101
rect	79	100	80	101
rect	80	100	81	101
rect	81	100	82	101
rect	82	100	83	101
rect	83	100	84	101
rect	84	100	85	101
rect	85	100	86	101
rect	86	100	87	101
rect	87	100	88	101
rect	88	100	89	101
rect	89	100	90	101
rect	90	100	91	101
rect	91	100	92	101
rect	92	100	93	101
rect	93	100	94	101
rect	94	100	95	101
rect	95	100	96	101
rect	96	100	97	101
rect	98	100	99	101
rect	99	100	100	101
rect	100	100	101	101
rect	101	100	102	101
rect	102	100	103	101
rect	103	100	104	101
rect	105	100	106	101
rect	106	100	107	101
rect	107	100	108	101
rect	108	100	109	101
rect	109	100	110	101
rect	110	100	111	101
rect	111	100	112	101
rect	112	100	113	101
rect	113	100	114	101
rect	114	100	115	101
rect	115	100	116	101
rect	116	100	117	101
rect	117	100	118	101
rect	118	100	119	101
rect	119	100	120	101
rect	120	100	121	101
rect	121	100	122	101
rect	122	100	123	101
rect	123	100	124	101
rect	124	100	125	101
rect	125	100	126	101
rect	126	100	127	101
rect	127	100	128	101
rect	128	100	129	101
rect	129	100	130	101
rect	130	100	131	101
rect	131	100	132	101
rect	132	100	133	101
rect	133	100	134	101
rect	134	100	135	101
rect	135	100	136	101
rect	136	100	137	101
rect	137	100	138	101
rect	138	100	139	101
rect	139	100	140	101
rect	140	100	141	101
rect	141	100	142	101
rect	142	100	143	101
rect	143	100	144	101
rect	144	100	145	101
rect	145	100	146	101
rect	146	100	147	101
rect	147	100	148	101
rect	148	100	149	101
rect	149	100	150	101
rect	150	100	151	101
rect	151	100	152	101
rect	152	100	153	101
rect	153	100	154	101
rect	154	100	155	101
rect	155	100	156	101
rect	156	100	157	101
rect	157	100	158	101
rect	158	100	159	101
rect	160	100	161	101
rect	161	100	162	101
rect	162	100	163	101
rect	163	100	164	101
rect	164	100	165	101
rect	165	100	166	101
rect	166	100	167	101
rect	167	100	168	101
rect	168	100	169	101
rect	169	100	170	101
rect	170	100	171	101
rect	171	100	172	101
rect	172	100	173	101
rect	173	100	174	101
rect	174	100	175	101
rect	175	100	176	101
rect	176	100	177	101
rect	177	100	178	101
rect	178	100	179	101
rect	179	100	180	101
rect	180	100	181	101
rect	181	100	182	101
rect	182	100	183	101
rect	183	100	184	101
rect	184	100	185	101
rect	185	100	186	101
rect	186	100	187	101
rect	187	100	188	101
rect	188	100	189	101
rect	189	100	190	101
rect	190	100	191	101
rect	191	100	192	101
rect	192	100	193	101
rect	193	100	194	101
rect	194	100	195	101
rect	195	100	196	101
rect	196	100	197	101
rect	197	100	198	101
rect	198	100	199	101
rect	199	100	200	101
rect	200	100	201	101
rect	201	100	202	101
rect	202	100	203	101
rect	203	100	204	101
rect	204	100	205	101
rect	205	100	206	101
rect	206	100	207	101
rect	207	100	208	101
rect	208	100	209	101
rect	209	100	210	101
rect	210	100	211	101
rect	212	100	213	101
rect	213	100	214	101
rect	214	100	215	101
rect	215	100	216	101
rect	216	100	217	101
rect	217	100	218	101
rect	218	100	219	101
rect	219	100	220	101
rect	220	100	221	101
rect	221	100	222	101
rect	222	100	223	101
rect	223	100	224	101
rect	224	100	225	101
rect	225	100	226	101
rect	226	100	227	101
rect	227	100	228	101
rect	228	100	229	101
rect	229	100	230	101
rect	230	100	231	101
rect	231	100	232	101
rect	232	100	233	101
rect	233	100	234	101
rect	234	100	235	101
rect	235	100	236	101
rect	236	100	237	101
rect	237	100	238	101
rect	238	100	239	101
rect	239	100	240	101
rect	240	100	241	101
rect	241	100	242	101
rect	242	100	243	101
rect	243	100	244	101
rect	244	100	245	101
rect	245	100	246	101
rect	246	100	247	101
rect	247	100	248	101
rect	248	100	249	101
rect	249	100	250	101
rect	250	100	251	101
rect	251	100	252	101
rect	252	100	253	101
rect	253	100	254	101
rect	254	100	255	101
rect	255	100	256	101
rect	256	100	257	101
rect	257	100	258	101
rect	258	100	259	101
rect	259	100	260	101
rect	260	100	261	101
rect	261	100	262	101
rect	262	100	263	101
rect	263	100	264	101
rect	264	100	265	101
rect	265	100	266	101
rect	266	100	267	101
rect	267	100	268	101
rect	268	100	269	101
rect	269	100	270	101
rect	270	100	271	101
rect	271	100	272	101
rect	272	100	273	101
rect	273	100	274	101
rect	274	100	275	101
rect	275	100	276	101
rect	276	100	277	101
rect	277	100	278	101
rect	278	100	279	101
rect	279	100	280	101
rect	280	100	281	101
rect	281	100	282	101
rect	282	100	283	101
rect	283	100	284	101
rect	284	100	285	101
rect	285	100	286	101
rect	286	100	287	101
rect	287	100	288	101
rect	288	100	289	101
rect	289	100	290	101
rect	290	100	291	101
rect	291	100	292	101
rect	292	100	293	101
rect	293	100	294	101
rect	294	100	295	101
rect	295	100	296	101
rect	296	100	297	101
rect	297	100	298	101
rect	298	100	299	101
rect	299	100	300	101
rect	300	100	301	101
rect	301	100	302	101
rect	302	100	303	101
rect	303	100	304	101
rect	304	100	305	101
rect	305	100	306	101
rect	306	100	307	101
rect	307	100	308	101
rect	308	100	309	101
rect	309	100	310	101
rect	310	100	311	101
rect	311	100	312	101
rect	312	100	313	101
rect	313	100	314	101
rect	314	100	315	101
rect	315	100	316	101
rect	316	100	317	101
rect	317	100	318	101
rect	318	100	319	101
rect	319	100	320	101
rect	320	100	321	101
rect	321	100	322	101
rect	322	100	323	101
rect	323	100	324	101
rect	324	100	325	101
rect	325	100	326	101
rect	326	100	327	101
rect	327	100	328	101
rect	328	100	329	101
rect	329	100	330	101
rect	330	100	331	101
rect	331	100	332	101
rect	332	100	333	101
rect	333	100	334	101
rect	334	100	335	101
rect	335	100	336	101
rect	336	100	337	101
rect	337	100	338	101
rect	338	100	339	101
rect	339	100	340	101
rect	340	100	341	101
rect	341	100	342	101
rect	342	100	343	101
rect	343	100	344	101
rect	344	100	345	101
rect	345	100	346	101
rect	346	100	347	101
rect	347	100	348	101
rect	348	100	349	101
rect	349	100	350	101
rect	350	100	351	101
rect	351	100	352	101
rect	352	100	353	101
rect	353	100	354	101
rect	354	100	355	101
rect	355	100	356	101
rect	356	100	357	101
rect	357	100	358	101
rect	358	100	359	101
rect	359	100	360	101
rect	360	100	361	101
rect	361	100	362	101
rect	362	100	363	101
rect	363	100	364	101
rect	364	100	365	101
rect	365	100	366	101
rect	366	100	367	101
rect	367	100	368	101
rect	368	100	369	101
rect	369	100	370	101
rect	370	100	371	101
rect	371	100	372	101
rect	372	100	373	101
rect	373	100	374	101
rect	374	100	375	101
rect	375	100	376	101
rect	376	100	377	101
rect	377	100	378	101
rect	378	100	379	101
rect	379	100	380	101
rect	380	100	381	101
rect	381	100	382	101
rect	382	100	383	101
rect	383	100	384	101
rect	384	100	385	101
rect	385	100	386	101
rect	386	100	387	101
rect	387	100	388	101
rect	388	100	389	101
rect	389	100	390	101
rect	390	100	391	101
rect	391	100	392	101
rect	392	100	393	101
rect	393	100	394	101
rect	394	100	395	101
rect	395	100	396	101
rect	396	100	397	101
rect	397	100	398	101
rect	398	100	399	101
rect	399	100	400	101
rect	400	100	401	101
rect	401	100	402	101
rect	402	100	403	101
rect	403	100	404	101
rect	0	101	1	102
rect	1	101	2	102
rect	2	101	3	102
rect	3	101	4	102
rect	4	101	5	102
rect	5	101	6	102
rect	7	101	8	102
rect	8	101	9	102
rect	9	101	10	102
rect	10	101	11	102
rect	11	101	12	102
rect	12	101	13	102
rect	14	101	15	102
rect	15	101	16	102
rect	16	101	17	102
rect	17	101	18	102
rect	18	101	19	102
rect	19	101	20	102
rect	21	101	22	102
rect	22	101	23	102
rect	23	101	24	102
rect	24	101	25	102
rect	25	101	26	102
rect	26	101	27	102
rect	27	101	28	102
rect	28	101	29	102
rect	29	101	30	102
rect	30	101	31	102
rect	31	101	32	102
rect	32	101	33	102
rect	33	101	34	102
rect	34	101	35	102
rect	35	101	36	102
rect	36	101	37	102
rect	37	101	38	102
rect	38	101	39	102
rect	39	101	40	102
rect	40	101	41	102
rect	41	101	42	102
rect	42	101	43	102
rect	43	101	44	102
rect	44	101	45	102
rect	45	101	46	102
rect	46	101	47	102
rect	47	101	48	102
rect	49	101	50	102
rect	50	101	51	102
rect	51	101	52	102
rect	52	101	53	102
rect	53	101	54	102
rect	54	101	55	102
rect	55	101	56	102
rect	56	101	57	102
rect	57	101	58	102
rect	58	101	59	102
rect	59	101	60	102
rect	60	101	61	102
rect	61	101	62	102
rect	62	101	63	102
rect	63	101	64	102
rect	64	101	65	102
rect	65	101	66	102
rect	66	101	67	102
rect	67	101	68	102
rect	68	101	69	102
rect	69	101	70	102
rect	70	101	71	102
rect	71	101	72	102
rect	72	101	73	102
rect	73	101	74	102
rect	74	101	75	102
rect	75	101	76	102
rect	76	101	77	102
rect	77	101	78	102
rect	78	101	79	102
rect	79	101	80	102
rect	80	101	81	102
rect	81	101	82	102
rect	82	101	83	102
rect	83	101	84	102
rect	84	101	85	102
rect	85	101	86	102
rect	86	101	87	102
rect	87	101	88	102
rect	88	101	89	102
rect	89	101	90	102
rect	90	101	91	102
rect	91	101	92	102
rect	92	101	93	102
rect	93	101	94	102
rect	94	101	95	102
rect	95	101	96	102
rect	96	101	97	102
rect	98	101	99	102
rect	99	101	100	102
rect	100	101	101	102
rect	101	101	102	102
rect	102	101	103	102
rect	103	101	104	102
rect	105	101	106	102
rect	106	101	107	102
rect	107	101	108	102
rect	108	101	109	102
rect	109	101	110	102
rect	110	101	111	102
rect	111	101	112	102
rect	112	101	113	102
rect	113	101	114	102
rect	114	101	115	102
rect	115	101	116	102
rect	116	101	117	102
rect	117	101	118	102
rect	118	101	119	102
rect	119	101	120	102
rect	120	101	121	102
rect	121	101	122	102
rect	122	101	123	102
rect	123	101	124	102
rect	124	101	125	102
rect	125	101	126	102
rect	126	101	127	102
rect	127	101	128	102
rect	128	101	129	102
rect	129	101	130	102
rect	130	101	131	102
rect	131	101	132	102
rect	132	101	133	102
rect	133	101	134	102
rect	134	101	135	102
rect	135	101	136	102
rect	136	101	137	102
rect	137	101	138	102
rect	138	101	139	102
rect	139	101	140	102
rect	140	101	141	102
rect	141	101	142	102
rect	142	101	143	102
rect	143	101	144	102
rect	144	101	145	102
rect	145	101	146	102
rect	146	101	147	102
rect	147	101	148	102
rect	148	101	149	102
rect	149	101	150	102
rect	150	101	151	102
rect	151	101	152	102
rect	152	101	153	102
rect	153	101	154	102
rect	154	101	155	102
rect	155	101	156	102
rect	156	101	157	102
rect	157	101	158	102
rect	158	101	159	102
rect	160	101	161	102
rect	161	101	162	102
rect	162	101	163	102
rect	163	101	164	102
rect	164	101	165	102
rect	165	101	166	102
rect	166	101	167	102
rect	167	101	168	102
rect	168	101	169	102
rect	169	101	170	102
rect	170	101	171	102
rect	171	101	172	102
rect	172	101	173	102
rect	173	101	174	102
rect	174	101	175	102
rect	175	101	176	102
rect	176	101	177	102
rect	177	101	178	102
rect	178	101	179	102
rect	179	101	180	102
rect	180	101	181	102
rect	181	101	182	102
rect	182	101	183	102
rect	183	101	184	102
rect	184	101	185	102
rect	185	101	186	102
rect	186	101	187	102
rect	187	101	188	102
rect	188	101	189	102
rect	189	101	190	102
rect	190	101	191	102
rect	191	101	192	102
rect	192	101	193	102
rect	193	101	194	102
rect	194	101	195	102
rect	195	101	196	102
rect	196	101	197	102
rect	197	101	198	102
rect	198	101	199	102
rect	199	101	200	102
rect	200	101	201	102
rect	201	101	202	102
rect	202	101	203	102
rect	203	101	204	102
rect	204	101	205	102
rect	205	101	206	102
rect	206	101	207	102
rect	207	101	208	102
rect	208	101	209	102
rect	209	101	210	102
rect	210	101	211	102
rect	212	101	213	102
rect	213	101	214	102
rect	214	101	215	102
rect	215	101	216	102
rect	216	101	217	102
rect	217	101	218	102
rect	218	101	219	102
rect	219	101	220	102
rect	220	101	221	102
rect	221	101	222	102
rect	222	101	223	102
rect	223	101	224	102
rect	224	101	225	102
rect	225	101	226	102
rect	226	101	227	102
rect	227	101	228	102
rect	228	101	229	102
rect	229	101	230	102
rect	230	101	231	102
rect	231	101	232	102
rect	232	101	233	102
rect	233	101	234	102
rect	234	101	235	102
rect	235	101	236	102
rect	236	101	237	102
rect	237	101	238	102
rect	238	101	239	102
rect	239	101	240	102
rect	240	101	241	102
rect	241	101	242	102
rect	242	101	243	102
rect	243	101	244	102
rect	244	101	245	102
rect	245	101	246	102
rect	246	101	247	102
rect	247	101	248	102
rect	248	101	249	102
rect	249	101	250	102
rect	250	101	251	102
rect	251	101	252	102
rect	252	101	253	102
rect	253	101	254	102
rect	254	101	255	102
rect	255	101	256	102
rect	256	101	257	102
rect	257	101	258	102
rect	258	101	259	102
rect	259	101	260	102
rect	260	101	261	102
rect	261	101	262	102
rect	262	101	263	102
rect	263	101	264	102
rect	264	101	265	102
rect	265	101	266	102
rect	266	101	267	102
rect	267	101	268	102
rect	268	101	269	102
rect	269	101	270	102
rect	270	101	271	102
rect	271	101	272	102
rect	272	101	273	102
rect	273	101	274	102
rect	274	101	275	102
rect	275	101	276	102
rect	276	101	277	102
rect	277	101	278	102
rect	278	101	279	102
rect	279	101	280	102
rect	280	101	281	102
rect	281	101	282	102
rect	282	101	283	102
rect	283	101	284	102
rect	284	101	285	102
rect	285	101	286	102
rect	286	101	287	102
rect	287	101	288	102
rect	288	101	289	102
rect	289	101	290	102
rect	290	101	291	102
rect	291	101	292	102
rect	292	101	293	102
rect	293	101	294	102
rect	294	101	295	102
rect	295	101	296	102
rect	296	101	297	102
rect	297	101	298	102
rect	298	101	299	102
rect	299	101	300	102
rect	300	101	301	102
rect	301	101	302	102
rect	302	101	303	102
rect	303	101	304	102
rect	304	101	305	102
rect	305	101	306	102
rect	306	101	307	102
rect	307	101	308	102
rect	308	101	309	102
rect	309	101	310	102
rect	310	101	311	102
rect	311	101	312	102
rect	312	101	313	102
rect	313	101	314	102
rect	314	101	315	102
rect	315	101	316	102
rect	316	101	317	102
rect	317	101	318	102
rect	318	101	319	102
rect	319	101	320	102
rect	320	101	321	102
rect	321	101	322	102
rect	322	101	323	102
rect	323	101	324	102
rect	324	101	325	102
rect	325	101	326	102
rect	326	101	327	102
rect	327	101	328	102
rect	328	101	329	102
rect	329	101	330	102
rect	330	101	331	102
rect	331	101	332	102
rect	332	101	333	102
rect	333	101	334	102
rect	334	101	335	102
rect	335	101	336	102
rect	336	101	337	102
rect	337	101	338	102
rect	338	101	339	102
rect	339	101	340	102
rect	340	101	341	102
rect	341	101	342	102
rect	342	101	343	102
rect	343	101	344	102
rect	344	101	345	102
rect	345	101	346	102
rect	346	101	347	102
rect	347	101	348	102
rect	348	101	349	102
rect	349	101	350	102
rect	350	101	351	102
rect	351	101	352	102
rect	352	101	353	102
rect	353	101	354	102
rect	354	101	355	102
rect	355	101	356	102
rect	356	101	357	102
rect	357	101	358	102
rect	358	101	359	102
rect	359	101	360	102
rect	360	101	361	102
rect	361	101	362	102
rect	362	101	363	102
rect	363	101	364	102
rect	364	101	365	102
rect	365	101	366	102
rect	366	101	367	102
rect	367	101	368	102
rect	368	101	369	102
rect	369	101	370	102
rect	370	101	371	102
rect	371	101	372	102
rect	372	101	373	102
rect	373	101	374	102
rect	374	101	375	102
rect	375	101	376	102
rect	376	101	377	102
rect	377	101	378	102
rect	378	101	379	102
rect	379	101	380	102
rect	380	101	381	102
rect	381	101	382	102
rect	382	101	383	102
rect	383	101	384	102
rect	384	101	385	102
rect	385	101	386	102
rect	386	101	387	102
rect	387	101	388	102
rect	388	101	389	102
rect	389	101	390	102
rect	390	101	391	102
rect	391	101	392	102
rect	392	101	393	102
rect	393	101	394	102
rect	394	101	395	102
rect	395	101	396	102
rect	396	101	397	102
rect	397	101	398	102
rect	398	101	399	102
rect	399	101	400	102
rect	400	101	401	102
rect	401	101	402	102
rect	402	101	403	102
rect	403	101	404	102
rect	0	102	1	103
rect	1	102	2	103
rect	2	102	3	103
rect	3	102	4	103
rect	4	102	5	103
rect	5	102	6	103
rect	7	102	8	103
rect	8	102	9	103
rect	9	102	10	103
rect	10	102	11	103
rect	11	102	12	103
rect	12	102	13	103
rect	14	102	15	103
rect	15	102	16	103
rect	16	102	17	103
rect	17	102	18	103
rect	18	102	19	103
rect	19	102	20	103
rect	21	102	22	103
rect	22	102	23	103
rect	23	102	24	103
rect	24	102	25	103
rect	25	102	26	103
rect	26	102	27	103
rect	27	102	28	103
rect	28	102	29	103
rect	29	102	30	103
rect	30	102	31	103
rect	31	102	32	103
rect	32	102	33	103
rect	33	102	34	103
rect	34	102	35	103
rect	35	102	36	103
rect	36	102	37	103
rect	37	102	38	103
rect	38	102	39	103
rect	39	102	40	103
rect	40	102	41	103
rect	41	102	42	103
rect	42	102	43	103
rect	43	102	44	103
rect	44	102	45	103
rect	45	102	46	103
rect	46	102	47	103
rect	47	102	48	103
rect	49	102	50	103
rect	50	102	51	103
rect	51	102	52	103
rect	52	102	53	103
rect	53	102	54	103
rect	54	102	55	103
rect	55	102	56	103
rect	56	102	57	103
rect	57	102	58	103
rect	58	102	59	103
rect	59	102	60	103
rect	60	102	61	103
rect	61	102	62	103
rect	62	102	63	103
rect	63	102	64	103
rect	64	102	65	103
rect	65	102	66	103
rect	66	102	67	103
rect	67	102	68	103
rect	68	102	69	103
rect	69	102	70	103
rect	70	102	71	103
rect	71	102	72	103
rect	72	102	73	103
rect	73	102	74	103
rect	74	102	75	103
rect	75	102	76	103
rect	76	102	77	103
rect	77	102	78	103
rect	78	102	79	103
rect	79	102	80	103
rect	80	102	81	103
rect	81	102	82	103
rect	82	102	83	103
rect	83	102	84	103
rect	84	102	85	103
rect	85	102	86	103
rect	86	102	87	103
rect	87	102	88	103
rect	88	102	89	103
rect	89	102	90	103
rect	90	102	91	103
rect	91	102	92	103
rect	92	102	93	103
rect	93	102	94	103
rect	94	102	95	103
rect	95	102	96	103
rect	96	102	97	103
rect	98	102	99	103
rect	99	102	100	103
rect	100	102	101	103
rect	101	102	102	103
rect	102	102	103	103
rect	103	102	104	103
rect	105	102	106	103
rect	106	102	107	103
rect	107	102	108	103
rect	108	102	109	103
rect	109	102	110	103
rect	110	102	111	103
rect	111	102	112	103
rect	112	102	113	103
rect	113	102	114	103
rect	114	102	115	103
rect	115	102	116	103
rect	116	102	117	103
rect	117	102	118	103
rect	118	102	119	103
rect	119	102	120	103
rect	120	102	121	103
rect	121	102	122	103
rect	122	102	123	103
rect	123	102	124	103
rect	124	102	125	103
rect	125	102	126	103
rect	126	102	127	103
rect	127	102	128	103
rect	128	102	129	103
rect	129	102	130	103
rect	130	102	131	103
rect	131	102	132	103
rect	132	102	133	103
rect	133	102	134	103
rect	134	102	135	103
rect	135	102	136	103
rect	136	102	137	103
rect	137	102	138	103
rect	138	102	139	103
rect	139	102	140	103
rect	140	102	141	103
rect	141	102	142	103
rect	142	102	143	103
rect	143	102	144	103
rect	144	102	145	103
rect	145	102	146	103
rect	146	102	147	103
rect	147	102	148	103
rect	148	102	149	103
rect	149	102	150	103
rect	150	102	151	103
rect	151	102	152	103
rect	152	102	153	103
rect	153	102	154	103
rect	154	102	155	103
rect	155	102	156	103
rect	156	102	157	103
rect	157	102	158	103
rect	158	102	159	103
rect	160	102	161	103
rect	161	102	162	103
rect	162	102	163	103
rect	163	102	164	103
rect	164	102	165	103
rect	165	102	166	103
rect	166	102	167	103
rect	167	102	168	103
rect	168	102	169	103
rect	169	102	170	103
rect	170	102	171	103
rect	171	102	172	103
rect	172	102	173	103
rect	173	102	174	103
rect	174	102	175	103
rect	175	102	176	103
rect	176	102	177	103
rect	177	102	178	103
rect	178	102	179	103
rect	179	102	180	103
rect	180	102	181	103
rect	181	102	182	103
rect	182	102	183	103
rect	183	102	184	103
rect	184	102	185	103
rect	185	102	186	103
rect	186	102	187	103
rect	187	102	188	103
rect	188	102	189	103
rect	189	102	190	103
rect	190	102	191	103
rect	191	102	192	103
rect	192	102	193	103
rect	193	102	194	103
rect	194	102	195	103
rect	195	102	196	103
rect	196	102	197	103
rect	197	102	198	103
rect	198	102	199	103
rect	199	102	200	103
rect	200	102	201	103
rect	201	102	202	103
rect	202	102	203	103
rect	203	102	204	103
rect	204	102	205	103
rect	205	102	206	103
rect	206	102	207	103
rect	207	102	208	103
rect	208	102	209	103
rect	209	102	210	103
rect	210	102	211	103
rect	212	102	213	103
rect	213	102	214	103
rect	214	102	215	103
rect	215	102	216	103
rect	216	102	217	103
rect	217	102	218	103
rect	218	102	219	103
rect	219	102	220	103
rect	220	102	221	103
rect	221	102	222	103
rect	222	102	223	103
rect	223	102	224	103
rect	224	102	225	103
rect	225	102	226	103
rect	226	102	227	103
rect	227	102	228	103
rect	228	102	229	103
rect	229	102	230	103
rect	230	102	231	103
rect	231	102	232	103
rect	232	102	233	103
rect	233	102	234	103
rect	234	102	235	103
rect	235	102	236	103
rect	236	102	237	103
rect	237	102	238	103
rect	238	102	239	103
rect	239	102	240	103
rect	240	102	241	103
rect	241	102	242	103
rect	242	102	243	103
rect	243	102	244	103
rect	244	102	245	103
rect	245	102	246	103
rect	246	102	247	103
rect	247	102	248	103
rect	248	102	249	103
rect	249	102	250	103
rect	250	102	251	103
rect	251	102	252	103
rect	252	102	253	103
rect	253	102	254	103
rect	254	102	255	103
rect	255	102	256	103
rect	256	102	257	103
rect	257	102	258	103
rect	258	102	259	103
rect	259	102	260	103
rect	260	102	261	103
rect	261	102	262	103
rect	262	102	263	103
rect	263	102	264	103
rect	264	102	265	103
rect	265	102	266	103
rect	266	102	267	103
rect	267	102	268	103
rect	268	102	269	103
rect	269	102	270	103
rect	270	102	271	103
rect	271	102	272	103
rect	272	102	273	103
rect	273	102	274	103
rect	274	102	275	103
rect	275	102	276	103
rect	276	102	277	103
rect	277	102	278	103
rect	278	102	279	103
rect	279	102	280	103
rect	280	102	281	103
rect	281	102	282	103
rect	282	102	283	103
rect	283	102	284	103
rect	284	102	285	103
rect	285	102	286	103
rect	286	102	287	103
rect	287	102	288	103
rect	288	102	289	103
rect	289	102	290	103
rect	290	102	291	103
rect	291	102	292	103
rect	292	102	293	103
rect	293	102	294	103
rect	294	102	295	103
rect	295	102	296	103
rect	296	102	297	103
rect	297	102	298	103
rect	298	102	299	103
rect	299	102	300	103
rect	300	102	301	103
rect	301	102	302	103
rect	302	102	303	103
rect	303	102	304	103
rect	304	102	305	103
rect	305	102	306	103
rect	306	102	307	103
rect	307	102	308	103
rect	308	102	309	103
rect	309	102	310	103
rect	310	102	311	103
rect	311	102	312	103
rect	312	102	313	103
rect	313	102	314	103
rect	314	102	315	103
rect	315	102	316	103
rect	316	102	317	103
rect	317	102	318	103
rect	318	102	319	103
rect	319	102	320	103
rect	320	102	321	103
rect	321	102	322	103
rect	322	102	323	103
rect	323	102	324	103
rect	324	102	325	103
rect	325	102	326	103
rect	326	102	327	103
rect	327	102	328	103
rect	328	102	329	103
rect	329	102	330	103
rect	330	102	331	103
rect	331	102	332	103
rect	332	102	333	103
rect	333	102	334	103
rect	334	102	335	103
rect	335	102	336	103
rect	336	102	337	103
rect	337	102	338	103
rect	338	102	339	103
rect	339	102	340	103
rect	340	102	341	103
rect	341	102	342	103
rect	342	102	343	103
rect	343	102	344	103
rect	344	102	345	103
rect	345	102	346	103
rect	346	102	347	103
rect	347	102	348	103
rect	348	102	349	103
rect	349	102	350	103
rect	350	102	351	103
rect	351	102	352	103
rect	352	102	353	103
rect	353	102	354	103
rect	354	102	355	103
rect	355	102	356	103
rect	356	102	357	103
rect	357	102	358	103
rect	358	102	359	103
rect	359	102	360	103
rect	360	102	361	103
rect	361	102	362	103
rect	362	102	363	103
rect	363	102	364	103
rect	364	102	365	103
rect	365	102	366	103
rect	366	102	367	103
rect	367	102	368	103
rect	368	102	369	103
rect	369	102	370	103
rect	370	102	371	103
rect	371	102	372	103
rect	372	102	373	103
rect	373	102	374	103
rect	374	102	375	103
rect	375	102	376	103
rect	376	102	377	103
rect	377	102	378	103
rect	378	102	379	103
rect	379	102	380	103
rect	380	102	381	103
rect	381	102	382	103
rect	382	102	383	103
rect	383	102	384	103
rect	384	102	385	103
rect	385	102	386	103
rect	386	102	387	103
rect	387	102	388	103
rect	388	102	389	103
rect	389	102	390	103
rect	390	102	391	103
rect	391	102	392	103
rect	392	102	393	103
rect	393	102	394	103
rect	394	102	395	103
rect	395	102	396	103
rect	396	102	397	103
rect	397	102	398	103
rect	398	102	399	103
rect	399	102	400	103
rect	400	102	401	103
rect	401	102	402	103
rect	402	102	403	103
rect	403	102	404	103
rect	0	128	1	129
rect	1	128	2	129
rect	2	128	3	129
rect	3	128	4	129
rect	4	128	5	129
rect	5	128	6	129
rect	7	128	8	129
rect	8	128	9	129
rect	9	128	10	129
rect	10	128	11	129
rect	11	128	12	129
rect	12	128	13	129
rect	14	128	15	129
rect	15	128	16	129
rect	16	128	17	129
rect	17	128	18	129
rect	18	128	19	129
rect	19	128	20	129
rect	20	128	21	129
rect	21	128	22	129
rect	22	128	23	129
rect	23	128	24	129
rect	24	128	25	129
rect	25	128	26	129
rect	26	128	27	129
rect	27	128	28	129
rect	28	128	29	129
rect	29	128	30	129
rect	30	128	31	129
rect	31	128	32	129
rect	32	128	33	129
rect	33	128	34	129
rect	34	128	35	129
rect	35	128	36	129
rect	36	128	37	129
rect	37	128	38	129
rect	38	128	39	129
rect	39	128	40	129
rect	40	128	41	129
rect	41	128	42	129
rect	42	128	43	129
rect	43	128	44	129
rect	44	128	45	129
rect	45	128	46	129
rect	46	128	47	129
rect	47	128	48	129
rect	48	128	49	129
rect	49	128	50	129
rect	51	128	52	129
rect	52	128	53	129
rect	53	128	54	129
rect	54	128	55	129
rect	55	128	56	129
rect	56	128	57	129
rect	57	128	58	129
rect	58	128	59	129
rect	59	128	60	129
rect	60	128	61	129
rect	61	128	62	129
rect	62	128	63	129
rect	63	128	64	129
rect	64	128	65	129
rect	65	128	66	129
rect	66	128	67	129
rect	67	128	68	129
rect	68	128	69	129
rect	69	128	70	129
rect	70	128	71	129
rect	71	128	72	129
rect	72	128	73	129
rect	73	128	74	129
rect	74	128	75	129
rect	75	128	76	129
rect	76	128	77	129
rect	77	128	78	129
rect	79	128	80	129
rect	80	128	81	129
rect	81	128	82	129
rect	82	128	83	129
rect	83	128	84	129
rect	84	128	85	129
rect	85	128	86	129
rect	86	128	87	129
rect	87	128	88	129
rect	88	128	89	129
rect	89	128	90	129
rect	90	128	91	129
rect	91	128	92	129
rect	92	128	93	129
rect	93	128	94	129
rect	94	128	95	129
rect	95	128	96	129
rect	96	128	97	129
rect	97	128	98	129
rect	98	128	99	129
rect	99	128	100	129
rect	101	128	102	129
rect	102	128	103	129
rect	103	128	104	129
rect	104	128	105	129
rect	105	128	106	129
rect	106	128	107	129
rect	108	128	109	129
rect	109	128	110	129
rect	110	128	111	129
rect	111	128	112	129
rect	112	128	113	129
rect	113	128	114	129
rect	114	128	115	129
rect	115	128	116	129
rect	116	128	117	129
rect	117	128	118	129
rect	118	128	119	129
rect	119	128	120	129
rect	120	128	121	129
rect	121	128	122	129
rect	122	128	123	129
rect	123	128	124	129
rect	124	128	125	129
rect	125	128	126	129
rect	126	128	127	129
rect	127	128	128	129
rect	128	128	129	129
rect	129	128	130	129
rect	130	128	131	129
rect	131	128	132	129
rect	132	128	133	129
rect	133	128	134	129
rect	134	128	135	129
rect	135	128	136	129
rect	136	128	137	129
rect	137	128	138	129
rect	138	128	139	129
rect	139	128	140	129
rect	140	128	141	129
rect	141	128	142	129
rect	142	128	143	129
rect	143	128	144	129
rect	145	128	146	129
rect	146	128	147	129
rect	147	128	148	129
rect	148	128	149	129
rect	149	128	150	129
rect	150	128	151	129
rect	151	128	152	129
rect	152	128	153	129
rect	153	128	154	129
rect	154	128	155	129
rect	155	128	156	129
rect	156	128	157	129
rect	157	128	158	129
rect	158	128	159	129
rect	159	128	160	129
rect	160	128	161	129
rect	161	128	162	129
rect	162	128	163	129
rect	163	128	164	129
rect	164	128	165	129
rect	165	128	166	129
rect	167	128	168	129
rect	168	128	169	129
rect	169	128	170	129
rect	170	128	171	129
rect	171	128	172	129
rect	172	128	173	129
rect	173	128	174	129
rect	174	128	175	129
rect	175	128	176	129
rect	176	128	177	129
rect	177	128	178	129
rect	178	128	179	129
rect	179	128	180	129
rect	180	128	181	129
rect	181	128	182	129
rect	182	128	183	129
rect	183	128	184	129
rect	184	128	185	129
rect	185	128	186	129
rect	186	128	187	129
rect	187	128	188	129
rect	188	128	189	129
rect	189	128	190	129
rect	190	128	191	129
rect	191	128	192	129
rect	192	128	193	129
rect	193	128	194	129
rect	194	128	195	129
rect	195	128	196	129
rect	196	128	197	129
rect	197	128	198	129
rect	198	128	199	129
rect	199	128	200	129
rect	200	128	201	129
rect	201	128	202	129
rect	202	128	203	129
rect	203	128	204	129
rect	204	128	205	129
rect	205	128	206	129
rect	206	128	207	129
rect	207	128	208	129
rect	208	128	209	129
rect	209	128	210	129
rect	210	128	211	129
rect	211	128	212	129
rect	212	128	213	129
rect	213	128	214	129
rect	214	128	215	129
rect	215	128	216	129
rect	216	128	217	129
rect	217	128	218	129
rect	218	128	219	129
rect	219	128	220	129
rect	220	128	221	129
rect	221	128	222	129
rect	222	128	223	129
rect	223	128	224	129
rect	224	128	225	129
rect	225	128	226	129
rect	226	128	227	129
rect	227	128	228	129
rect	228	128	229	129
rect	229	128	230	129
rect	230	128	231	129
rect	231	128	232	129
rect	232	128	233	129
rect	233	128	234	129
rect	234	128	235	129
rect	235	128	236	129
rect	236	128	237	129
rect	237	128	238	129
rect	238	128	239	129
rect	239	128	240	129
rect	240	128	241	129
rect	241	128	242	129
rect	242	128	243	129
rect	243	128	244	129
rect	244	128	245	129
rect	245	128	246	129
rect	246	128	247	129
rect	247	128	248	129
rect	248	128	249	129
rect	249	128	250	129
rect	250	128	251	129
rect	251	128	252	129
rect	252	128	253	129
rect	253	128	254	129
rect	254	128	255	129
rect	255	128	256	129
rect	256	128	257	129
rect	257	128	258	129
rect	258	128	259	129
rect	259	128	260	129
rect	260	128	261	129
rect	261	128	262	129
rect	262	128	263	129
rect	263	128	264	129
rect	264	128	265	129
rect	265	128	266	129
rect	266	128	267	129
rect	267	128	268	129
rect	268	128	269	129
rect	269	128	270	129
rect	270	128	271	129
rect	271	128	272	129
rect	272	128	273	129
rect	273	128	274	129
rect	274	128	275	129
rect	275	128	276	129
rect	276	128	277	129
rect	277	128	278	129
rect	278	128	279	129
rect	279	128	280	129
rect	280	128	281	129
rect	281	128	282	129
rect	282	128	283	129
rect	283	128	284	129
rect	284	128	285	129
rect	285	128	286	129
rect	286	128	287	129
rect	287	128	288	129
rect	288	128	289	129
rect	289	128	290	129
rect	290	128	291	129
rect	291	128	292	129
rect	292	128	293	129
rect	293	128	294	129
rect	294	128	295	129
rect	295	128	296	129
rect	296	128	297	129
rect	297	128	298	129
rect	298	128	299	129
rect	299	128	300	129
rect	300	128	301	129
rect	301	128	302	129
rect	302	128	303	129
rect	303	128	304	129
rect	304	128	305	129
rect	305	128	306	129
rect	306	128	307	129
rect	307	128	308	129
rect	308	128	309	129
rect	309	128	310	129
rect	310	128	311	129
rect	311	128	312	129
rect	312	128	313	129
rect	313	128	314	129
rect	314	128	315	129
rect	315	128	316	129
rect	316	128	317	129
rect	317	128	318	129
rect	318	128	319	129
rect	319	128	320	129
rect	320	128	321	129
rect	321	128	322	129
rect	322	128	323	129
rect	323	128	324	129
rect	324	128	325	129
rect	325	128	326	129
rect	326	128	327	129
rect	327	128	328	129
rect	328	128	329	129
rect	329	128	330	129
rect	330	128	331	129
rect	331	128	332	129
rect	332	128	333	129
rect	333	128	334	129
rect	334	128	335	129
rect	335	128	336	129
rect	336	128	337	129
rect	337	128	338	129
rect	338	128	339	129
rect	339	128	340	129
rect	340	128	341	129
rect	341	128	342	129
rect	342	128	343	129
rect	343	128	344	129
rect	344	128	345	129
rect	345	128	346	129
rect	346	128	347	129
rect	347	128	348	129
rect	348	128	349	129
rect	349	128	350	129
rect	350	128	351	129
rect	351	128	352	129
rect	352	128	353	129
rect	353	128	354	129
rect	354	128	355	129
rect	355	128	356	129
rect	356	128	357	129
rect	357	128	358	129
rect	358	128	359	129
rect	359	128	360	129
rect	360	128	361	129
rect	361	128	362	129
rect	362	128	363	129
rect	363	128	364	129
rect	364	128	365	129
rect	365	128	366	129
rect	366	128	367	129
rect	367	128	368	129
rect	368	128	369	129
rect	369	128	370	129
rect	370	128	371	129
rect	371	128	372	129
rect	372	128	373	129
rect	373	128	374	129
rect	374	128	375	129
rect	375	128	376	129
rect	376	128	377	129
rect	377	128	378	129
rect	378	128	379	129
rect	379	128	380	129
rect	380	128	381	129
rect	381	128	382	129
rect	382	128	383	129
rect	383	128	384	129
rect	384	128	385	129
rect	385	128	386	129
rect	386	128	387	129
rect	387	128	388	129
rect	388	128	389	129
rect	389	128	390	129
rect	390	128	391	129
rect	391	128	392	129
rect	392	128	393	129
rect	393	128	394	129
rect	394	128	395	129
rect	395	128	396	129
rect	396	128	397	129
rect	397	128	398	129
rect	398	128	399	129
rect	399	128	400	129
rect	400	128	401	129
rect	401	128	402	129
rect	402	128	403	129
rect	403	128	404	129
rect	405	128	406	129
rect	406	128	407	129
rect	407	128	408	129
rect	408	128	409	129
rect	409	128	410	129
rect	410	128	411	129
rect	412	128	413	129
rect	413	128	414	129
rect	414	128	415	129
rect	415	128	416	129
rect	416	128	417	129
rect	417	128	418	129
rect	418	128	419	129
rect	419	128	420	129
rect	420	128	421	129
rect	0	129	1	130
rect	1	129	2	130
rect	2	129	3	130
rect	3	129	4	130
rect	4	129	5	130
rect	5	129	6	130
rect	7	129	8	130
rect	8	129	9	130
rect	9	129	10	130
rect	10	129	11	130
rect	11	129	12	130
rect	12	129	13	130
rect	14	129	15	130
rect	15	129	16	130
rect	16	129	17	130
rect	17	129	18	130
rect	18	129	19	130
rect	19	129	20	130
rect	20	129	21	130
rect	21	129	22	130
rect	22	129	23	130
rect	23	129	24	130
rect	24	129	25	130
rect	25	129	26	130
rect	26	129	27	130
rect	27	129	28	130
rect	28	129	29	130
rect	29	129	30	130
rect	30	129	31	130
rect	31	129	32	130
rect	32	129	33	130
rect	33	129	34	130
rect	34	129	35	130
rect	35	129	36	130
rect	36	129	37	130
rect	37	129	38	130
rect	38	129	39	130
rect	39	129	40	130
rect	40	129	41	130
rect	41	129	42	130
rect	42	129	43	130
rect	43	129	44	130
rect	44	129	45	130
rect	45	129	46	130
rect	46	129	47	130
rect	47	129	48	130
rect	48	129	49	130
rect	49	129	50	130
rect	51	129	52	130
rect	52	129	53	130
rect	53	129	54	130
rect	54	129	55	130
rect	55	129	56	130
rect	56	129	57	130
rect	57	129	58	130
rect	58	129	59	130
rect	59	129	60	130
rect	60	129	61	130
rect	61	129	62	130
rect	62	129	63	130
rect	63	129	64	130
rect	64	129	65	130
rect	65	129	66	130
rect	66	129	67	130
rect	67	129	68	130
rect	68	129	69	130
rect	69	129	70	130
rect	70	129	71	130
rect	71	129	72	130
rect	72	129	73	130
rect	73	129	74	130
rect	74	129	75	130
rect	75	129	76	130
rect	76	129	77	130
rect	77	129	78	130
rect	79	129	80	130
rect	80	129	81	130
rect	81	129	82	130
rect	82	129	83	130
rect	83	129	84	130
rect	84	129	85	130
rect	85	129	86	130
rect	86	129	87	130
rect	87	129	88	130
rect	88	129	89	130
rect	89	129	90	130
rect	90	129	91	130
rect	91	129	92	130
rect	92	129	93	130
rect	93	129	94	130
rect	94	129	95	130
rect	95	129	96	130
rect	96	129	97	130
rect	97	129	98	130
rect	98	129	99	130
rect	99	129	100	130
rect	101	129	102	130
rect	102	129	103	130
rect	103	129	104	130
rect	104	129	105	130
rect	105	129	106	130
rect	106	129	107	130
rect	108	129	109	130
rect	109	129	110	130
rect	110	129	111	130
rect	111	129	112	130
rect	112	129	113	130
rect	113	129	114	130
rect	114	129	115	130
rect	115	129	116	130
rect	116	129	117	130
rect	117	129	118	130
rect	118	129	119	130
rect	119	129	120	130
rect	120	129	121	130
rect	121	129	122	130
rect	122	129	123	130
rect	123	129	124	130
rect	124	129	125	130
rect	125	129	126	130
rect	126	129	127	130
rect	127	129	128	130
rect	128	129	129	130
rect	129	129	130	130
rect	130	129	131	130
rect	131	129	132	130
rect	132	129	133	130
rect	133	129	134	130
rect	134	129	135	130
rect	135	129	136	130
rect	136	129	137	130
rect	137	129	138	130
rect	138	129	139	130
rect	139	129	140	130
rect	140	129	141	130
rect	141	129	142	130
rect	142	129	143	130
rect	143	129	144	130
rect	145	129	146	130
rect	146	129	147	130
rect	147	129	148	130
rect	148	129	149	130
rect	149	129	150	130
rect	150	129	151	130
rect	151	129	152	130
rect	152	129	153	130
rect	153	129	154	130
rect	154	129	155	130
rect	155	129	156	130
rect	156	129	157	130
rect	157	129	158	130
rect	158	129	159	130
rect	159	129	160	130
rect	160	129	161	130
rect	161	129	162	130
rect	162	129	163	130
rect	163	129	164	130
rect	164	129	165	130
rect	165	129	166	130
rect	167	129	168	130
rect	168	129	169	130
rect	169	129	170	130
rect	170	129	171	130
rect	171	129	172	130
rect	172	129	173	130
rect	173	129	174	130
rect	174	129	175	130
rect	175	129	176	130
rect	176	129	177	130
rect	177	129	178	130
rect	178	129	179	130
rect	179	129	180	130
rect	180	129	181	130
rect	181	129	182	130
rect	182	129	183	130
rect	183	129	184	130
rect	184	129	185	130
rect	185	129	186	130
rect	186	129	187	130
rect	187	129	188	130
rect	188	129	189	130
rect	189	129	190	130
rect	190	129	191	130
rect	191	129	192	130
rect	192	129	193	130
rect	193	129	194	130
rect	194	129	195	130
rect	195	129	196	130
rect	196	129	197	130
rect	197	129	198	130
rect	198	129	199	130
rect	199	129	200	130
rect	200	129	201	130
rect	201	129	202	130
rect	202	129	203	130
rect	203	129	204	130
rect	204	129	205	130
rect	205	129	206	130
rect	206	129	207	130
rect	207	129	208	130
rect	208	129	209	130
rect	209	129	210	130
rect	210	129	211	130
rect	211	129	212	130
rect	212	129	213	130
rect	213	129	214	130
rect	214	129	215	130
rect	215	129	216	130
rect	216	129	217	130
rect	217	129	218	130
rect	218	129	219	130
rect	219	129	220	130
rect	220	129	221	130
rect	221	129	222	130
rect	222	129	223	130
rect	223	129	224	130
rect	224	129	225	130
rect	225	129	226	130
rect	226	129	227	130
rect	227	129	228	130
rect	228	129	229	130
rect	229	129	230	130
rect	230	129	231	130
rect	231	129	232	130
rect	232	129	233	130
rect	233	129	234	130
rect	234	129	235	130
rect	235	129	236	130
rect	236	129	237	130
rect	237	129	238	130
rect	238	129	239	130
rect	239	129	240	130
rect	240	129	241	130
rect	241	129	242	130
rect	242	129	243	130
rect	243	129	244	130
rect	244	129	245	130
rect	245	129	246	130
rect	246	129	247	130
rect	247	129	248	130
rect	248	129	249	130
rect	249	129	250	130
rect	250	129	251	130
rect	251	129	252	130
rect	252	129	253	130
rect	253	129	254	130
rect	254	129	255	130
rect	255	129	256	130
rect	256	129	257	130
rect	257	129	258	130
rect	258	129	259	130
rect	259	129	260	130
rect	260	129	261	130
rect	261	129	262	130
rect	262	129	263	130
rect	263	129	264	130
rect	264	129	265	130
rect	265	129	266	130
rect	266	129	267	130
rect	267	129	268	130
rect	268	129	269	130
rect	269	129	270	130
rect	270	129	271	130
rect	271	129	272	130
rect	272	129	273	130
rect	273	129	274	130
rect	274	129	275	130
rect	275	129	276	130
rect	276	129	277	130
rect	277	129	278	130
rect	278	129	279	130
rect	279	129	280	130
rect	280	129	281	130
rect	281	129	282	130
rect	282	129	283	130
rect	283	129	284	130
rect	284	129	285	130
rect	285	129	286	130
rect	286	129	287	130
rect	287	129	288	130
rect	288	129	289	130
rect	289	129	290	130
rect	290	129	291	130
rect	291	129	292	130
rect	292	129	293	130
rect	293	129	294	130
rect	294	129	295	130
rect	295	129	296	130
rect	296	129	297	130
rect	297	129	298	130
rect	298	129	299	130
rect	299	129	300	130
rect	300	129	301	130
rect	301	129	302	130
rect	302	129	303	130
rect	303	129	304	130
rect	304	129	305	130
rect	305	129	306	130
rect	306	129	307	130
rect	307	129	308	130
rect	308	129	309	130
rect	309	129	310	130
rect	310	129	311	130
rect	311	129	312	130
rect	312	129	313	130
rect	313	129	314	130
rect	314	129	315	130
rect	315	129	316	130
rect	316	129	317	130
rect	317	129	318	130
rect	318	129	319	130
rect	319	129	320	130
rect	320	129	321	130
rect	321	129	322	130
rect	322	129	323	130
rect	323	129	324	130
rect	324	129	325	130
rect	325	129	326	130
rect	326	129	327	130
rect	327	129	328	130
rect	328	129	329	130
rect	329	129	330	130
rect	330	129	331	130
rect	331	129	332	130
rect	332	129	333	130
rect	333	129	334	130
rect	334	129	335	130
rect	335	129	336	130
rect	336	129	337	130
rect	337	129	338	130
rect	338	129	339	130
rect	339	129	340	130
rect	340	129	341	130
rect	341	129	342	130
rect	342	129	343	130
rect	343	129	344	130
rect	344	129	345	130
rect	345	129	346	130
rect	346	129	347	130
rect	347	129	348	130
rect	348	129	349	130
rect	349	129	350	130
rect	350	129	351	130
rect	351	129	352	130
rect	352	129	353	130
rect	353	129	354	130
rect	354	129	355	130
rect	355	129	356	130
rect	356	129	357	130
rect	357	129	358	130
rect	358	129	359	130
rect	359	129	360	130
rect	360	129	361	130
rect	361	129	362	130
rect	362	129	363	130
rect	363	129	364	130
rect	364	129	365	130
rect	365	129	366	130
rect	366	129	367	130
rect	367	129	368	130
rect	368	129	369	130
rect	369	129	370	130
rect	370	129	371	130
rect	371	129	372	130
rect	372	129	373	130
rect	373	129	374	130
rect	374	129	375	130
rect	375	129	376	130
rect	376	129	377	130
rect	377	129	378	130
rect	378	129	379	130
rect	379	129	380	130
rect	380	129	381	130
rect	381	129	382	130
rect	382	129	383	130
rect	383	129	384	130
rect	384	129	385	130
rect	385	129	386	130
rect	386	129	387	130
rect	387	129	388	130
rect	388	129	389	130
rect	389	129	390	130
rect	390	129	391	130
rect	391	129	392	130
rect	392	129	393	130
rect	393	129	394	130
rect	394	129	395	130
rect	395	129	396	130
rect	396	129	397	130
rect	397	129	398	130
rect	398	129	399	130
rect	399	129	400	130
rect	400	129	401	130
rect	401	129	402	130
rect	402	129	403	130
rect	403	129	404	130
rect	405	129	406	130
rect	406	129	407	130
rect	407	129	408	130
rect	408	129	409	130
rect	409	129	410	130
rect	410	129	411	130
rect	412	129	413	130
rect	413	129	414	130
rect	414	129	415	130
rect	415	129	416	130
rect	416	129	417	130
rect	417	129	418	130
rect	418	129	419	130
rect	419	129	420	130
rect	420	129	421	130
rect	0	130	1	131
rect	1	130	2	131
rect	2	130	3	131
rect	3	130	4	131
rect	4	130	5	131
rect	5	130	6	131
rect	7	130	8	131
rect	8	130	9	131
rect	9	130	10	131
rect	10	130	11	131
rect	11	130	12	131
rect	12	130	13	131
rect	14	130	15	131
rect	15	130	16	131
rect	16	130	17	131
rect	17	130	18	131
rect	18	130	19	131
rect	19	130	20	131
rect	20	130	21	131
rect	21	130	22	131
rect	22	130	23	131
rect	23	130	24	131
rect	24	130	25	131
rect	25	130	26	131
rect	26	130	27	131
rect	27	130	28	131
rect	28	130	29	131
rect	29	130	30	131
rect	30	130	31	131
rect	31	130	32	131
rect	32	130	33	131
rect	33	130	34	131
rect	34	130	35	131
rect	35	130	36	131
rect	36	130	37	131
rect	37	130	38	131
rect	38	130	39	131
rect	39	130	40	131
rect	40	130	41	131
rect	41	130	42	131
rect	42	130	43	131
rect	43	130	44	131
rect	44	130	45	131
rect	45	130	46	131
rect	46	130	47	131
rect	47	130	48	131
rect	48	130	49	131
rect	49	130	50	131
rect	51	130	52	131
rect	52	130	53	131
rect	53	130	54	131
rect	54	130	55	131
rect	55	130	56	131
rect	56	130	57	131
rect	57	130	58	131
rect	58	130	59	131
rect	59	130	60	131
rect	60	130	61	131
rect	61	130	62	131
rect	62	130	63	131
rect	63	130	64	131
rect	64	130	65	131
rect	65	130	66	131
rect	66	130	67	131
rect	67	130	68	131
rect	68	130	69	131
rect	69	130	70	131
rect	70	130	71	131
rect	71	130	72	131
rect	72	130	73	131
rect	73	130	74	131
rect	74	130	75	131
rect	75	130	76	131
rect	76	130	77	131
rect	77	130	78	131
rect	79	130	80	131
rect	80	130	81	131
rect	81	130	82	131
rect	82	130	83	131
rect	83	130	84	131
rect	84	130	85	131
rect	85	130	86	131
rect	86	130	87	131
rect	87	130	88	131
rect	88	130	89	131
rect	89	130	90	131
rect	90	130	91	131
rect	91	130	92	131
rect	92	130	93	131
rect	93	130	94	131
rect	94	130	95	131
rect	95	130	96	131
rect	96	130	97	131
rect	97	130	98	131
rect	98	130	99	131
rect	99	130	100	131
rect	101	130	102	131
rect	102	130	103	131
rect	103	130	104	131
rect	104	130	105	131
rect	105	130	106	131
rect	106	130	107	131
rect	108	130	109	131
rect	109	130	110	131
rect	110	130	111	131
rect	111	130	112	131
rect	112	130	113	131
rect	113	130	114	131
rect	114	130	115	131
rect	115	130	116	131
rect	116	130	117	131
rect	117	130	118	131
rect	118	130	119	131
rect	119	130	120	131
rect	120	130	121	131
rect	121	130	122	131
rect	122	130	123	131
rect	123	130	124	131
rect	124	130	125	131
rect	125	130	126	131
rect	126	130	127	131
rect	127	130	128	131
rect	128	130	129	131
rect	129	130	130	131
rect	130	130	131	131
rect	131	130	132	131
rect	132	130	133	131
rect	133	130	134	131
rect	134	130	135	131
rect	135	130	136	131
rect	136	130	137	131
rect	137	130	138	131
rect	138	130	139	131
rect	139	130	140	131
rect	140	130	141	131
rect	141	130	142	131
rect	142	130	143	131
rect	143	130	144	131
rect	145	130	146	131
rect	146	130	147	131
rect	147	130	148	131
rect	148	130	149	131
rect	149	130	150	131
rect	150	130	151	131
rect	151	130	152	131
rect	152	130	153	131
rect	153	130	154	131
rect	154	130	155	131
rect	155	130	156	131
rect	156	130	157	131
rect	157	130	158	131
rect	158	130	159	131
rect	159	130	160	131
rect	160	130	161	131
rect	161	130	162	131
rect	162	130	163	131
rect	163	130	164	131
rect	164	130	165	131
rect	165	130	166	131
rect	167	130	168	131
rect	168	130	169	131
rect	169	130	170	131
rect	170	130	171	131
rect	171	130	172	131
rect	172	130	173	131
rect	173	130	174	131
rect	174	130	175	131
rect	175	130	176	131
rect	176	130	177	131
rect	177	130	178	131
rect	178	130	179	131
rect	179	130	180	131
rect	180	130	181	131
rect	181	130	182	131
rect	182	130	183	131
rect	183	130	184	131
rect	184	130	185	131
rect	185	130	186	131
rect	186	130	187	131
rect	187	130	188	131
rect	188	130	189	131
rect	189	130	190	131
rect	190	130	191	131
rect	191	130	192	131
rect	192	130	193	131
rect	193	130	194	131
rect	194	130	195	131
rect	195	130	196	131
rect	196	130	197	131
rect	197	130	198	131
rect	198	130	199	131
rect	199	130	200	131
rect	200	130	201	131
rect	201	130	202	131
rect	202	130	203	131
rect	203	130	204	131
rect	204	130	205	131
rect	205	130	206	131
rect	206	130	207	131
rect	207	130	208	131
rect	208	130	209	131
rect	209	130	210	131
rect	210	130	211	131
rect	211	130	212	131
rect	212	130	213	131
rect	213	130	214	131
rect	214	130	215	131
rect	215	130	216	131
rect	216	130	217	131
rect	217	130	218	131
rect	218	130	219	131
rect	219	130	220	131
rect	220	130	221	131
rect	221	130	222	131
rect	222	130	223	131
rect	223	130	224	131
rect	224	130	225	131
rect	225	130	226	131
rect	226	130	227	131
rect	227	130	228	131
rect	228	130	229	131
rect	229	130	230	131
rect	230	130	231	131
rect	231	130	232	131
rect	232	130	233	131
rect	233	130	234	131
rect	234	130	235	131
rect	235	130	236	131
rect	236	130	237	131
rect	237	130	238	131
rect	238	130	239	131
rect	239	130	240	131
rect	240	130	241	131
rect	241	130	242	131
rect	242	130	243	131
rect	243	130	244	131
rect	244	130	245	131
rect	245	130	246	131
rect	246	130	247	131
rect	247	130	248	131
rect	248	130	249	131
rect	249	130	250	131
rect	250	130	251	131
rect	251	130	252	131
rect	252	130	253	131
rect	253	130	254	131
rect	254	130	255	131
rect	255	130	256	131
rect	256	130	257	131
rect	257	130	258	131
rect	258	130	259	131
rect	259	130	260	131
rect	260	130	261	131
rect	261	130	262	131
rect	262	130	263	131
rect	263	130	264	131
rect	264	130	265	131
rect	265	130	266	131
rect	266	130	267	131
rect	267	130	268	131
rect	268	130	269	131
rect	269	130	270	131
rect	270	130	271	131
rect	271	130	272	131
rect	272	130	273	131
rect	273	130	274	131
rect	274	130	275	131
rect	275	130	276	131
rect	276	130	277	131
rect	277	130	278	131
rect	278	130	279	131
rect	279	130	280	131
rect	280	130	281	131
rect	281	130	282	131
rect	282	130	283	131
rect	283	130	284	131
rect	284	130	285	131
rect	285	130	286	131
rect	286	130	287	131
rect	287	130	288	131
rect	288	130	289	131
rect	289	130	290	131
rect	290	130	291	131
rect	291	130	292	131
rect	292	130	293	131
rect	293	130	294	131
rect	294	130	295	131
rect	295	130	296	131
rect	296	130	297	131
rect	297	130	298	131
rect	298	130	299	131
rect	299	130	300	131
rect	300	130	301	131
rect	301	130	302	131
rect	302	130	303	131
rect	303	130	304	131
rect	304	130	305	131
rect	305	130	306	131
rect	306	130	307	131
rect	307	130	308	131
rect	308	130	309	131
rect	309	130	310	131
rect	310	130	311	131
rect	311	130	312	131
rect	312	130	313	131
rect	313	130	314	131
rect	314	130	315	131
rect	315	130	316	131
rect	316	130	317	131
rect	317	130	318	131
rect	318	130	319	131
rect	319	130	320	131
rect	320	130	321	131
rect	321	130	322	131
rect	322	130	323	131
rect	323	130	324	131
rect	324	130	325	131
rect	325	130	326	131
rect	326	130	327	131
rect	327	130	328	131
rect	328	130	329	131
rect	329	130	330	131
rect	330	130	331	131
rect	331	130	332	131
rect	332	130	333	131
rect	333	130	334	131
rect	334	130	335	131
rect	335	130	336	131
rect	336	130	337	131
rect	337	130	338	131
rect	338	130	339	131
rect	339	130	340	131
rect	340	130	341	131
rect	341	130	342	131
rect	342	130	343	131
rect	343	130	344	131
rect	344	130	345	131
rect	345	130	346	131
rect	346	130	347	131
rect	347	130	348	131
rect	348	130	349	131
rect	349	130	350	131
rect	350	130	351	131
rect	351	130	352	131
rect	352	130	353	131
rect	353	130	354	131
rect	354	130	355	131
rect	355	130	356	131
rect	356	130	357	131
rect	357	130	358	131
rect	358	130	359	131
rect	359	130	360	131
rect	360	130	361	131
rect	361	130	362	131
rect	362	130	363	131
rect	363	130	364	131
rect	364	130	365	131
rect	365	130	366	131
rect	366	130	367	131
rect	367	130	368	131
rect	368	130	369	131
rect	369	130	370	131
rect	370	130	371	131
rect	371	130	372	131
rect	372	130	373	131
rect	373	130	374	131
rect	374	130	375	131
rect	375	130	376	131
rect	376	130	377	131
rect	377	130	378	131
rect	378	130	379	131
rect	379	130	380	131
rect	380	130	381	131
rect	381	130	382	131
rect	382	130	383	131
rect	383	130	384	131
rect	384	130	385	131
rect	385	130	386	131
rect	386	130	387	131
rect	387	130	388	131
rect	388	130	389	131
rect	389	130	390	131
rect	390	130	391	131
rect	391	130	392	131
rect	392	130	393	131
rect	393	130	394	131
rect	394	130	395	131
rect	395	130	396	131
rect	396	130	397	131
rect	397	130	398	131
rect	398	130	399	131
rect	399	130	400	131
rect	400	130	401	131
rect	401	130	402	131
rect	402	130	403	131
rect	403	130	404	131
rect	405	130	406	131
rect	406	130	407	131
rect	407	130	408	131
rect	408	130	409	131
rect	409	130	410	131
rect	410	130	411	131
rect	412	130	413	131
rect	413	130	414	131
rect	414	130	415	131
rect	415	130	416	131
rect	416	130	417	131
rect	417	130	418	131
rect	418	130	419	131
rect	419	130	420	131
rect	420	130	421	131
rect	0	131	1	132
rect	1	131	2	132
rect	2	131	3	132
rect	3	131	4	132
rect	4	131	5	132
rect	5	131	6	132
rect	7	131	8	132
rect	8	131	9	132
rect	9	131	10	132
rect	10	131	11	132
rect	11	131	12	132
rect	12	131	13	132
rect	14	131	15	132
rect	15	131	16	132
rect	16	131	17	132
rect	17	131	18	132
rect	18	131	19	132
rect	19	131	20	132
rect	20	131	21	132
rect	21	131	22	132
rect	22	131	23	132
rect	23	131	24	132
rect	24	131	25	132
rect	25	131	26	132
rect	26	131	27	132
rect	27	131	28	132
rect	28	131	29	132
rect	29	131	30	132
rect	30	131	31	132
rect	31	131	32	132
rect	32	131	33	132
rect	33	131	34	132
rect	34	131	35	132
rect	35	131	36	132
rect	36	131	37	132
rect	37	131	38	132
rect	38	131	39	132
rect	39	131	40	132
rect	40	131	41	132
rect	41	131	42	132
rect	42	131	43	132
rect	43	131	44	132
rect	44	131	45	132
rect	45	131	46	132
rect	46	131	47	132
rect	47	131	48	132
rect	48	131	49	132
rect	49	131	50	132
rect	51	131	52	132
rect	52	131	53	132
rect	53	131	54	132
rect	54	131	55	132
rect	55	131	56	132
rect	56	131	57	132
rect	57	131	58	132
rect	58	131	59	132
rect	59	131	60	132
rect	60	131	61	132
rect	61	131	62	132
rect	62	131	63	132
rect	63	131	64	132
rect	64	131	65	132
rect	65	131	66	132
rect	66	131	67	132
rect	67	131	68	132
rect	68	131	69	132
rect	69	131	70	132
rect	70	131	71	132
rect	71	131	72	132
rect	72	131	73	132
rect	73	131	74	132
rect	74	131	75	132
rect	75	131	76	132
rect	76	131	77	132
rect	77	131	78	132
rect	79	131	80	132
rect	80	131	81	132
rect	81	131	82	132
rect	82	131	83	132
rect	83	131	84	132
rect	84	131	85	132
rect	85	131	86	132
rect	86	131	87	132
rect	87	131	88	132
rect	88	131	89	132
rect	89	131	90	132
rect	90	131	91	132
rect	91	131	92	132
rect	92	131	93	132
rect	93	131	94	132
rect	94	131	95	132
rect	95	131	96	132
rect	96	131	97	132
rect	97	131	98	132
rect	98	131	99	132
rect	99	131	100	132
rect	101	131	102	132
rect	102	131	103	132
rect	103	131	104	132
rect	104	131	105	132
rect	105	131	106	132
rect	106	131	107	132
rect	108	131	109	132
rect	109	131	110	132
rect	110	131	111	132
rect	111	131	112	132
rect	112	131	113	132
rect	113	131	114	132
rect	114	131	115	132
rect	115	131	116	132
rect	116	131	117	132
rect	117	131	118	132
rect	118	131	119	132
rect	119	131	120	132
rect	120	131	121	132
rect	121	131	122	132
rect	122	131	123	132
rect	123	131	124	132
rect	124	131	125	132
rect	125	131	126	132
rect	126	131	127	132
rect	127	131	128	132
rect	128	131	129	132
rect	129	131	130	132
rect	130	131	131	132
rect	131	131	132	132
rect	132	131	133	132
rect	133	131	134	132
rect	134	131	135	132
rect	135	131	136	132
rect	136	131	137	132
rect	137	131	138	132
rect	138	131	139	132
rect	139	131	140	132
rect	140	131	141	132
rect	141	131	142	132
rect	142	131	143	132
rect	143	131	144	132
rect	145	131	146	132
rect	146	131	147	132
rect	147	131	148	132
rect	148	131	149	132
rect	149	131	150	132
rect	150	131	151	132
rect	151	131	152	132
rect	152	131	153	132
rect	153	131	154	132
rect	154	131	155	132
rect	155	131	156	132
rect	156	131	157	132
rect	157	131	158	132
rect	158	131	159	132
rect	159	131	160	132
rect	160	131	161	132
rect	161	131	162	132
rect	162	131	163	132
rect	163	131	164	132
rect	164	131	165	132
rect	165	131	166	132
rect	167	131	168	132
rect	168	131	169	132
rect	169	131	170	132
rect	170	131	171	132
rect	171	131	172	132
rect	172	131	173	132
rect	173	131	174	132
rect	174	131	175	132
rect	175	131	176	132
rect	176	131	177	132
rect	177	131	178	132
rect	178	131	179	132
rect	179	131	180	132
rect	180	131	181	132
rect	181	131	182	132
rect	182	131	183	132
rect	183	131	184	132
rect	184	131	185	132
rect	185	131	186	132
rect	186	131	187	132
rect	187	131	188	132
rect	188	131	189	132
rect	189	131	190	132
rect	190	131	191	132
rect	191	131	192	132
rect	192	131	193	132
rect	193	131	194	132
rect	194	131	195	132
rect	195	131	196	132
rect	196	131	197	132
rect	197	131	198	132
rect	198	131	199	132
rect	199	131	200	132
rect	200	131	201	132
rect	201	131	202	132
rect	202	131	203	132
rect	203	131	204	132
rect	204	131	205	132
rect	205	131	206	132
rect	206	131	207	132
rect	207	131	208	132
rect	208	131	209	132
rect	209	131	210	132
rect	210	131	211	132
rect	211	131	212	132
rect	212	131	213	132
rect	213	131	214	132
rect	214	131	215	132
rect	215	131	216	132
rect	216	131	217	132
rect	217	131	218	132
rect	218	131	219	132
rect	219	131	220	132
rect	220	131	221	132
rect	221	131	222	132
rect	222	131	223	132
rect	223	131	224	132
rect	224	131	225	132
rect	225	131	226	132
rect	226	131	227	132
rect	227	131	228	132
rect	228	131	229	132
rect	229	131	230	132
rect	230	131	231	132
rect	231	131	232	132
rect	232	131	233	132
rect	233	131	234	132
rect	234	131	235	132
rect	235	131	236	132
rect	236	131	237	132
rect	237	131	238	132
rect	238	131	239	132
rect	239	131	240	132
rect	240	131	241	132
rect	241	131	242	132
rect	242	131	243	132
rect	243	131	244	132
rect	244	131	245	132
rect	245	131	246	132
rect	246	131	247	132
rect	247	131	248	132
rect	248	131	249	132
rect	249	131	250	132
rect	250	131	251	132
rect	251	131	252	132
rect	252	131	253	132
rect	253	131	254	132
rect	254	131	255	132
rect	255	131	256	132
rect	256	131	257	132
rect	257	131	258	132
rect	258	131	259	132
rect	259	131	260	132
rect	260	131	261	132
rect	261	131	262	132
rect	262	131	263	132
rect	263	131	264	132
rect	264	131	265	132
rect	265	131	266	132
rect	266	131	267	132
rect	267	131	268	132
rect	268	131	269	132
rect	269	131	270	132
rect	270	131	271	132
rect	271	131	272	132
rect	272	131	273	132
rect	273	131	274	132
rect	274	131	275	132
rect	275	131	276	132
rect	276	131	277	132
rect	277	131	278	132
rect	278	131	279	132
rect	279	131	280	132
rect	280	131	281	132
rect	281	131	282	132
rect	282	131	283	132
rect	283	131	284	132
rect	284	131	285	132
rect	285	131	286	132
rect	286	131	287	132
rect	287	131	288	132
rect	288	131	289	132
rect	289	131	290	132
rect	290	131	291	132
rect	291	131	292	132
rect	292	131	293	132
rect	293	131	294	132
rect	294	131	295	132
rect	295	131	296	132
rect	296	131	297	132
rect	297	131	298	132
rect	298	131	299	132
rect	299	131	300	132
rect	300	131	301	132
rect	301	131	302	132
rect	302	131	303	132
rect	303	131	304	132
rect	304	131	305	132
rect	305	131	306	132
rect	306	131	307	132
rect	307	131	308	132
rect	308	131	309	132
rect	309	131	310	132
rect	310	131	311	132
rect	311	131	312	132
rect	312	131	313	132
rect	313	131	314	132
rect	314	131	315	132
rect	315	131	316	132
rect	316	131	317	132
rect	317	131	318	132
rect	318	131	319	132
rect	319	131	320	132
rect	320	131	321	132
rect	321	131	322	132
rect	322	131	323	132
rect	323	131	324	132
rect	324	131	325	132
rect	325	131	326	132
rect	326	131	327	132
rect	327	131	328	132
rect	328	131	329	132
rect	329	131	330	132
rect	330	131	331	132
rect	331	131	332	132
rect	332	131	333	132
rect	333	131	334	132
rect	334	131	335	132
rect	335	131	336	132
rect	336	131	337	132
rect	337	131	338	132
rect	338	131	339	132
rect	339	131	340	132
rect	340	131	341	132
rect	341	131	342	132
rect	342	131	343	132
rect	343	131	344	132
rect	344	131	345	132
rect	345	131	346	132
rect	346	131	347	132
rect	347	131	348	132
rect	348	131	349	132
rect	349	131	350	132
rect	350	131	351	132
rect	351	131	352	132
rect	352	131	353	132
rect	353	131	354	132
rect	354	131	355	132
rect	355	131	356	132
rect	356	131	357	132
rect	357	131	358	132
rect	358	131	359	132
rect	359	131	360	132
rect	360	131	361	132
rect	361	131	362	132
rect	362	131	363	132
rect	363	131	364	132
rect	364	131	365	132
rect	365	131	366	132
rect	366	131	367	132
rect	367	131	368	132
rect	368	131	369	132
rect	369	131	370	132
rect	370	131	371	132
rect	371	131	372	132
rect	372	131	373	132
rect	373	131	374	132
rect	374	131	375	132
rect	375	131	376	132
rect	376	131	377	132
rect	377	131	378	132
rect	378	131	379	132
rect	379	131	380	132
rect	380	131	381	132
rect	381	131	382	132
rect	382	131	383	132
rect	383	131	384	132
rect	384	131	385	132
rect	385	131	386	132
rect	386	131	387	132
rect	387	131	388	132
rect	388	131	389	132
rect	389	131	390	132
rect	390	131	391	132
rect	391	131	392	132
rect	392	131	393	132
rect	393	131	394	132
rect	394	131	395	132
rect	395	131	396	132
rect	396	131	397	132
rect	397	131	398	132
rect	398	131	399	132
rect	399	131	400	132
rect	400	131	401	132
rect	401	131	402	132
rect	402	131	403	132
rect	403	131	404	132
rect	405	131	406	132
rect	406	131	407	132
rect	407	131	408	132
rect	408	131	409	132
rect	409	131	410	132
rect	410	131	411	132
rect	412	131	413	132
rect	413	131	414	132
rect	414	131	415	132
rect	415	131	416	132
rect	416	131	417	132
rect	417	131	418	132
rect	418	131	419	132
rect	419	131	420	132
rect	420	131	421	132
rect	0	132	1	133
rect	1	132	2	133
rect	2	132	3	133
rect	3	132	4	133
rect	4	132	5	133
rect	5	132	6	133
rect	7	132	8	133
rect	8	132	9	133
rect	9	132	10	133
rect	10	132	11	133
rect	11	132	12	133
rect	12	132	13	133
rect	14	132	15	133
rect	15	132	16	133
rect	16	132	17	133
rect	17	132	18	133
rect	18	132	19	133
rect	19	132	20	133
rect	20	132	21	133
rect	21	132	22	133
rect	22	132	23	133
rect	23	132	24	133
rect	24	132	25	133
rect	25	132	26	133
rect	26	132	27	133
rect	27	132	28	133
rect	28	132	29	133
rect	29	132	30	133
rect	30	132	31	133
rect	31	132	32	133
rect	32	132	33	133
rect	33	132	34	133
rect	34	132	35	133
rect	35	132	36	133
rect	36	132	37	133
rect	37	132	38	133
rect	38	132	39	133
rect	39	132	40	133
rect	40	132	41	133
rect	41	132	42	133
rect	42	132	43	133
rect	43	132	44	133
rect	44	132	45	133
rect	45	132	46	133
rect	46	132	47	133
rect	47	132	48	133
rect	48	132	49	133
rect	49	132	50	133
rect	51	132	52	133
rect	52	132	53	133
rect	53	132	54	133
rect	54	132	55	133
rect	55	132	56	133
rect	56	132	57	133
rect	57	132	58	133
rect	58	132	59	133
rect	59	132	60	133
rect	60	132	61	133
rect	61	132	62	133
rect	62	132	63	133
rect	63	132	64	133
rect	64	132	65	133
rect	65	132	66	133
rect	66	132	67	133
rect	67	132	68	133
rect	68	132	69	133
rect	69	132	70	133
rect	70	132	71	133
rect	71	132	72	133
rect	72	132	73	133
rect	73	132	74	133
rect	74	132	75	133
rect	75	132	76	133
rect	76	132	77	133
rect	77	132	78	133
rect	79	132	80	133
rect	80	132	81	133
rect	81	132	82	133
rect	82	132	83	133
rect	83	132	84	133
rect	84	132	85	133
rect	85	132	86	133
rect	86	132	87	133
rect	87	132	88	133
rect	88	132	89	133
rect	89	132	90	133
rect	90	132	91	133
rect	91	132	92	133
rect	92	132	93	133
rect	93	132	94	133
rect	94	132	95	133
rect	95	132	96	133
rect	96	132	97	133
rect	97	132	98	133
rect	98	132	99	133
rect	99	132	100	133
rect	101	132	102	133
rect	102	132	103	133
rect	103	132	104	133
rect	104	132	105	133
rect	105	132	106	133
rect	106	132	107	133
rect	108	132	109	133
rect	109	132	110	133
rect	110	132	111	133
rect	111	132	112	133
rect	112	132	113	133
rect	113	132	114	133
rect	114	132	115	133
rect	115	132	116	133
rect	116	132	117	133
rect	117	132	118	133
rect	118	132	119	133
rect	119	132	120	133
rect	120	132	121	133
rect	121	132	122	133
rect	122	132	123	133
rect	123	132	124	133
rect	124	132	125	133
rect	125	132	126	133
rect	126	132	127	133
rect	127	132	128	133
rect	128	132	129	133
rect	129	132	130	133
rect	130	132	131	133
rect	131	132	132	133
rect	132	132	133	133
rect	133	132	134	133
rect	134	132	135	133
rect	135	132	136	133
rect	136	132	137	133
rect	137	132	138	133
rect	138	132	139	133
rect	139	132	140	133
rect	140	132	141	133
rect	141	132	142	133
rect	142	132	143	133
rect	143	132	144	133
rect	145	132	146	133
rect	146	132	147	133
rect	147	132	148	133
rect	148	132	149	133
rect	149	132	150	133
rect	150	132	151	133
rect	151	132	152	133
rect	152	132	153	133
rect	153	132	154	133
rect	154	132	155	133
rect	155	132	156	133
rect	156	132	157	133
rect	157	132	158	133
rect	158	132	159	133
rect	159	132	160	133
rect	160	132	161	133
rect	161	132	162	133
rect	162	132	163	133
rect	163	132	164	133
rect	164	132	165	133
rect	165	132	166	133
rect	167	132	168	133
rect	168	132	169	133
rect	169	132	170	133
rect	170	132	171	133
rect	171	132	172	133
rect	172	132	173	133
rect	173	132	174	133
rect	174	132	175	133
rect	175	132	176	133
rect	176	132	177	133
rect	177	132	178	133
rect	178	132	179	133
rect	179	132	180	133
rect	180	132	181	133
rect	181	132	182	133
rect	182	132	183	133
rect	183	132	184	133
rect	184	132	185	133
rect	185	132	186	133
rect	186	132	187	133
rect	187	132	188	133
rect	188	132	189	133
rect	189	132	190	133
rect	190	132	191	133
rect	191	132	192	133
rect	192	132	193	133
rect	193	132	194	133
rect	194	132	195	133
rect	195	132	196	133
rect	196	132	197	133
rect	197	132	198	133
rect	198	132	199	133
rect	199	132	200	133
rect	200	132	201	133
rect	201	132	202	133
rect	202	132	203	133
rect	203	132	204	133
rect	204	132	205	133
rect	205	132	206	133
rect	206	132	207	133
rect	207	132	208	133
rect	208	132	209	133
rect	209	132	210	133
rect	210	132	211	133
rect	211	132	212	133
rect	212	132	213	133
rect	213	132	214	133
rect	214	132	215	133
rect	215	132	216	133
rect	216	132	217	133
rect	217	132	218	133
rect	218	132	219	133
rect	219	132	220	133
rect	220	132	221	133
rect	221	132	222	133
rect	222	132	223	133
rect	223	132	224	133
rect	224	132	225	133
rect	225	132	226	133
rect	226	132	227	133
rect	227	132	228	133
rect	228	132	229	133
rect	229	132	230	133
rect	230	132	231	133
rect	231	132	232	133
rect	232	132	233	133
rect	233	132	234	133
rect	234	132	235	133
rect	235	132	236	133
rect	236	132	237	133
rect	237	132	238	133
rect	238	132	239	133
rect	239	132	240	133
rect	240	132	241	133
rect	241	132	242	133
rect	242	132	243	133
rect	243	132	244	133
rect	244	132	245	133
rect	245	132	246	133
rect	246	132	247	133
rect	247	132	248	133
rect	248	132	249	133
rect	249	132	250	133
rect	250	132	251	133
rect	251	132	252	133
rect	252	132	253	133
rect	253	132	254	133
rect	254	132	255	133
rect	255	132	256	133
rect	256	132	257	133
rect	257	132	258	133
rect	258	132	259	133
rect	259	132	260	133
rect	260	132	261	133
rect	261	132	262	133
rect	262	132	263	133
rect	263	132	264	133
rect	264	132	265	133
rect	265	132	266	133
rect	266	132	267	133
rect	267	132	268	133
rect	268	132	269	133
rect	269	132	270	133
rect	270	132	271	133
rect	271	132	272	133
rect	272	132	273	133
rect	273	132	274	133
rect	274	132	275	133
rect	275	132	276	133
rect	276	132	277	133
rect	277	132	278	133
rect	278	132	279	133
rect	279	132	280	133
rect	280	132	281	133
rect	281	132	282	133
rect	282	132	283	133
rect	283	132	284	133
rect	284	132	285	133
rect	285	132	286	133
rect	286	132	287	133
rect	287	132	288	133
rect	288	132	289	133
rect	289	132	290	133
rect	290	132	291	133
rect	291	132	292	133
rect	292	132	293	133
rect	293	132	294	133
rect	294	132	295	133
rect	295	132	296	133
rect	296	132	297	133
rect	297	132	298	133
rect	298	132	299	133
rect	299	132	300	133
rect	300	132	301	133
rect	301	132	302	133
rect	302	132	303	133
rect	303	132	304	133
rect	304	132	305	133
rect	305	132	306	133
rect	306	132	307	133
rect	307	132	308	133
rect	308	132	309	133
rect	309	132	310	133
rect	310	132	311	133
rect	311	132	312	133
rect	312	132	313	133
rect	313	132	314	133
rect	314	132	315	133
rect	315	132	316	133
rect	316	132	317	133
rect	317	132	318	133
rect	318	132	319	133
rect	319	132	320	133
rect	320	132	321	133
rect	321	132	322	133
rect	322	132	323	133
rect	323	132	324	133
rect	324	132	325	133
rect	325	132	326	133
rect	326	132	327	133
rect	327	132	328	133
rect	328	132	329	133
rect	329	132	330	133
rect	330	132	331	133
rect	331	132	332	133
rect	332	132	333	133
rect	333	132	334	133
rect	334	132	335	133
rect	335	132	336	133
rect	336	132	337	133
rect	337	132	338	133
rect	338	132	339	133
rect	339	132	340	133
rect	340	132	341	133
rect	341	132	342	133
rect	342	132	343	133
rect	343	132	344	133
rect	344	132	345	133
rect	345	132	346	133
rect	346	132	347	133
rect	347	132	348	133
rect	348	132	349	133
rect	349	132	350	133
rect	350	132	351	133
rect	351	132	352	133
rect	352	132	353	133
rect	353	132	354	133
rect	354	132	355	133
rect	355	132	356	133
rect	356	132	357	133
rect	357	132	358	133
rect	358	132	359	133
rect	359	132	360	133
rect	360	132	361	133
rect	361	132	362	133
rect	362	132	363	133
rect	363	132	364	133
rect	364	132	365	133
rect	365	132	366	133
rect	366	132	367	133
rect	367	132	368	133
rect	368	132	369	133
rect	369	132	370	133
rect	370	132	371	133
rect	371	132	372	133
rect	372	132	373	133
rect	373	132	374	133
rect	374	132	375	133
rect	375	132	376	133
rect	376	132	377	133
rect	377	132	378	133
rect	378	132	379	133
rect	379	132	380	133
rect	380	132	381	133
rect	381	132	382	133
rect	382	132	383	133
rect	383	132	384	133
rect	384	132	385	133
rect	385	132	386	133
rect	386	132	387	133
rect	387	132	388	133
rect	388	132	389	133
rect	389	132	390	133
rect	390	132	391	133
rect	391	132	392	133
rect	392	132	393	133
rect	393	132	394	133
rect	394	132	395	133
rect	395	132	396	133
rect	396	132	397	133
rect	397	132	398	133
rect	398	132	399	133
rect	399	132	400	133
rect	400	132	401	133
rect	401	132	402	133
rect	402	132	403	133
rect	403	132	404	133
rect	405	132	406	133
rect	406	132	407	133
rect	407	132	408	133
rect	408	132	409	133
rect	409	132	410	133
rect	410	132	411	133
rect	412	132	413	133
rect	413	132	414	133
rect	414	132	415	133
rect	415	132	416	133
rect	416	132	417	133
rect	417	132	418	133
rect	418	132	419	133
rect	419	132	420	133
rect	420	132	421	133
rect	0	133	1	134
rect	1	133	2	134
rect	2	133	3	134
rect	3	133	4	134
rect	4	133	5	134
rect	5	133	6	134
rect	7	133	8	134
rect	8	133	9	134
rect	9	133	10	134
rect	10	133	11	134
rect	11	133	12	134
rect	12	133	13	134
rect	14	133	15	134
rect	15	133	16	134
rect	16	133	17	134
rect	17	133	18	134
rect	18	133	19	134
rect	19	133	20	134
rect	20	133	21	134
rect	21	133	22	134
rect	22	133	23	134
rect	23	133	24	134
rect	24	133	25	134
rect	25	133	26	134
rect	26	133	27	134
rect	27	133	28	134
rect	28	133	29	134
rect	29	133	30	134
rect	30	133	31	134
rect	31	133	32	134
rect	32	133	33	134
rect	33	133	34	134
rect	34	133	35	134
rect	35	133	36	134
rect	36	133	37	134
rect	37	133	38	134
rect	38	133	39	134
rect	39	133	40	134
rect	40	133	41	134
rect	41	133	42	134
rect	42	133	43	134
rect	43	133	44	134
rect	44	133	45	134
rect	45	133	46	134
rect	46	133	47	134
rect	47	133	48	134
rect	48	133	49	134
rect	49	133	50	134
rect	51	133	52	134
rect	52	133	53	134
rect	53	133	54	134
rect	54	133	55	134
rect	55	133	56	134
rect	56	133	57	134
rect	57	133	58	134
rect	58	133	59	134
rect	59	133	60	134
rect	60	133	61	134
rect	61	133	62	134
rect	62	133	63	134
rect	63	133	64	134
rect	64	133	65	134
rect	65	133	66	134
rect	66	133	67	134
rect	67	133	68	134
rect	68	133	69	134
rect	69	133	70	134
rect	70	133	71	134
rect	71	133	72	134
rect	72	133	73	134
rect	73	133	74	134
rect	74	133	75	134
rect	75	133	76	134
rect	76	133	77	134
rect	77	133	78	134
rect	79	133	80	134
rect	80	133	81	134
rect	81	133	82	134
rect	82	133	83	134
rect	83	133	84	134
rect	84	133	85	134
rect	85	133	86	134
rect	86	133	87	134
rect	87	133	88	134
rect	88	133	89	134
rect	89	133	90	134
rect	90	133	91	134
rect	91	133	92	134
rect	92	133	93	134
rect	93	133	94	134
rect	94	133	95	134
rect	95	133	96	134
rect	96	133	97	134
rect	97	133	98	134
rect	98	133	99	134
rect	99	133	100	134
rect	101	133	102	134
rect	102	133	103	134
rect	103	133	104	134
rect	104	133	105	134
rect	105	133	106	134
rect	106	133	107	134
rect	108	133	109	134
rect	109	133	110	134
rect	110	133	111	134
rect	111	133	112	134
rect	112	133	113	134
rect	113	133	114	134
rect	114	133	115	134
rect	115	133	116	134
rect	116	133	117	134
rect	117	133	118	134
rect	118	133	119	134
rect	119	133	120	134
rect	120	133	121	134
rect	121	133	122	134
rect	122	133	123	134
rect	123	133	124	134
rect	124	133	125	134
rect	125	133	126	134
rect	126	133	127	134
rect	127	133	128	134
rect	128	133	129	134
rect	129	133	130	134
rect	130	133	131	134
rect	131	133	132	134
rect	132	133	133	134
rect	133	133	134	134
rect	134	133	135	134
rect	135	133	136	134
rect	136	133	137	134
rect	137	133	138	134
rect	138	133	139	134
rect	139	133	140	134
rect	140	133	141	134
rect	141	133	142	134
rect	142	133	143	134
rect	143	133	144	134
rect	145	133	146	134
rect	146	133	147	134
rect	147	133	148	134
rect	148	133	149	134
rect	149	133	150	134
rect	150	133	151	134
rect	151	133	152	134
rect	152	133	153	134
rect	153	133	154	134
rect	154	133	155	134
rect	155	133	156	134
rect	156	133	157	134
rect	157	133	158	134
rect	158	133	159	134
rect	159	133	160	134
rect	160	133	161	134
rect	161	133	162	134
rect	162	133	163	134
rect	163	133	164	134
rect	164	133	165	134
rect	165	133	166	134
rect	167	133	168	134
rect	168	133	169	134
rect	169	133	170	134
rect	170	133	171	134
rect	171	133	172	134
rect	172	133	173	134
rect	173	133	174	134
rect	174	133	175	134
rect	175	133	176	134
rect	176	133	177	134
rect	177	133	178	134
rect	178	133	179	134
rect	179	133	180	134
rect	180	133	181	134
rect	181	133	182	134
rect	182	133	183	134
rect	183	133	184	134
rect	184	133	185	134
rect	185	133	186	134
rect	186	133	187	134
rect	187	133	188	134
rect	188	133	189	134
rect	189	133	190	134
rect	190	133	191	134
rect	191	133	192	134
rect	192	133	193	134
rect	193	133	194	134
rect	194	133	195	134
rect	195	133	196	134
rect	196	133	197	134
rect	197	133	198	134
rect	198	133	199	134
rect	199	133	200	134
rect	200	133	201	134
rect	201	133	202	134
rect	202	133	203	134
rect	203	133	204	134
rect	204	133	205	134
rect	205	133	206	134
rect	206	133	207	134
rect	207	133	208	134
rect	208	133	209	134
rect	209	133	210	134
rect	210	133	211	134
rect	211	133	212	134
rect	212	133	213	134
rect	213	133	214	134
rect	214	133	215	134
rect	215	133	216	134
rect	216	133	217	134
rect	217	133	218	134
rect	218	133	219	134
rect	219	133	220	134
rect	220	133	221	134
rect	221	133	222	134
rect	222	133	223	134
rect	223	133	224	134
rect	224	133	225	134
rect	225	133	226	134
rect	226	133	227	134
rect	227	133	228	134
rect	228	133	229	134
rect	229	133	230	134
rect	230	133	231	134
rect	231	133	232	134
rect	232	133	233	134
rect	233	133	234	134
rect	234	133	235	134
rect	235	133	236	134
rect	236	133	237	134
rect	237	133	238	134
rect	238	133	239	134
rect	239	133	240	134
rect	240	133	241	134
rect	241	133	242	134
rect	242	133	243	134
rect	243	133	244	134
rect	244	133	245	134
rect	245	133	246	134
rect	246	133	247	134
rect	247	133	248	134
rect	248	133	249	134
rect	249	133	250	134
rect	250	133	251	134
rect	251	133	252	134
rect	252	133	253	134
rect	253	133	254	134
rect	254	133	255	134
rect	255	133	256	134
rect	256	133	257	134
rect	257	133	258	134
rect	258	133	259	134
rect	259	133	260	134
rect	260	133	261	134
rect	261	133	262	134
rect	262	133	263	134
rect	263	133	264	134
rect	264	133	265	134
rect	265	133	266	134
rect	266	133	267	134
rect	267	133	268	134
rect	268	133	269	134
rect	269	133	270	134
rect	270	133	271	134
rect	271	133	272	134
rect	272	133	273	134
rect	273	133	274	134
rect	274	133	275	134
rect	275	133	276	134
rect	276	133	277	134
rect	277	133	278	134
rect	278	133	279	134
rect	279	133	280	134
rect	280	133	281	134
rect	281	133	282	134
rect	282	133	283	134
rect	283	133	284	134
rect	284	133	285	134
rect	285	133	286	134
rect	286	133	287	134
rect	287	133	288	134
rect	288	133	289	134
rect	289	133	290	134
rect	290	133	291	134
rect	291	133	292	134
rect	292	133	293	134
rect	293	133	294	134
rect	294	133	295	134
rect	295	133	296	134
rect	296	133	297	134
rect	297	133	298	134
rect	298	133	299	134
rect	299	133	300	134
rect	300	133	301	134
rect	301	133	302	134
rect	302	133	303	134
rect	303	133	304	134
rect	304	133	305	134
rect	305	133	306	134
rect	306	133	307	134
rect	307	133	308	134
rect	308	133	309	134
rect	309	133	310	134
rect	310	133	311	134
rect	311	133	312	134
rect	312	133	313	134
rect	313	133	314	134
rect	314	133	315	134
rect	315	133	316	134
rect	316	133	317	134
rect	317	133	318	134
rect	318	133	319	134
rect	319	133	320	134
rect	320	133	321	134
rect	321	133	322	134
rect	322	133	323	134
rect	323	133	324	134
rect	324	133	325	134
rect	325	133	326	134
rect	326	133	327	134
rect	327	133	328	134
rect	328	133	329	134
rect	329	133	330	134
rect	330	133	331	134
rect	331	133	332	134
rect	332	133	333	134
rect	333	133	334	134
rect	334	133	335	134
rect	335	133	336	134
rect	336	133	337	134
rect	337	133	338	134
rect	338	133	339	134
rect	339	133	340	134
rect	340	133	341	134
rect	341	133	342	134
rect	342	133	343	134
rect	343	133	344	134
rect	344	133	345	134
rect	345	133	346	134
rect	346	133	347	134
rect	347	133	348	134
rect	348	133	349	134
rect	349	133	350	134
rect	350	133	351	134
rect	351	133	352	134
rect	352	133	353	134
rect	353	133	354	134
rect	354	133	355	134
rect	355	133	356	134
rect	356	133	357	134
rect	357	133	358	134
rect	358	133	359	134
rect	359	133	360	134
rect	360	133	361	134
rect	361	133	362	134
rect	362	133	363	134
rect	363	133	364	134
rect	364	133	365	134
rect	365	133	366	134
rect	366	133	367	134
rect	367	133	368	134
rect	368	133	369	134
rect	369	133	370	134
rect	370	133	371	134
rect	371	133	372	134
rect	372	133	373	134
rect	373	133	374	134
rect	374	133	375	134
rect	375	133	376	134
rect	376	133	377	134
rect	377	133	378	134
rect	378	133	379	134
rect	379	133	380	134
rect	380	133	381	134
rect	381	133	382	134
rect	382	133	383	134
rect	383	133	384	134
rect	384	133	385	134
rect	385	133	386	134
rect	386	133	387	134
rect	387	133	388	134
rect	388	133	389	134
rect	389	133	390	134
rect	390	133	391	134
rect	391	133	392	134
rect	392	133	393	134
rect	393	133	394	134
rect	394	133	395	134
rect	395	133	396	134
rect	396	133	397	134
rect	397	133	398	134
rect	398	133	399	134
rect	399	133	400	134
rect	400	133	401	134
rect	401	133	402	134
rect	402	133	403	134
rect	403	133	404	134
rect	405	133	406	134
rect	406	133	407	134
rect	407	133	408	134
rect	408	133	409	134
rect	409	133	410	134
rect	410	133	411	134
rect	412	133	413	134
rect	413	133	414	134
rect	414	133	415	134
rect	415	133	416	134
rect	416	133	417	134
rect	417	133	418	134
rect	418	133	419	134
rect	419	133	420	134
rect	420	133	421	134
rect	0	157	1	158
rect	1	157	2	158
rect	2	157	3	158
rect	3	157	4	158
rect	4	157	5	158
rect	5	157	6	158
rect	7	157	8	158
rect	8	157	9	158
rect	9	157	10	158
rect	10	157	11	158
rect	11	157	12	158
rect	12	157	13	158
rect	14	157	15	158
rect	15	157	16	158
rect	16	157	17	158
rect	17	157	18	158
rect	18	157	19	158
rect	19	157	20	158
rect	21	157	22	158
rect	22	157	23	158
rect	23	157	24	158
rect	24	157	25	158
rect	25	157	26	158
rect	26	157	27	158
rect	28	157	29	158
rect	29	157	30	158
rect	30	157	31	158
rect	31	157	32	158
rect	32	157	33	158
rect	33	157	34	158
rect	34	157	35	158
rect	35	157	36	158
rect	36	157	37	158
rect	37	157	38	158
rect	38	157	39	158
rect	39	157	40	158
rect	40	157	41	158
rect	41	157	42	158
rect	42	157	43	158
rect	43	157	44	158
rect	44	157	45	158
rect	45	157	46	158
rect	46	157	47	158
rect	47	157	48	158
rect	48	157	49	158
rect	49	157	50	158
rect	50	157	51	158
rect	51	157	52	158
rect	52	157	53	158
rect	53	157	54	158
rect	54	157	55	158
rect	55	157	56	158
rect	56	157	57	158
rect	57	157	58	158
rect	58	157	59	158
rect	59	157	60	158
rect	60	157	61	158
rect	61	157	62	158
rect	62	157	63	158
rect	63	157	64	158
rect	64	157	65	158
rect	65	157	66	158
rect	66	157	67	158
rect	67	157	68	158
rect	68	157	69	158
rect	69	157	70	158
rect	70	157	71	158
rect	71	157	72	158
rect	72	157	73	158
rect	74	157	75	158
rect	75	157	76	158
rect	76	157	77	158
rect	77	157	78	158
rect	78	157	79	158
rect	79	157	80	158
rect	81	157	82	158
rect	82	157	83	158
rect	83	157	84	158
rect	84	157	85	158
rect	85	157	86	158
rect	86	157	87	158
rect	88	157	89	158
rect	89	157	90	158
rect	90	157	91	158
rect	91	157	92	158
rect	92	157	93	158
rect	93	157	94	158
rect	94	157	95	158
rect	95	157	96	158
rect	96	157	97	158
rect	97	157	98	158
rect	98	157	99	158
rect	99	157	100	158
rect	100	157	101	158
rect	101	157	102	158
rect	102	157	103	158
rect	103	157	104	158
rect	104	157	105	158
rect	105	157	106	158
rect	106	157	107	158
rect	107	157	108	158
rect	108	157	109	158
rect	109	157	110	158
rect	110	157	111	158
rect	111	157	112	158
rect	112	157	113	158
rect	113	157	114	158
rect	114	157	115	158
rect	115	157	116	158
rect	116	157	117	158
rect	117	157	118	158
rect	118	157	119	158
rect	119	157	120	158
rect	120	157	121	158
rect	121	157	122	158
rect	122	157	123	158
rect	123	157	124	158
rect	124	157	125	158
rect	125	157	126	158
rect	126	157	127	158
rect	127	157	128	158
rect	128	157	129	158
rect	129	157	130	158
rect	130	157	131	158
rect	131	157	132	158
rect	132	157	133	158
rect	133	157	134	158
rect	134	157	135	158
rect	135	157	136	158
rect	136	157	137	158
rect	137	157	138	158
rect	138	157	139	158
rect	139	157	140	158
rect	140	157	141	158
rect	141	157	142	158
rect	142	157	143	158
rect	143	157	144	158
rect	144	157	145	158
rect	145	157	146	158
rect	146	157	147	158
rect	147	157	148	158
rect	148	157	149	158
rect	149	157	150	158
rect	150	157	151	158
rect	151	157	152	158
rect	152	157	153	158
rect	153	157	154	158
rect	154	157	155	158
rect	155	157	156	158
rect	156	157	157	158
rect	157	157	158	158
rect	158	157	159	158
rect	159	157	160	158
rect	160	157	161	158
rect	161	157	162	158
rect	162	157	163	158
rect	163	157	164	158
rect	164	157	165	158
rect	165	157	166	158
rect	166	157	167	158
rect	167	157	168	158
rect	168	157	169	158
rect	169	157	170	158
rect	170	157	171	158
rect	171	157	172	158
rect	172	157	173	158
rect	173	157	174	158
rect	174	157	175	158
rect	176	157	177	158
rect	177	157	178	158
rect	178	157	179	158
rect	179	157	180	158
rect	180	157	181	158
rect	181	157	182	158
rect	182	157	183	158
rect	183	157	184	158
rect	184	157	185	158
rect	185	157	186	158
rect	186	157	187	158
rect	187	157	188	158
rect	188	157	189	158
rect	189	157	190	158
rect	190	157	191	158
rect	191	157	192	158
rect	192	157	193	158
rect	193	157	194	158
rect	194	157	195	158
rect	195	157	196	158
rect	196	157	197	158
rect	197	157	198	158
rect	198	157	199	158
rect	199	157	200	158
rect	200	157	201	158
rect	201	157	202	158
rect	202	157	203	158
rect	203	157	204	158
rect	204	157	205	158
rect	205	157	206	158
rect	206	157	207	158
rect	207	157	208	158
rect	208	157	209	158
rect	209	157	210	158
rect	210	157	211	158
rect	211	157	212	158
rect	212	157	213	158
rect	213	157	214	158
rect	214	157	215	158
rect	215	157	216	158
rect	216	157	217	158
rect	217	157	218	158
rect	218	157	219	158
rect	219	157	220	158
rect	220	157	221	158
rect	221	157	222	158
rect	222	157	223	158
rect	223	157	224	158
rect	224	157	225	158
rect	225	157	226	158
rect	226	157	227	158
rect	227	157	228	158
rect	228	157	229	158
rect	229	157	230	158
rect	230	157	231	158
rect	231	157	232	158
rect	232	157	233	158
rect	233	157	234	158
rect	234	157	235	158
rect	235	157	236	158
rect	236	157	237	158
rect	237	157	238	158
rect	238	157	239	158
rect	239	157	240	158
rect	240	157	241	158
rect	241	157	242	158
rect	242	157	243	158
rect	243	157	244	158
rect	244	157	245	158
rect	245	157	246	158
rect	246	157	247	158
rect	247	157	248	158
rect	248	157	249	158
rect	249	157	250	158
rect	250	157	251	158
rect	251	157	252	158
rect	252	157	253	158
rect	253	157	254	158
rect	254	157	255	158
rect	255	157	256	158
rect	256	157	257	158
rect	257	157	258	158
rect	258	157	259	158
rect	259	157	260	158
rect	260	157	261	158
rect	261	157	262	158
rect	262	157	263	158
rect	263	157	264	158
rect	264	157	265	158
rect	265	157	266	158
rect	266	157	267	158
rect	267	157	268	158
rect	268	157	269	158
rect	269	157	270	158
rect	270	157	271	158
rect	271	157	272	158
rect	272	157	273	158
rect	273	157	274	158
rect	274	157	275	158
rect	275	157	276	158
rect	276	157	277	158
rect	277	157	278	158
rect	278	157	279	158
rect	279	157	280	158
rect	280	157	281	158
rect	281	157	282	158
rect	282	157	283	158
rect	283	157	284	158
rect	284	157	285	158
rect	285	157	286	158
rect	286	157	287	158
rect	287	157	288	158
rect	288	157	289	158
rect	289	157	290	158
rect	290	157	291	158
rect	291	157	292	158
rect	292	157	293	158
rect	293	157	294	158
rect	294	157	295	158
rect	295	157	296	158
rect	296	157	297	158
rect	297	157	298	158
rect	298	157	299	158
rect	299	157	300	158
rect	300	157	301	158
rect	301	157	302	158
rect	302	157	303	158
rect	303	157	304	158
rect	304	157	305	158
rect	305	157	306	158
rect	306	157	307	158
rect	307	157	308	158
rect	308	157	309	158
rect	309	157	310	158
rect	310	157	311	158
rect	311	157	312	158
rect	312	157	313	158
rect	313	157	314	158
rect	314	157	315	158
rect	315	157	316	158
rect	316	157	317	158
rect	317	157	318	158
rect	318	157	319	158
rect	319	157	320	158
rect	320	157	321	158
rect	321	157	322	158
rect	322	157	323	158
rect	323	157	324	158
rect	324	157	325	158
rect	325	157	326	158
rect	326	157	327	158
rect	327	157	328	158
rect	328	157	329	158
rect	329	157	330	158
rect	330	157	331	158
rect	331	157	332	158
rect	332	157	333	158
rect	333	157	334	158
rect	334	157	335	158
rect	335	157	336	158
rect	336	157	337	158
rect	337	157	338	158
rect	339	157	340	158
rect	340	157	341	158
rect	341	157	342	158
rect	342	157	343	158
rect	343	157	344	158
rect	344	157	345	158
rect	345	157	346	158
rect	346	157	347	158
rect	347	157	348	158
rect	348	157	349	158
rect	349	157	350	158
rect	350	157	351	158
rect	351	157	352	158
rect	352	157	353	158
rect	353	157	354	158
rect	354	157	355	158
rect	355	157	356	158
rect	356	157	357	158
rect	357	157	358	158
rect	358	157	359	158
rect	359	157	360	158
rect	360	157	361	158
rect	361	157	362	158
rect	362	157	363	158
rect	363	157	364	158
rect	364	157	365	158
rect	365	157	366	158
rect	366	157	367	158
rect	367	157	368	158
rect	368	157	369	158
rect	369	157	370	158
rect	370	157	371	158
rect	371	157	372	158
rect	372	157	373	158
rect	373	157	374	158
rect	374	157	375	158
rect	375	157	376	158
rect	376	157	377	158
rect	377	157	378	158
rect	378	157	379	158
rect	379	157	380	158
rect	380	157	381	158
rect	381	157	382	158
rect	382	157	383	158
rect	383	157	384	158
rect	384	157	385	158
rect	385	157	386	158
rect	386	157	387	158
rect	387	157	388	158
rect	388	157	389	158
rect	389	157	390	158
rect	390	157	391	158
rect	391	157	392	158
rect	392	157	393	158
rect	393	157	394	158
rect	394	157	395	158
rect	395	157	396	158
rect	396	157	397	158
rect	397	157	398	158
rect	398	157	399	158
rect	399	157	400	158
rect	400	157	401	158
rect	401	157	402	158
rect	403	157	404	158
rect	404	157	405	158
rect	405	157	406	158
rect	406	157	407	158
rect	407	157	408	158
rect	408	157	409	158
rect	409	157	410	158
rect	410	157	411	158
rect	411	157	412	158
rect	412	157	413	158
rect	413	157	414	158
rect	414	157	415	158
rect	0	158	1	159
rect	1	158	2	159
rect	2	158	3	159
rect	3	158	4	159
rect	4	158	5	159
rect	5	158	6	159
rect	7	158	8	159
rect	8	158	9	159
rect	9	158	10	159
rect	10	158	11	159
rect	11	158	12	159
rect	12	158	13	159
rect	14	158	15	159
rect	15	158	16	159
rect	16	158	17	159
rect	17	158	18	159
rect	18	158	19	159
rect	19	158	20	159
rect	21	158	22	159
rect	22	158	23	159
rect	23	158	24	159
rect	24	158	25	159
rect	25	158	26	159
rect	26	158	27	159
rect	28	158	29	159
rect	29	158	30	159
rect	30	158	31	159
rect	31	158	32	159
rect	32	158	33	159
rect	33	158	34	159
rect	34	158	35	159
rect	35	158	36	159
rect	36	158	37	159
rect	37	158	38	159
rect	38	158	39	159
rect	39	158	40	159
rect	40	158	41	159
rect	41	158	42	159
rect	42	158	43	159
rect	43	158	44	159
rect	44	158	45	159
rect	45	158	46	159
rect	46	158	47	159
rect	47	158	48	159
rect	48	158	49	159
rect	49	158	50	159
rect	50	158	51	159
rect	51	158	52	159
rect	52	158	53	159
rect	53	158	54	159
rect	54	158	55	159
rect	55	158	56	159
rect	56	158	57	159
rect	57	158	58	159
rect	58	158	59	159
rect	59	158	60	159
rect	60	158	61	159
rect	61	158	62	159
rect	62	158	63	159
rect	63	158	64	159
rect	64	158	65	159
rect	65	158	66	159
rect	66	158	67	159
rect	67	158	68	159
rect	68	158	69	159
rect	69	158	70	159
rect	70	158	71	159
rect	71	158	72	159
rect	72	158	73	159
rect	74	158	75	159
rect	75	158	76	159
rect	76	158	77	159
rect	77	158	78	159
rect	78	158	79	159
rect	79	158	80	159
rect	81	158	82	159
rect	82	158	83	159
rect	83	158	84	159
rect	84	158	85	159
rect	85	158	86	159
rect	86	158	87	159
rect	88	158	89	159
rect	89	158	90	159
rect	90	158	91	159
rect	91	158	92	159
rect	92	158	93	159
rect	93	158	94	159
rect	94	158	95	159
rect	95	158	96	159
rect	96	158	97	159
rect	97	158	98	159
rect	98	158	99	159
rect	99	158	100	159
rect	100	158	101	159
rect	101	158	102	159
rect	102	158	103	159
rect	103	158	104	159
rect	104	158	105	159
rect	105	158	106	159
rect	106	158	107	159
rect	107	158	108	159
rect	108	158	109	159
rect	109	158	110	159
rect	110	158	111	159
rect	111	158	112	159
rect	112	158	113	159
rect	113	158	114	159
rect	114	158	115	159
rect	115	158	116	159
rect	116	158	117	159
rect	117	158	118	159
rect	118	158	119	159
rect	119	158	120	159
rect	120	158	121	159
rect	121	158	122	159
rect	122	158	123	159
rect	123	158	124	159
rect	124	158	125	159
rect	125	158	126	159
rect	126	158	127	159
rect	127	158	128	159
rect	128	158	129	159
rect	129	158	130	159
rect	130	158	131	159
rect	131	158	132	159
rect	132	158	133	159
rect	133	158	134	159
rect	134	158	135	159
rect	135	158	136	159
rect	136	158	137	159
rect	137	158	138	159
rect	138	158	139	159
rect	139	158	140	159
rect	140	158	141	159
rect	141	158	142	159
rect	142	158	143	159
rect	143	158	144	159
rect	144	158	145	159
rect	145	158	146	159
rect	146	158	147	159
rect	147	158	148	159
rect	148	158	149	159
rect	149	158	150	159
rect	150	158	151	159
rect	151	158	152	159
rect	152	158	153	159
rect	153	158	154	159
rect	154	158	155	159
rect	155	158	156	159
rect	156	158	157	159
rect	157	158	158	159
rect	158	158	159	159
rect	159	158	160	159
rect	160	158	161	159
rect	161	158	162	159
rect	162	158	163	159
rect	163	158	164	159
rect	164	158	165	159
rect	165	158	166	159
rect	166	158	167	159
rect	167	158	168	159
rect	168	158	169	159
rect	169	158	170	159
rect	170	158	171	159
rect	171	158	172	159
rect	172	158	173	159
rect	173	158	174	159
rect	174	158	175	159
rect	176	158	177	159
rect	177	158	178	159
rect	178	158	179	159
rect	179	158	180	159
rect	180	158	181	159
rect	181	158	182	159
rect	182	158	183	159
rect	183	158	184	159
rect	184	158	185	159
rect	185	158	186	159
rect	186	158	187	159
rect	187	158	188	159
rect	188	158	189	159
rect	189	158	190	159
rect	190	158	191	159
rect	191	158	192	159
rect	192	158	193	159
rect	193	158	194	159
rect	194	158	195	159
rect	195	158	196	159
rect	196	158	197	159
rect	197	158	198	159
rect	198	158	199	159
rect	199	158	200	159
rect	200	158	201	159
rect	201	158	202	159
rect	202	158	203	159
rect	203	158	204	159
rect	204	158	205	159
rect	205	158	206	159
rect	206	158	207	159
rect	207	158	208	159
rect	208	158	209	159
rect	209	158	210	159
rect	210	158	211	159
rect	211	158	212	159
rect	212	158	213	159
rect	213	158	214	159
rect	214	158	215	159
rect	215	158	216	159
rect	216	158	217	159
rect	217	158	218	159
rect	218	158	219	159
rect	219	158	220	159
rect	220	158	221	159
rect	221	158	222	159
rect	222	158	223	159
rect	223	158	224	159
rect	224	158	225	159
rect	225	158	226	159
rect	226	158	227	159
rect	227	158	228	159
rect	228	158	229	159
rect	229	158	230	159
rect	230	158	231	159
rect	231	158	232	159
rect	232	158	233	159
rect	233	158	234	159
rect	234	158	235	159
rect	235	158	236	159
rect	236	158	237	159
rect	237	158	238	159
rect	238	158	239	159
rect	239	158	240	159
rect	240	158	241	159
rect	241	158	242	159
rect	242	158	243	159
rect	243	158	244	159
rect	244	158	245	159
rect	245	158	246	159
rect	246	158	247	159
rect	247	158	248	159
rect	248	158	249	159
rect	249	158	250	159
rect	250	158	251	159
rect	251	158	252	159
rect	252	158	253	159
rect	253	158	254	159
rect	254	158	255	159
rect	255	158	256	159
rect	256	158	257	159
rect	257	158	258	159
rect	258	158	259	159
rect	259	158	260	159
rect	260	158	261	159
rect	261	158	262	159
rect	262	158	263	159
rect	263	158	264	159
rect	264	158	265	159
rect	265	158	266	159
rect	266	158	267	159
rect	267	158	268	159
rect	268	158	269	159
rect	269	158	270	159
rect	270	158	271	159
rect	271	158	272	159
rect	272	158	273	159
rect	273	158	274	159
rect	274	158	275	159
rect	275	158	276	159
rect	276	158	277	159
rect	277	158	278	159
rect	278	158	279	159
rect	279	158	280	159
rect	280	158	281	159
rect	281	158	282	159
rect	282	158	283	159
rect	283	158	284	159
rect	284	158	285	159
rect	285	158	286	159
rect	286	158	287	159
rect	287	158	288	159
rect	288	158	289	159
rect	289	158	290	159
rect	290	158	291	159
rect	291	158	292	159
rect	292	158	293	159
rect	293	158	294	159
rect	294	158	295	159
rect	295	158	296	159
rect	296	158	297	159
rect	297	158	298	159
rect	298	158	299	159
rect	299	158	300	159
rect	300	158	301	159
rect	301	158	302	159
rect	302	158	303	159
rect	303	158	304	159
rect	304	158	305	159
rect	305	158	306	159
rect	306	158	307	159
rect	307	158	308	159
rect	308	158	309	159
rect	309	158	310	159
rect	310	158	311	159
rect	311	158	312	159
rect	312	158	313	159
rect	313	158	314	159
rect	314	158	315	159
rect	315	158	316	159
rect	316	158	317	159
rect	317	158	318	159
rect	318	158	319	159
rect	319	158	320	159
rect	320	158	321	159
rect	321	158	322	159
rect	322	158	323	159
rect	323	158	324	159
rect	324	158	325	159
rect	325	158	326	159
rect	326	158	327	159
rect	327	158	328	159
rect	328	158	329	159
rect	329	158	330	159
rect	330	158	331	159
rect	331	158	332	159
rect	332	158	333	159
rect	333	158	334	159
rect	334	158	335	159
rect	335	158	336	159
rect	336	158	337	159
rect	337	158	338	159
rect	339	158	340	159
rect	340	158	341	159
rect	341	158	342	159
rect	342	158	343	159
rect	343	158	344	159
rect	344	158	345	159
rect	345	158	346	159
rect	346	158	347	159
rect	347	158	348	159
rect	348	158	349	159
rect	349	158	350	159
rect	350	158	351	159
rect	351	158	352	159
rect	352	158	353	159
rect	353	158	354	159
rect	354	158	355	159
rect	355	158	356	159
rect	356	158	357	159
rect	357	158	358	159
rect	358	158	359	159
rect	359	158	360	159
rect	360	158	361	159
rect	361	158	362	159
rect	362	158	363	159
rect	363	158	364	159
rect	364	158	365	159
rect	365	158	366	159
rect	366	158	367	159
rect	367	158	368	159
rect	368	158	369	159
rect	369	158	370	159
rect	370	158	371	159
rect	371	158	372	159
rect	372	158	373	159
rect	373	158	374	159
rect	374	158	375	159
rect	375	158	376	159
rect	376	158	377	159
rect	377	158	378	159
rect	378	158	379	159
rect	379	158	380	159
rect	380	158	381	159
rect	381	158	382	159
rect	382	158	383	159
rect	383	158	384	159
rect	384	158	385	159
rect	385	158	386	159
rect	386	158	387	159
rect	387	158	388	159
rect	388	158	389	159
rect	389	158	390	159
rect	390	158	391	159
rect	391	158	392	159
rect	392	158	393	159
rect	393	158	394	159
rect	394	158	395	159
rect	395	158	396	159
rect	396	158	397	159
rect	397	158	398	159
rect	398	158	399	159
rect	399	158	400	159
rect	400	158	401	159
rect	401	158	402	159
rect	403	158	404	159
rect	404	158	405	159
rect	405	158	406	159
rect	406	158	407	159
rect	407	158	408	159
rect	408	158	409	159
rect	409	158	410	159
rect	410	158	411	159
rect	411	158	412	159
rect	412	158	413	159
rect	413	158	414	159
rect	414	158	415	159
rect	0	159	1	160
rect	1	159	2	160
rect	2	159	3	160
rect	3	159	4	160
rect	4	159	5	160
rect	5	159	6	160
rect	7	159	8	160
rect	8	159	9	160
rect	9	159	10	160
rect	10	159	11	160
rect	11	159	12	160
rect	12	159	13	160
rect	14	159	15	160
rect	15	159	16	160
rect	16	159	17	160
rect	17	159	18	160
rect	18	159	19	160
rect	19	159	20	160
rect	21	159	22	160
rect	22	159	23	160
rect	23	159	24	160
rect	24	159	25	160
rect	25	159	26	160
rect	26	159	27	160
rect	28	159	29	160
rect	29	159	30	160
rect	30	159	31	160
rect	31	159	32	160
rect	32	159	33	160
rect	33	159	34	160
rect	34	159	35	160
rect	35	159	36	160
rect	36	159	37	160
rect	37	159	38	160
rect	38	159	39	160
rect	39	159	40	160
rect	40	159	41	160
rect	41	159	42	160
rect	42	159	43	160
rect	43	159	44	160
rect	44	159	45	160
rect	45	159	46	160
rect	46	159	47	160
rect	47	159	48	160
rect	48	159	49	160
rect	49	159	50	160
rect	50	159	51	160
rect	51	159	52	160
rect	52	159	53	160
rect	53	159	54	160
rect	54	159	55	160
rect	55	159	56	160
rect	56	159	57	160
rect	57	159	58	160
rect	58	159	59	160
rect	59	159	60	160
rect	60	159	61	160
rect	61	159	62	160
rect	62	159	63	160
rect	63	159	64	160
rect	64	159	65	160
rect	65	159	66	160
rect	66	159	67	160
rect	67	159	68	160
rect	68	159	69	160
rect	69	159	70	160
rect	70	159	71	160
rect	71	159	72	160
rect	72	159	73	160
rect	74	159	75	160
rect	75	159	76	160
rect	76	159	77	160
rect	77	159	78	160
rect	78	159	79	160
rect	79	159	80	160
rect	81	159	82	160
rect	82	159	83	160
rect	83	159	84	160
rect	84	159	85	160
rect	85	159	86	160
rect	86	159	87	160
rect	88	159	89	160
rect	89	159	90	160
rect	90	159	91	160
rect	91	159	92	160
rect	92	159	93	160
rect	93	159	94	160
rect	94	159	95	160
rect	95	159	96	160
rect	96	159	97	160
rect	97	159	98	160
rect	98	159	99	160
rect	99	159	100	160
rect	100	159	101	160
rect	101	159	102	160
rect	102	159	103	160
rect	103	159	104	160
rect	104	159	105	160
rect	105	159	106	160
rect	106	159	107	160
rect	107	159	108	160
rect	108	159	109	160
rect	109	159	110	160
rect	110	159	111	160
rect	111	159	112	160
rect	112	159	113	160
rect	113	159	114	160
rect	114	159	115	160
rect	115	159	116	160
rect	116	159	117	160
rect	117	159	118	160
rect	118	159	119	160
rect	119	159	120	160
rect	120	159	121	160
rect	121	159	122	160
rect	122	159	123	160
rect	123	159	124	160
rect	124	159	125	160
rect	125	159	126	160
rect	126	159	127	160
rect	127	159	128	160
rect	128	159	129	160
rect	129	159	130	160
rect	130	159	131	160
rect	131	159	132	160
rect	132	159	133	160
rect	133	159	134	160
rect	134	159	135	160
rect	135	159	136	160
rect	136	159	137	160
rect	137	159	138	160
rect	138	159	139	160
rect	139	159	140	160
rect	140	159	141	160
rect	141	159	142	160
rect	142	159	143	160
rect	143	159	144	160
rect	144	159	145	160
rect	145	159	146	160
rect	146	159	147	160
rect	147	159	148	160
rect	148	159	149	160
rect	149	159	150	160
rect	150	159	151	160
rect	151	159	152	160
rect	152	159	153	160
rect	153	159	154	160
rect	154	159	155	160
rect	155	159	156	160
rect	156	159	157	160
rect	157	159	158	160
rect	158	159	159	160
rect	159	159	160	160
rect	160	159	161	160
rect	161	159	162	160
rect	162	159	163	160
rect	163	159	164	160
rect	164	159	165	160
rect	165	159	166	160
rect	166	159	167	160
rect	167	159	168	160
rect	168	159	169	160
rect	169	159	170	160
rect	170	159	171	160
rect	171	159	172	160
rect	172	159	173	160
rect	173	159	174	160
rect	174	159	175	160
rect	176	159	177	160
rect	177	159	178	160
rect	178	159	179	160
rect	179	159	180	160
rect	180	159	181	160
rect	181	159	182	160
rect	182	159	183	160
rect	183	159	184	160
rect	184	159	185	160
rect	185	159	186	160
rect	186	159	187	160
rect	187	159	188	160
rect	188	159	189	160
rect	189	159	190	160
rect	190	159	191	160
rect	191	159	192	160
rect	192	159	193	160
rect	193	159	194	160
rect	194	159	195	160
rect	195	159	196	160
rect	196	159	197	160
rect	197	159	198	160
rect	198	159	199	160
rect	199	159	200	160
rect	200	159	201	160
rect	201	159	202	160
rect	202	159	203	160
rect	203	159	204	160
rect	204	159	205	160
rect	205	159	206	160
rect	206	159	207	160
rect	207	159	208	160
rect	208	159	209	160
rect	209	159	210	160
rect	210	159	211	160
rect	211	159	212	160
rect	212	159	213	160
rect	213	159	214	160
rect	214	159	215	160
rect	215	159	216	160
rect	216	159	217	160
rect	217	159	218	160
rect	218	159	219	160
rect	219	159	220	160
rect	220	159	221	160
rect	221	159	222	160
rect	222	159	223	160
rect	223	159	224	160
rect	224	159	225	160
rect	225	159	226	160
rect	226	159	227	160
rect	227	159	228	160
rect	228	159	229	160
rect	229	159	230	160
rect	230	159	231	160
rect	231	159	232	160
rect	232	159	233	160
rect	233	159	234	160
rect	234	159	235	160
rect	235	159	236	160
rect	236	159	237	160
rect	237	159	238	160
rect	238	159	239	160
rect	239	159	240	160
rect	240	159	241	160
rect	241	159	242	160
rect	242	159	243	160
rect	243	159	244	160
rect	244	159	245	160
rect	245	159	246	160
rect	246	159	247	160
rect	247	159	248	160
rect	248	159	249	160
rect	249	159	250	160
rect	250	159	251	160
rect	251	159	252	160
rect	252	159	253	160
rect	253	159	254	160
rect	254	159	255	160
rect	255	159	256	160
rect	256	159	257	160
rect	257	159	258	160
rect	258	159	259	160
rect	259	159	260	160
rect	260	159	261	160
rect	261	159	262	160
rect	262	159	263	160
rect	263	159	264	160
rect	264	159	265	160
rect	265	159	266	160
rect	266	159	267	160
rect	267	159	268	160
rect	268	159	269	160
rect	269	159	270	160
rect	270	159	271	160
rect	271	159	272	160
rect	272	159	273	160
rect	273	159	274	160
rect	274	159	275	160
rect	275	159	276	160
rect	276	159	277	160
rect	277	159	278	160
rect	278	159	279	160
rect	279	159	280	160
rect	280	159	281	160
rect	281	159	282	160
rect	282	159	283	160
rect	283	159	284	160
rect	284	159	285	160
rect	285	159	286	160
rect	286	159	287	160
rect	287	159	288	160
rect	288	159	289	160
rect	289	159	290	160
rect	290	159	291	160
rect	291	159	292	160
rect	292	159	293	160
rect	293	159	294	160
rect	294	159	295	160
rect	295	159	296	160
rect	296	159	297	160
rect	297	159	298	160
rect	298	159	299	160
rect	299	159	300	160
rect	300	159	301	160
rect	301	159	302	160
rect	302	159	303	160
rect	303	159	304	160
rect	304	159	305	160
rect	305	159	306	160
rect	306	159	307	160
rect	307	159	308	160
rect	308	159	309	160
rect	309	159	310	160
rect	310	159	311	160
rect	311	159	312	160
rect	312	159	313	160
rect	313	159	314	160
rect	314	159	315	160
rect	315	159	316	160
rect	316	159	317	160
rect	317	159	318	160
rect	318	159	319	160
rect	319	159	320	160
rect	320	159	321	160
rect	321	159	322	160
rect	322	159	323	160
rect	323	159	324	160
rect	324	159	325	160
rect	325	159	326	160
rect	326	159	327	160
rect	327	159	328	160
rect	328	159	329	160
rect	329	159	330	160
rect	330	159	331	160
rect	331	159	332	160
rect	332	159	333	160
rect	333	159	334	160
rect	334	159	335	160
rect	335	159	336	160
rect	336	159	337	160
rect	337	159	338	160
rect	339	159	340	160
rect	340	159	341	160
rect	341	159	342	160
rect	342	159	343	160
rect	343	159	344	160
rect	344	159	345	160
rect	345	159	346	160
rect	346	159	347	160
rect	347	159	348	160
rect	348	159	349	160
rect	349	159	350	160
rect	350	159	351	160
rect	351	159	352	160
rect	352	159	353	160
rect	353	159	354	160
rect	354	159	355	160
rect	355	159	356	160
rect	356	159	357	160
rect	357	159	358	160
rect	358	159	359	160
rect	359	159	360	160
rect	360	159	361	160
rect	361	159	362	160
rect	362	159	363	160
rect	363	159	364	160
rect	364	159	365	160
rect	365	159	366	160
rect	366	159	367	160
rect	367	159	368	160
rect	368	159	369	160
rect	369	159	370	160
rect	370	159	371	160
rect	371	159	372	160
rect	372	159	373	160
rect	373	159	374	160
rect	374	159	375	160
rect	375	159	376	160
rect	376	159	377	160
rect	377	159	378	160
rect	378	159	379	160
rect	379	159	380	160
rect	380	159	381	160
rect	381	159	382	160
rect	382	159	383	160
rect	383	159	384	160
rect	384	159	385	160
rect	385	159	386	160
rect	386	159	387	160
rect	387	159	388	160
rect	388	159	389	160
rect	389	159	390	160
rect	390	159	391	160
rect	391	159	392	160
rect	392	159	393	160
rect	393	159	394	160
rect	394	159	395	160
rect	395	159	396	160
rect	396	159	397	160
rect	397	159	398	160
rect	398	159	399	160
rect	399	159	400	160
rect	400	159	401	160
rect	401	159	402	160
rect	403	159	404	160
rect	404	159	405	160
rect	405	159	406	160
rect	406	159	407	160
rect	407	159	408	160
rect	408	159	409	160
rect	409	159	410	160
rect	410	159	411	160
rect	411	159	412	160
rect	412	159	413	160
rect	413	159	414	160
rect	414	159	415	160
rect	0	160	1	161
rect	1	160	2	161
rect	2	160	3	161
rect	3	160	4	161
rect	4	160	5	161
rect	5	160	6	161
rect	7	160	8	161
rect	8	160	9	161
rect	9	160	10	161
rect	10	160	11	161
rect	11	160	12	161
rect	12	160	13	161
rect	14	160	15	161
rect	15	160	16	161
rect	16	160	17	161
rect	17	160	18	161
rect	18	160	19	161
rect	19	160	20	161
rect	21	160	22	161
rect	22	160	23	161
rect	23	160	24	161
rect	24	160	25	161
rect	25	160	26	161
rect	26	160	27	161
rect	28	160	29	161
rect	29	160	30	161
rect	30	160	31	161
rect	31	160	32	161
rect	32	160	33	161
rect	33	160	34	161
rect	34	160	35	161
rect	35	160	36	161
rect	36	160	37	161
rect	37	160	38	161
rect	38	160	39	161
rect	39	160	40	161
rect	40	160	41	161
rect	41	160	42	161
rect	42	160	43	161
rect	43	160	44	161
rect	44	160	45	161
rect	45	160	46	161
rect	46	160	47	161
rect	47	160	48	161
rect	48	160	49	161
rect	49	160	50	161
rect	50	160	51	161
rect	51	160	52	161
rect	52	160	53	161
rect	53	160	54	161
rect	54	160	55	161
rect	55	160	56	161
rect	56	160	57	161
rect	57	160	58	161
rect	58	160	59	161
rect	59	160	60	161
rect	60	160	61	161
rect	61	160	62	161
rect	62	160	63	161
rect	63	160	64	161
rect	64	160	65	161
rect	65	160	66	161
rect	66	160	67	161
rect	67	160	68	161
rect	68	160	69	161
rect	69	160	70	161
rect	70	160	71	161
rect	71	160	72	161
rect	72	160	73	161
rect	74	160	75	161
rect	75	160	76	161
rect	76	160	77	161
rect	77	160	78	161
rect	78	160	79	161
rect	79	160	80	161
rect	81	160	82	161
rect	82	160	83	161
rect	83	160	84	161
rect	84	160	85	161
rect	85	160	86	161
rect	86	160	87	161
rect	88	160	89	161
rect	89	160	90	161
rect	90	160	91	161
rect	91	160	92	161
rect	92	160	93	161
rect	93	160	94	161
rect	94	160	95	161
rect	95	160	96	161
rect	96	160	97	161
rect	97	160	98	161
rect	98	160	99	161
rect	99	160	100	161
rect	100	160	101	161
rect	101	160	102	161
rect	102	160	103	161
rect	103	160	104	161
rect	104	160	105	161
rect	105	160	106	161
rect	106	160	107	161
rect	107	160	108	161
rect	108	160	109	161
rect	109	160	110	161
rect	110	160	111	161
rect	111	160	112	161
rect	112	160	113	161
rect	113	160	114	161
rect	114	160	115	161
rect	115	160	116	161
rect	116	160	117	161
rect	117	160	118	161
rect	118	160	119	161
rect	119	160	120	161
rect	120	160	121	161
rect	121	160	122	161
rect	122	160	123	161
rect	123	160	124	161
rect	124	160	125	161
rect	125	160	126	161
rect	126	160	127	161
rect	127	160	128	161
rect	128	160	129	161
rect	129	160	130	161
rect	130	160	131	161
rect	131	160	132	161
rect	132	160	133	161
rect	133	160	134	161
rect	134	160	135	161
rect	135	160	136	161
rect	136	160	137	161
rect	137	160	138	161
rect	138	160	139	161
rect	139	160	140	161
rect	140	160	141	161
rect	141	160	142	161
rect	142	160	143	161
rect	143	160	144	161
rect	144	160	145	161
rect	145	160	146	161
rect	146	160	147	161
rect	147	160	148	161
rect	148	160	149	161
rect	149	160	150	161
rect	150	160	151	161
rect	151	160	152	161
rect	152	160	153	161
rect	153	160	154	161
rect	154	160	155	161
rect	155	160	156	161
rect	156	160	157	161
rect	157	160	158	161
rect	158	160	159	161
rect	159	160	160	161
rect	160	160	161	161
rect	161	160	162	161
rect	162	160	163	161
rect	163	160	164	161
rect	164	160	165	161
rect	165	160	166	161
rect	166	160	167	161
rect	167	160	168	161
rect	168	160	169	161
rect	169	160	170	161
rect	170	160	171	161
rect	171	160	172	161
rect	172	160	173	161
rect	173	160	174	161
rect	174	160	175	161
rect	176	160	177	161
rect	177	160	178	161
rect	178	160	179	161
rect	179	160	180	161
rect	180	160	181	161
rect	181	160	182	161
rect	182	160	183	161
rect	183	160	184	161
rect	184	160	185	161
rect	185	160	186	161
rect	186	160	187	161
rect	187	160	188	161
rect	188	160	189	161
rect	189	160	190	161
rect	190	160	191	161
rect	191	160	192	161
rect	192	160	193	161
rect	193	160	194	161
rect	194	160	195	161
rect	195	160	196	161
rect	196	160	197	161
rect	197	160	198	161
rect	198	160	199	161
rect	199	160	200	161
rect	200	160	201	161
rect	201	160	202	161
rect	202	160	203	161
rect	203	160	204	161
rect	204	160	205	161
rect	205	160	206	161
rect	206	160	207	161
rect	207	160	208	161
rect	208	160	209	161
rect	209	160	210	161
rect	210	160	211	161
rect	211	160	212	161
rect	212	160	213	161
rect	213	160	214	161
rect	214	160	215	161
rect	215	160	216	161
rect	216	160	217	161
rect	217	160	218	161
rect	218	160	219	161
rect	219	160	220	161
rect	220	160	221	161
rect	221	160	222	161
rect	222	160	223	161
rect	223	160	224	161
rect	224	160	225	161
rect	225	160	226	161
rect	226	160	227	161
rect	227	160	228	161
rect	228	160	229	161
rect	229	160	230	161
rect	230	160	231	161
rect	231	160	232	161
rect	232	160	233	161
rect	233	160	234	161
rect	234	160	235	161
rect	235	160	236	161
rect	236	160	237	161
rect	237	160	238	161
rect	238	160	239	161
rect	239	160	240	161
rect	240	160	241	161
rect	241	160	242	161
rect	242	160	243	161
rect	243	160	244	161
rect	244	160	245	161
rect	245	160	246	161
rect	246	160	247	161
rect	247	160	248	161
rect	248	160	249	161
rect	249	160	250	161
rect	250	160	251	161
rect	251	160	252	161
rect	252	160	253	161
rect	253	160	254	161
rect	254	160	255	161
rect	255	160	256	161
rect	256	160	257	161
rect	257	160	258	161
rect	258	160	259	161
rect	259	160	260	161
rect	260	160	261	161
rect	261	160	262	161
rect	262	160	263	161
rect	263	160	264	161
rect	264	160	265	161
rect	265	160	266	161
rect	266	160	267	161
rect	267	160	268	161
rect	268	160	269	161
rect	269	160	270	161
rect	270	160	271	161
rect	271	160	272	161
rect	272	160	273	161
rect	273	160	274	161
rect	274	160	275	161
rect	275	160	276	161
rect	276	160	277	161
rect	277	160	278	161
rect	278	160	279	161
rect	279	160	280	161
rect	280	160	281	161
rect	281	160	282	161
rect	282	160	283	161
rect	283	160	284	161
rect	284	160	285	161
rect	285	160	286	161
rect	286	160	287	161
rect	287	160	288	161
rect	288	160	289	161
rect	289	160	290	161
rect	290	160	291	161
rect	291	160	292	161
rect	292	160	293	161
rect	293	160	294	161
rect	294	160	295	161
rect	295	160	296	161
rect	296	160	297	161
rect	297	160	298	161
rect	298	160	299	161
rect	299	160	300	161
rect	300	160	301	161
rect	301	160	302	161
rect	302	160	303	161
rect	303	160	304	161
rect	304	160	305	161
rect	305	160	306	161
rect	306	160	307	161
rect	307	160	308	161
rect	308	160	309	161
rect	309	160	310	161
rect	310	160	311	161
rect	311	160	312	161
rect	312	160	313	161
rect	313	160	314	161
rect	314	160	315	161
rect	315	160	316	161
rect	316	160	317	161
rect	317	160	318	161
rect	318	160	319	161
rect	319	160	320	161
rect	320	160	321	161
rect	321	160	322	161
rect	322	160	323	161
rect	323	160	324	161
rect	324	160	325	161
rect	325	160	326	161
rect	326	160	327	161
rect	327	160	328	161
rect	328	160	329	161
rect	329	160	330	161
rect	330	160	331	161
rect	331	160	332	161
rect	332	160	333	161
rect	333	160	334	161
rect	334	160	335	161
rect	335	160	336	161
rect	336	160	337	161
rect	337	160	338	161
rect	339	160	340	161
rect	340	160	341	161
rect	341	160	342	161
rect	342	160	343	161
rect	343	160	344	161
rect	344	160	345	161
rect	345	160	346	161
rect	346	160	347	161
rect	347	160	348	161
rect	348	160	349	161
rect	349	160	350	161
rect	350	160	351	161
rect	351	160	352	161
rect	352	160	353	161
rect	353	160	354	161
rect	354	160	355	161
rect	355	160	356	161
rect	356	160	357	161
rect	357	160	358	161
rect	358	160	359	161
rect	359	160	360	161
rect	360	160	361	161
rect	361	160	362	161
rect	362	160	363	161
rect	363	160	364	161
rect	364	160	365	161
rect	365	160	366	161
rect	366	160	367	161
rect	367	160	368	161
rect	368	160	369	161
rect	369	160	370	161
rect	370	160	371	161
rect	371	160	372	161
rect	372	160	373	161
rect	373	160	374	161
rect	374	160	375	161
rect	375	160	376	161
rect	376	160	377	161
rect	377	160	378	161
rect	378	160	379	161
rect	379	160	380	161
rect	380	160	381	161
rect	381	160	382	161
rect	382	160	383	161
rect	383	160	384	161
rect	384	160	385	161
rect	385	160	386	161
rect	386	160	387	161
rect	387	160	388	161
rect	388	160	389	161
rect	389	160	390	161
rect	390	160	391	161
rect	391	160	392	161
rect	392	160	393	161
rect	393	160	394	161
rect	394	160	395	161
rect	395	160	396	161
rect	396	160	397	161
rect	397	160	398	161
rect	398	160	399	161
rect	399	160	400	161
rect	400	160	401	161
rect	401	160	402	161
rect	403	160	404	161
rect	404	160	405	161
rect	405	160	406	161
rect	406	160	407	161
rect	407	160	408	161
rect	408	160	409	161
rect	409	160	410	161
rect	410	160	411	161
rect	411	160	412	161
rect	412	160	413	161
rect	413	160	414	161
rect	414	160	415	161
rect	0	161	1	162
rect	1	161	2	162
rect	2	161	3	162
rect	3	161	4	162
rect	4	161	5	162
rect	5	161	6	162
rect	7	161	8	162
rect	8	161	9	162
rect	9	161	10	162
rect	10	161	11	162
rect	11	161	12	162
rect	12	161	13	162
rect	14	161	15	162
rect	15	161	16	162
rect	16	161	17	162
rect	17	161	18	162
rect	18	161	19	162
rect	19	161	20	162
rect	21	161	22	162
rect	22	161	23	162
rect	23	161	24	162
rect	24	161	25	162
rect	25	161	26	162
rect	26	161	27	162
rect	28	161	29	162
rect	29	161	30	162
rect	30	161	31	162
rect	31	161	32	162
rect	32	161	33	162
rect	33	161	34	162
rect	34	161	35	162
rect	35	161	36	162
rect	36	161	37	162
rect	37	161	38	162
rect	38	161	39	162
rect	39	161	40	162
rect	40	161	41	162
rect	41	161	42	162
rect	42	161	43	162
rect	43	161	44	162
rect	44	161	45	162
rect	45	161	46	162
rect	46	161	47	162
rect	47	161	48	162
rect	48	161	49	162
rect	49	161	50	162
rect	50	161	51	162
rect	51	161	52	162
rect	52	161	53	162
rect	53	161	54	162
rect	54	161	55	162
rect	55	161	56	162
rect	56	161	57	162
rect	57	161	58	162
rect	58	161	59	162
rect	59	161	60	162
rect	60	161	61	162
rect	61	161	62	162
rect	62	161	63	162
rect	63	161	64	162
rect	64	161	65	162
rect	65	161	66	162
rect	66	161	67	162
rect	67	161	68	162
rect	68	161	69	162
rect	69	161	70	162
rect	70	161	71	162
rect	71	161	72	162
rect	72	161	73	162
rect	74	161	75	162
rect	75	161	76	162
rect	76	161	77	162
rect	77	161	78	162
rect	78	161	79	162
rect	79	161	80	162
rect	81	161	82	162
rect	82	161	83	162
rect	83	161	84	162
rect	84	161	85	162
rect	85	161	86	162
rect	86	161	87	162
rect	88	161	89	162
rect	89	161	90	162
rect	90	161	91	162
rect	91	161	92	162
rect	92	161	93	162
rect	93	161	94	162
rect	94	161	95	162
rect	95	161	96	162
rect	96	161	97	162
rect	97	161	98	162
rect	98	161	99	162
rect	99	161	100	162
rect	100	161	101	162
rect	101	161	102	162
rect	102	161	103	162
rect	103	161	104	162
rect	104	161	105	162
rect	105	161	106	162
rect	106	161	107	162
rect	107	161	108	162
rect	108	161	109	162
rect	109	161	110	162
rect	110	161	111	162
rect	111	161	112	162
rect	112	161	113	162
rect	113	161	114	162
rect	114	161	115	162
rect	115	161	116	162
rect	116	161	117	162
rect	117	161	118	162
rect	118	161	119	162
rect	119	161	120	162
rect	120	161	121	162
rect	121	161	122	162
rect	122	161	123	162
rect	123	161	124	162
rect	124	161	125	162
rect	125	161	126	162
rect	126	161	127	162
rect	127	161	128	162
rect	128	161	129	162
rect	129	161	130	162
rect	130	161	131	162
rect	131	161	132	162
rect	132	161	133	162
rect	133	161	134	162
rect	134	161	135	162
rect	135	161	136	162
rect	136	161	137	162
rect	137	161	138	162
rect	138	161	139	162
rect	139	161	140	162
rect	140	161	141	162
rect	141	161	142	162
rect	142	161	143	162
rect	143	161	144	162
rect	144	161	145	162
rect	145	161	146	162
rect	146	161	147	162
rect	147	161	148	162
rect	148	161	149	162
rect	149	161	150	162
rect	150	161	151	162
rect	151	161	152	162
rect	152	161	153	162
rect	153	161	154	162
rect	154	161	155	162
rect	155	161	156	162
rect	156	161	157	162
rect	157	161	158	162
rect	158	161	159	162
rect	159	161	160	162
rect	160	161	161	162
rect	161	161	162	162
rect	162	161	163	162
rect	163	161	164	162
rect	164	161	165	162
rect	165	161	166	162
rect	166	161	167	162
rect	167	161	168	162
rect	168	161	169	162
rect	169	161	170	162
rect	170	161	171	162
rect	171	161	172	162
rect	172	161	173	162
rect	173	161	174	162
rect	174	161	175	162
rect	176	161	177	162
rect	177	161	178	162
rect	178	161	179	162
rect	179	161	180	162
rect	180	161	181	162
rect	181	161	182	162
rect	182	161	183	162
rect	183	161	184	162
rect	184	161	185	162
rect	185	161	186	162
rect	186	161	187	162
rect	187	161	188	162
rect	188	161	189	162
rect	189	161	190	162
rect	190	161	191	162
rect	191	161	192	162
rect	192	161	193	162
rect	193	161	194	162
rect	194	161	195	162
rect	195	161	196	162
rect	196	161	197	162
rect	197	161	198	162
rect	198	161	199	162
rect	199	161	200	162
rect	200	161	201	162
rect	201	161	202	162
rect	202	161	203	162
rect	203	161	204	162
rect	204	161	205	162
rect	205	161	206	162
rect	206	161	207	162
rect	207	161	208	162
rect	208	161	209	162
rect	209	161	210	162
rect	210	161	211	162
rect	211	161	212	162
rect	212	161	213	162
rect	213	161	214	162
rect	214	161	215	162
rect	215	161	216	162
rect	216	161	217	162
rect	217	161	218	162
rect	218	161	219	162
rect	219	161	220	162
rect	220	161	221	162
rect	221	161	222	162
rect	222	161	223	162
rect	223	161	224	162
rect	224	161	225	162
rect	225	161	226	162
rect	226	161	227	162
rect	227	161	228	162
rect	228	161	229	162
rect	229	161	230	162
rect	230	161	231	162
rect	231	161	232	162
rect	232	161	233	162
rect	233	161	234	162
rect	234	161	235	162
rect	235	161	236	162
rect	236	161	237	162
rect	237	161	238	162
rect	238	161	239	162
rect	239	161	240	162
rect	240	161	241	162
rect	241	161	242	162
rect	242	161	243	162
rect	243	161	244	162
rect	244	161	245	162
rect	245	161	246	162
rect	246	161	247	162
rect	247	161	248	162
rect	248	161	249	162
rect	249	161	250	162
rect	250	161	251	162
rect	251	161	252	162
rect	252	161	253	162
rect	253	161	254	162
rect	254	161	255	162
rect	255	161	256	162
rect	256	161	257	162
rect	257	161	258	162
rect	258	161	259	162
rect	259	161	260	162
rect	260	161	261	162
rect	261	161	262	162
rect	262	161	263	162
rect	263	161	264	162
rect	264	161	265	162
rect	265	161	266	162
rect	266	161	267	162
rect	267	161	268	162
rect	268	161	269	162
rect	269	161	270	162
rect	270	161	271	162
rect	271	161	272	162
rect	272	161	273	162
rect	273	161	274	162
rect	274	161	275	162
rect	275	161	276	162
rect	276	161	277	162
rect	277	161	278	162
rect	278	161	279	162
rect	279	161	280	162
rect	280	161	281	162
rect	281	161	282	162
rect	282	161	283	162
rect	283	161	284	162
rect	284	161	285	162
rect	285	161	286	162
rect	286	161	287	162
rect	287	161	288	162
rect	288	161	289	162
rect	289	161	290	162
rect	290	161	291	162
rect	291	161	292	162
rect	292	161	293	162
rect	293	161	294	162
rect	294	161	295	162
rect	295	161	296	162
rect	296	161	297	162
rect	297	161	298	162
rect	298	161	299	162
rect	299	161	300	162
rect	300	161	301	162
rect	301	161	302	162
rect	302	161	303	162
rect	303	161	304	162
rect	304	161	305	162
rect	305	161	306	162
rect	306	161	307	162
rect	307	161	308	162
rect	308	161	309	162
rect	309	161	310	162
rect	310	161	311	162
rect	311	161	312	162
rect	312	161	313	162
rect	313	161	314	162
rect	314	161	315	162
rect	315	161	316	162
rect	316	161	317	162
rect	317	161	318	162
rect	318	161	319	162
rect	319	161	320	162
rect	320	161	321	162
rect	321	161	322	162
rect	322	161	323	162
rect	323	161	324	162
rect	324	161	325	162
rect	325	161	326	162
rect	326	161	327	162
rect	327	161	328	162
rect	328	161	329	162
rect	329	161	330	162
rect	330	161	331	162
rect	331	161	332	162
rect	332	161	333	162
rect	333	161	334	162
rect	334	161	335	162
rect	335	161	336	162
rect	336	161	337	162
rect	337	161	338	162
rect	339	161	340	162
rect	340	161	341	162
rect	341	161	342	162
rect	342	161	343	162
rect	343	161	344	162
rect	344	161	345	162
rect	345	161	346	162
rect	346	161	347	162
rect	347	161	348	162
rect	348	161	349	162
rect	349	161	350	162
rect	350	161	351	162
rect	351	161	352	162
rect	352	161	353	162
rect	353	161	354	162
rect	354	161	355	162
rect	355	161	356	162
rect	356	161	357	162
rect	357	161	358	162
rect	358	161	359	162
rect	359	161	360	162
rect	360	161	361	162
rect	361	161	362	162
rect	362	161	363	162
rect	363	161	364	162
rect	364	161	365	162
rect	365	161	366	162
rect	366	161	367	162
rect	367	161	368	162
rect	368	161	369	162
rect	369	161	370	162
rect	370	161	371	162
rect	371	161	372	162
rect	372	161	373	162
rect	373	161	374	162
rect	374	161	375	162
rect	375	161	376	162
rect	376	161	377	162
rect	377	161	378	162
rect	378	161	379	162
rect	379	161	380	162
rect	380	161	381	162
rect	381	161	382	162
rect	382	161	383	162
rect	383	161	384	162
rect	384	161	385	162
rect	385	161	386	162
rect	386	161	387	162
rect	387	161	388	162
rect	388	161	389	162
rect	389	161	390	162
rect	390	161	391	162
rect	391	161	392	162
rect	392	161	393	162
rect	393	161	394	162
rect	394	161	395	162
rect	395	161	396	162
rect	396	161	397	162
rect	397	161	398	162
rect	398	161	399	162
rect	399	161	400	162
rect	400	161	401	162
rect	401	161	402	162
rect	403	161	404	162
rect	404	161	405	162
rect	405	161	406	162
rect	406	161	407	162
rect	407	161	408	162
rect	408	161	409	162
rect	409	161	410	162
rect	410	161	411	162
rect	411	161	412	162
rect	412	161	413	162
rect	413	161	414	162
rect	414	161	415	162
rect	0	162	1	163
rect	1	162	2	163
rect	2	162	3	163
rect	3	162	4	163
rect	4	162	5	163
rect	5	162	6	163
rect	7	162	8	163
rect	8	162	9	163
rect	9	162	10	163
rect	10	162	11	163
rect	11	162	12	163
rect	12	162	13	163
rect	14	162	15	163
rect	15	162	16	163
rect	16	162	17	163
rect	17	162	18	163
rect	18	162	19	163
rect	19	162	20	163
rect	21	162	22	163
rect	22	162	23	163
rect	23	162	24	163
rect	24	162	25	163
rect	25	162	26	163
rect	26	162	27	163
rect	28	162	29	163
rect	29	162	30	163
rect	30	162	31	163
rect	31	162	32	163
rect	32	162	33	163
rect	33	162	34	163
rect	34	162	35	163
rect	35	162	36	163
rect	36	162	37	163
rect	37	162	38	163
rect	38	162	39	163
rect	39	162	40	163
rect	40	162	41	163
rect	41	162	42	163
rect	42	162	43	163
rect	43	162	44	163
rect	44	162	45	163
rect	45	162	46	163
rect	46	162	47	163
rect	47	162	48	163
rect	48	162	49	163
rect	49	162	50	163
rect	50	162	51	163
rect	51	162	52	163
rect	52	162	53	163
rect	53	162	54	163
rect	54	162	55	163
rect	55	162	56	163
rect	56	162	57	163
rect	57	162	58	163
rect	58	162	59	163
rect	59	162	60	163
rect	60	162	61	163
rect	61	162	62	163
rect	62	162	63	163
rect	63	162	64	163
rect	64	162	65	163
rect	65	162	66	163
rect	66	162	67	163
rect	67	162	68	163
rect	68	162	69	163
rect	69	162	70	163
rect	70	162	71	163
rect	71	162	72	163
rect	72	162	73	163
rect	74	162	75	163
rect	75	162	76	163
rect	76	162	77	163
rect	77	162	78	163
rect	78	162	79	163
rect	79	162	80	163
rect	81	162	82	163
rect	82	162	83	163
rect	83	162	84	163
rect	84	162	85	163
rect	85	162	86	163
rect	86	162	87	163
rect	88	162	89	163
rect	89	162	90	163
rect	90	162	91	163
rect	91	162	92	163
rect	92	162	93	163
rect	93	162	94	163
rect	94	162	95	163
rect	95	162	96	163
rect	96	162	97	163
rect	97	162	98	163
rect	98	162	99	163
rect	99	162	100	163
rect	100	162	101	163
rect	101	162	102	163
rect	102	162	103	163
rect	103	162	104	163
rect	104	162	105	163
rect	105	162	106	163
rect	106	162	107	163
rect	107	162	108	163
rect	108	162	109	163
rect	109	162	110	163
rect	110	162	111	163
rect	111	162	112	163
rect	112	162	113	163
rect	113	162	114	163
rect	114	162	115	163
rect	115	162	116	163
rect	116	162	117	163
rect	117	162	118	163
rect	118	162	119	163
rect	119	162	120	163
rect	120	162	121	163
rect	121	162	122	163
rect	122	162	123	163
rect	123	162	124	163
rect	124	162	125	163
rect	125	162	126	163
rect	126	162	127	163
rect	127	162	128	163
rect	128	162	129	163
rect	129	162	130	163
rect	130	162	131	163
rect	131	162	132	163
rect	132	162	133	163
rect	133	162	134	163
rect	134	162	135	163
rect	135	162	136	163
rect	136	162	137	163
rect	137	162	138	163
rect	138	162	139	163
rect	139	162	140	163
rect	140	162	141	163
rect	141	162	142	163
rect	142	162	143	163
rect	143	162	144	163
rect	144	162	145	163
rect	145	162	146	163
rect	146	162	147	163
rect	147	162	148	163
rect	148	162	149	163
rect	149	162	150	163
rect	150	162	151	163
rect	151	162	152	163
rect	152	162	153	163
rect	153	162	154	163
rect	154	162	155	163
rect	155	162	156	163
rect	156	162	157	163
rect	157	162	158	163
rect	158	162	159	163
rect	159	162	160	163
rect	160	162	161	163
rect	161	162	162	163
rect	162	162	163	163
rect	163	162	164	163
rect	164	162	165	163
rect	165	162	166	163
rect	166	162	167	163
rect	167	162	168	163
rect	168	162	169	163
rect	169	162	170	163
rect	170	162	171	163
rect	171	162	172	163
rect	172	162	173	163
rect	173	162	174	163
rect	174	162	175	163
rect	176	162	177	163
rect	177	162	178	163
rect	178	162	179	163
rect	179	162	180	163
rect	180	162	181	163
rect	181	162	182	163
rect	182	162	183	163
rect	183	162	184	163
rect	184	162	185	163
rect	185	162	186	163
rect	186	162	187	163
rect	187	162	188	163
rect	188	162	189	163
rect	189	162	190	163
rect	190	162	191	163
rect	191	162	192	163
rect	192	162	193	163
rect	193	162	194	163
rect	194	162	195	163
rect	195	162	196	163
rect	196	162	197	163
rect	197	162	198	163
rect	198	162	199	163
rect	199	162	200	163
rect	200	162	201	163
rect	201	162	202	163
rect	202	162	203	163
rect	203	162	204	163
rect	204	162	205	163
rect	205	162	206	163
rect	206	162	207	163
rect	207	162	208	163
rect	208	162	209	163
rect	209	162	210	163
rect	210	162	211	163
rect	211	162	212	163
rect	212	162	213	163
rect	213	162	214	163
rect	214	162	215	163
rect	215	162	216	163
rect	216	162	217	163
rect	217	162	218	163
rect	218	162	219	163
rect	219	162	220	163
rect	220	162	221	163
rect	221	162	222	163
rect	222	162	223	163
rect	223	162	224	163
rect	224	162	225	163
rect	225	162	226	163
rect	226	162	227	163
rect	227	162	228	163
rect	228	162	229	163
rect	229	162	230	163
rect	230	162	231	163
rect	231	162	232	163
rect	232	162	233	163
rect	233	162	234	163
rect	234	162	235	163
rect	235	162	236	163
rect	236	162	237	163
rect	237	162	238	163
rect	238	162	239	163
rect	239	162	240	163
rect	240	162	241	163
rect	241	162	242	163
rect	242	162	243	163
rect	243	162	244	163
rect	244	162	245	163
rect	245	162	246	163
rect	246	162	247	163
rect	247	162	248	163
rect	248	162	249	163
rect	249	162	250	163
rect	250	162	251	163
rect	251	162	252	163
rect	252	162	253	163
rect	253	162	254	163
rect	254	162	255	163
rect	255	162	256	163
rect	256	162	257	163
rect	257	162	258	163
rect	258	162	259	163
rect	259	162	260	163
rect	260	162	261	163
rect	261	162	262	163
rect	262	162	263	163
rect	263	162	264	163
rect	264	162	265	163
rect	265	162	266	163
rect	266	162	267	163
rect	267	162	268	163
rect	268	162	269	163
rect	269	162	270	163
rect	270	162	271	163
rect	271	162	272	163
rect	272	162	273	163
rect	273	162	274	163
rect	274	162	275	163
rect	275	162	276	163
rect	276	162	277	163
rect	277	162	278	163
rect	278	162	279	163
rect	279	162	280	163
rect	280	162	281	163
rect	281	162	282	163
rect	282	162	283	163
rect	283	162	284	163
rect	284	162	285	163
rect	285	162	286	163
rect	286	162	287	163
rect	287	162	288	163
rect	288	162	289	163
rect	289	162	290	163
rect	290	162	291	163
rect	291	162	292	163
rect	292	162	293	163
rect	293	162	294	163
rect	294	162	295	163
rect	295	162	296	163
rect	296	162	297	163
rect	297	162	298	163
rect	298	162	299	163
rect	299	162	300	163
rect	300	162	301	163
rect	301	162	302	163
rect	302	162	303	163
rect	303	162	304	163
rect	304	162	305	163
rect	305	162	306	163
rect	306	162	307	163
rect	307	162	308	163
rect	308	162	309	163
rect	309	162	310	163
rect	310	162	311	163
rect	311	162	312	163
rect	312	162	313	163
rect	313	162	314	163
rect	314	162	315	163
rect	315	162	316	163
rect	316	162	317	163
rect	317	162	318	163
rect	318	162	319	163
rect	319	162	320	163
rect	320	162	321	163
rect	321	162	322	163
rect	322	162	323	163
rect	323	162	324	163
rect	324	162	325	163
rect	325	162	326	163
rect	326	162	327	163
rect	327	162	328	163
rect	328	162	329	163
rect	329	162	330	163
rect	330	162	331	163
rect	331	162	332	163
rect	332	162	333	163
rect	333	162	334	163
rect	334	162	335	163
rect	335	162	336	163
rect	336	162	337	163
rect	337	162	338	163
rect	339	162	340	163
rect	340	162	341	163
rect	341	162	342	163
rect	342	162	343	163
rect	343	162	344	163
rect	344	162	345	163
rect	345	162	346	163
rect	346	162	347	163
rect	347	162	348	163
rect	348	162	349	163
rect	349	162	350	163
rect	350	162	351	163
rect	351	162	352	163
rect	352	162	353	163
rect	353	162	354	163
rect	354	162	355	163
rect	355	162	356	163
rect	356	162	357	163
rect	357	162	358	163
rect	358	162	359	163
rect	359	162	360	163
rect	360	162	361	163
rect	361	162	362	163
rect	362	162	363	163
rect	363	162	364	163
rect	364	162	365	163
rect	365	162	366	163
rect	366	162	367	163
rect	367	162	368	163
rect	368	162	369	163
rect	369	162	370	163
rect	370	162	371	163
rect	371	162	372	163
rect	372	162	373	163
rect	373	162	374	163
rect	374	162	375	163
rect	375	162	376	163
rect	376	162	377	163
rect	377	162	378	163
rect	378	162	379	163
rect	379	162	380	163
rect	380	162	381	163
rect	381	162	382	163
rect	382	162	383	163
rect	383	162	384	163
rect	384	162	385	163
rect	385	162	386	163
rect	386	162	387	163
rect	387	162	388	163
rect	388	162	389	163
rect	389	162	390	163
rect	390	162	391	163
rect	391	162	392	163
rect	392	162	393	163
rect	393	162	394	163
rect	394	162	395	163
rect	395	162	396	163
rect	396	162	397	163
rect	397	162	398	163
rect	398	162	399	163
rect	399	162	400	163
rect	400	162	401	163
rect	401	162	402	163
rect	403	162	404	163
rect	404	162	405	163
rect	405	162	406	163
rect	406	162	407	163
rect	407	162	408	163
rect	408	162	409	163
rect	409	162	410	163
rect	410	162	411	163
rect	411	162	412	163
rect	412	162	413	163
rect	413	162	414	163
rect	414	162	415	163
rect	0	186	1	187
rect	1	186	2	187
rect	2	186	3	187
rect	3	186	4	187
rect	4	186	5	187
rect	5	186	6	187
rect	7	186	8	187
rect	8	186	9	187
rect	9	186	10	187
rect	10	186	11	187
rect	11	186	12	187
rect	12	186	13	187
rect	13	186	14	187
rect	14	186	15	187
rect	15	186	16	187
rect	16	186	17	187
rect	17	186	18	187
rect	18	186	19	187
rect	19	186	20	187
rect	20	186	21	187
rect	21	186	22	187
rect	23	186	24	187
rect	24	186	25	187
rect	25	186	26	187
rect	26	186	27	187
rect	27	186	28	187
rect	28	186	29	187
rect	29	186	30	187
rect	30	186	31	187
rect	31	186	32	187
rect	32	186	33	187
rect	33	186	34	187
rect	34	186	35	187
rect	35	186	36	187
rect	36	186	37	187
rect	37	186	38	187
rect	38	186	39	187
rect	39	186	40	187
rect	40	186	41	187
rect	41	186	42	187
rect	42	186	43	187
rect	43	186	44	187
rect	44	186	45	187
rect	45	186	46	187
rect	46	186	47	187
rect	47	186	48	187
rect	48	186	49	187
rect	49	186	50	187
rect	50	186	51	187
rect	51	186	52	187
rect	52	186	53	187
rect	53	186	54	187
rect	54	186	55	187
rect	55	186	56	187
rect	56	186	57	187
rect	57	186	58	187
rect	58	186	59	187
rect	60	186	61	187
rect	61	186	62	187
rect	62	186	63	187
rect	63	186	64	187
rect	64	186	65	187
rect	65	186	66	187
rect	66	186	67	187
rect	67	186	68	187
rect	68	186	69	187
rect	69	186	70	187
rect	70	186	71	187
rect	71	186	72	187
rect	72	186	73	187
rect	73	186	74	187
rect	74	186	75	187
rect	76	186	77	187
rect	77	186	78	187
rect	78	186	79	187
rect	79	186	80	187
rect	80	186	81	187
rect	81	186	82	187
rect	83	186	84	187
rect	84	186	85	187
rect	85	186	86	187
rect	86	186	87	187
rect	87	186	88	187
rect	88	186	89	187
rect	90	186	91	187
rect	91	186	92	187
rect	92	186	93	187
rect	93	186	94	187
rect	94	186	95	187
rect	95	186	96	187
rect	96	186	97	187
rect	97	186	98	187
rect	98	186	99	187
rect	99	186	100	187
rect	100	186	101	187
rect	101	186	102	187
rect	102	186	103	187
rect	103	186	104	187
rect	104	186	105	187
rect	105	186	106	187
rect	106	186	107	187
rect	107	186	108	187
rect	109	186	110	187
rect	110	186	111	187
rect	111	186	112	187
rect	112	186	113	187
rect	113	186	114	187
rect	114	186	115	187
rect	115	186	116	187
rect	116	186	117	187
rect	117	186	118	187
rect	118	186	119	187
rect	119	186	120	187
rect	120	186	121	187
rect	121	186	122	187
rect	122	186	123	187
rect	123	186	124	187
rect	124	186	125	187
rect	125	186	126	187
rect	126	186	127	187
rect	127	186	128	187
rect	128	186	129	187
rect	129	186	130	187
rect	130	186	131	187
rect	131	186	132	187
rect	132	186	133	187
rect	133	186	134	187
rect	134	186	135	187
rect	135	186	136	187
rect	136	186	137	187
rect	137	186	138	187
rect	138	186	139	187
rect	139	186	140	187
rect	140	186	141	187
rect	141	186	142	187
rect	142	186	143	187
rect	143	186	144	187
rect	144	186	145	187
rect	145	186	146	187
rect	146	186	147	187
rect	147	186	148	187
rect	148	186	149	187
rect	149	186	150	187
rect	150	186	151	187
rect	151	186	152	187
rect	152	186	153	187
rect	153	186	154	187
rect	154	186	155	187
rect	155	186	156	187
rect	156	186	157	187
rect	157	186	158	187
rect	158	186	159	187
rect	159	186	160	187
rect	161	186	162	187
rect	162	186	163	187
rect	163	186	164	187
rect	164	186	165	187
rect	165	186	166	187
rect	166	186	167	187
rect	167	186	168	187
rect	168	186	169	187
rect	169	186	170	187
rect	170	186	171	187
rect	171	186	172	187
rect	172	186	173	187
rect	173	186	174	187
rect	174	186	175	187
rect	175	186	176	187
rect	176	186	177	187
rect	177	186	178	187
rect	178	186	179	187
rect	179	186	180	187
rect	180	186	181	187
rect	181	186	182	187
rect	182	186	183	187
rect	183	186	184	187
rect	184	186	185	187
rect	185	186	186	187
rect	186	186	187	187
rect	187	186	188	187
rect	188	186	189	187
rect	189	186	190	187
rect	190	186	191	187
rect	191	186	192	187
rect	192	186	193	187
rect	193	186	194	187
rect	195	186	196	187
rect	196	186	197	187
rect	197	186	198	187
rect	198	186	199	187
rect	199	186	200	187
rect	200	186	201	187
rect	201	186	202	187
rect	202	186	203	187
rect	203	186	204	187
rect	204	186	205	187
rect	205	186	206	187
rect	206	186	207	187
rect	207	186	208	187
rect	208	186	209	187
rect	209	186	210	187
rect	210	186	211	187
rect	211	186	212	187
rect	212	186	213	187
rect	213	186	214	187
rect	214	186	215	187
rect	215	186	216	187
rect	216	186	217	187
rect	217	186	218	187
rect	218	186	219	187
rect	219	186	220	187
rect	220	186	221	187
rect	221	186	222	187
rect	223	186	224	187
rect	224	186	225	187
rect	225	186	226	187
rect	226	186	227	187
rect	227	186	228	187
rect	228	186	229	187
rect	229	186	230	187
rect	230	186	231	187
rect	231	186	232	187
rect	232	186	233	187
rect	233	186	234	187
rect	234	186	235	187
rect	235	186	236	187
rect	236	186	237	187
rect	237	186	238	187
rect	238	186	239	187
rect	239	186	240	187
rect	240	186	241	187
rect	241	186	242	187
rect	242	186	243	187
rect	243	186	244	187
rect	244	186	245	187
rect	245	186	246	187
rect	246	186	247	187
rect	247	186	248	187
rect	248	186	249	187
rect	249	186	250	187
rect	250	186	251	187
rect	251	186	252	187
rect	252	186	253	187
rect	253	186	254	187
rect	254	186	255	187
rect	255	186	256	187
rect	256	186	257	187
rect	257	186	258	187
rect	258	186	259	187
rect	259	186	260	187
rect	260	186	261	187
rect	261	186	262	187
rect	262	186	263	187
rect	263	186	264	187
rect	264	186	265	187
rect	265	186	266	187
rect	266	186	267	187
rect	267	186	268	187
rect	268	186	269	187
rect	269	186	270	187
rect	270	186	271	187
rect	271	186	272	187
rect	272	186	273	187
rect	273	186	274	187
rect	274	186	275	187
rect	275	186	276	187
rect	276	186	277	187
rect	277	186	278	187
rect	278	186	279	187
rect	279	186	280	187
rect	280	186	281	187
rect	281	186	282	187
rect	282	186	283	187
rect	283	186	284	187
rect	284	186	285	187
rect	285	186	286	187
rect	286	186	287	187
rect	287	186	288	187
rect	288	186	289	187
rect	289	186	290	187
rect	290	186	291	187
rect	291	186	292	187
rect	292	186	293	187
rect	293	186	294	187
rect	294	186	295	187
rect	295	186	296	187
rect	296	186	297	187
rect	297	186	298	187
rect	298	186	299	187
rect	299	186	300	187
rect	300	186	301	187
rect	301	186	302	187
rect	302	186	303	187
rect	303	186	304	187
rect	304	186	305	187
rect	305	186	306	187
rect	306	186	307	187
rect	307	186	308	187
rect	308	186	309	187
rect	309	186	310	187
rect	310	186	311	187
rect	311	186	312	187
rect	312	186	313	187
rect	313	186	314	187
rect	314	186	315	187
rect	315	186	316	187
rect	316	186	317	187
rect	317	186	318	187
rect	318	186	319	187
rect	319	186	320	187
rect	320	186	321	187
rect	321	186	322	187
rect	322	186	323	187
rect	323	186	324	187
rect	324	186	325	187
rect	325	186	326	187
rect	326	186	327	187
rect	327	186	328	187
rect	328	186	329	187
rect	329	186	330	187
rect	330	186	331	187
rect	331	186	332	187
rect	332	186	333	187
rect	333	186	334	187
rect	334	186	335	187
rect	335	186	336	187
rect	336	186	337	187
rect	337	186	338	187
rect	338	186	339	187
rect	339	186	340	187
rect	340	186	341	187
rect	341	186	342	187
rect	342	186	343	187
rect	343	186	344	187
rect	344	186	345	187
rect	345	186	346	187
rect	346	186	347	187
rect	347	186	348	187
rect	348	186	349	187
rect	349	186	350	187
rect	350	186	351	187
rect	351	186	352	187
rect	352	186	353	187
rect	353	186	354	187
rect	354	186	355	187
rect	355	186	356	187
rect	356	186	357	187
rect	357	186	358	187
rect	358	186	359	187
rect	359	186	360	187
rect	360	186	361	187
rect	361	186	362	187
rect	362	186	363	187
rect	363	186	364	187
rect	364	186	365	187
rect	365	186	366	187
rect	366	186	367	187
rect	367	186	368	187
rect	368	186	369	187
rect	369	186	370	187
rect	370	186	371	187
rect	371	186	372	187
rect	372	186	373	187
rect	373	186	374	187
rect	374	186	375	187
rect	375	186	376	187
rect	377	186	378	187
rect	378	186	379	187
rect	379	186	380	187
rect	380	186	381	187
rect	381	186	382	187
rect	382	186	383	187
rect	384	186	385	187
rect	385	186	386	187
rect	386	186	387	187
rect	387	186	388	187
rect	388	186	389	187
rect	389	186	390	187
rect	390	186	391	187
rect	391	186	392	187
rect	392	186	393	187
rect	393	186	394	187
rect	394	186	395	187
rect	395	186	396	187
rect	396	186	397	187
rect	397	186	398	187
rect	398	186	399	187
rect	0	187	1	188
rect	1	187	2	188
rect	2	187	3	188
rect	3	187	4	188
rect	4	187	5	188
rect	5	187	6	188
rect	7	187	8	188
rect	8	187	9	188
rect	9	187	10	188
rect	10	187	11	188
rect	11	187	12	188
rect	12	187	13	188
rect	13	187	14	188
rect	14	187	15	188
rect	15	187	16	188
rect	16	187	17	188
rect	17	187	18	188
rect	18	187	19	188
rect	19	187	20	188
rect	20	187	21	188
rect	21	187	22	188
rect	23	187	24	188
rect	24	187	25	188
rect	25	187	26	188
rect	26	187	27	188
rect	27	187	28	188
rect	28	187	29	188
rect	29	187	30	188
rect	30	187	31	188
rect	31	187	32	188
rect	32	187	33	188
rect	33	187	34	188
rect	34	187	35	188
rect	35	187	36	188
rect	36	187	37	188
rect	37	187	38	188
rect	38	187	39	188
rect	39	187	40	188
rect	40	187	41	188
rect	41	187	42	188
rect	42	187	43	188
rect	43	187	44	188
rect	44	187	45	188
rect	45	187	46	188
rect	46	187	47	188
rect	47	187	48	188
rect	48	187	49	188
rect	49	187	50	188
rect	50	187	51	188
rect	51	187	52	188
rect	52	187	53	188
rect	53	187	54	188
rect	54	187	55	188
rect	55	187	56	188
rect	56	187	57	188
rect	57	187	58	188
rect	58	187	59	188
rect	60	187	61	188
rect	61	187	62	188
rect	62	187	63	188
rect	63	187	64	188
rect	64	187	65	188
rect	65	187	66	188
rect	66	187	67	188
rect	67	187	68	188
rect	68	187	69	188
rect	69	187	70	188
rect	70	187	71	188
rect	71	187	72	188
rect	72	187	73	188
rect	73	187	74	188
rect	74	187	75	188
rect	76	187	77	188
rect	77	187	78	188
rect	78	187	79	188
rect	79	187	80	188
rect	80	187	81	188
rect	81	187	82	188
rect	83	187	84	188
rect	84	187	85	188
rect	85	187	86	188
rect	86	187	87	188
rect	87	187	88	188
rect	88	187	89	188
rect	90	187	91	188
rect	91	187	92	188
rect	92	187	93	188
rect	93	187	94	188
rect	94	187	95	188
rect	95	187	96	188
rect	96	187	97	188
rect	97	187	98	188
rect	98	187	99	188
rect	99	187	100	188
rect	100	187	101	188
rect	101	187	102	188
rect	102	187	103	188
rect	103	187	104	188
rect	104	187	105	188
rect	105	187	106	188
rect	106	187	107	188
rect	107	187	108	188
rect	109	187	110	188
rect	110	187	111	188
rect	111	187	112	188
rect	112	187	113	188
rect	113	187	114	188
rect	114	187	115	188
rect	115	187	116	188
rect	116	187	117	188
rect	117	187	118	188
rect	118	187	119	188
rect	119	187	120	188
rect	120	187	121	188
rect	121	187	122	188
rect	122	187	123	188
rect	123	187	124	188
rect	124	187	125	188
rect	125	187	126	188
rect	126	187	127	188
rect	127	187	128	188
rect	128	187	129	188
rect	129	187	130	188
rect	130	187	131	188
rect	131	187	132	188
rect	132	187	133	188
rect	133	187	134	188
rect	134	187	135	188
rect	135	187	136	188
rect	136	187	137	188
rect	137	187	138	188
rect	138	187	139	188
rect	139	187	140	188
rect	140	187	141	188
rect	141	187	142	188
rect	142	187	143	188
rect	143	187	144	188
rect	144	187	145	188
rect	145	187	146	188
rect	146	187	147	188
rect	147	187	148	188
rect	148	187	149	188
rect	149	187	150	188
rect	150	187	151	188
rect	151	187	152	188
rect	152	187	153	188
rect	153	187	154	188
rect	154	187	155	188
rect	155	187	156	188
rect	156	187	157	188
rect	157	187	158	188
rect	158	187	159	188
rect	159	187	160	188
rect	161	187	162	188
rect	162	187	163	188
rect	163	187	164	188
rect	164	187	165	188
rect	165	187	166	188
rect	166	187	167	188
rect	167	187	168	188
rect	168	187	169	188
rect	169	187	170	188
rect	170	187	171	188
rect	171	187	172	188
rect	172	187	173	188
rect	173	187	174	188
rect	174	187	175	188
rect	175	187	176	188
rect	176	187	177	188
rect	177	187	178	188
rect	178	187	179	188
rect	179	187	180	188
rect	180	187	181	188
rect	181	187	182	188
rect	182	187	183	188
rect	183	187	184	188
rect	184	187	185	188
rect	185	187	186	188
rect	186	187	187	188
rect	187	187	188	188
rect	188	187	189	188
rect	189	187	190	188
rect	190	187	191	188
rect	191	187	192	188
rect	192	187	193	188
rect	193	187	194	188
rect	195	187	196	188
rect	196	187	197	188
rect	197	187	198	188
rect	198	187	199	188
rect	199	187	200	188
rect	200	187	201	188
rect	201	187	202	188
rect	202	187	203	188
rect	203	187	204	188
rect	204	187	205	188
rect	205	187	206	188
rect	206	187	207	188
rect	207	187	208	188
rect	208	187	209	188
rect	209	187	210	188
rect	210	187	211	188
rect	211	187	212	188
rect	212	187	213	188
rect	213	187	214	188
rect	214	187	215	188
rect	215	187	216	188
rect	216	187	217	188
rect	217	187	218	188
rect	218	187	219	188
rect	219	187	220	188
rect	220	187	221	188
rect	221	187	222	188
rect	223	187	224	188
rect	224	187	225	188
rect	225	187	226	188
rect	226	187	227	188
rect	227	187	228	188
rect	228	187	229	188
rect	229	187	230	188
rect	230	187	231	188
rect	231	187	232	188
rect	232	187	233	188
rect	233	187	234	188
rect	234	187	235	188
rect	235	187	236	188
rect	236	187	237	188
rect	237	187	238	188
rect	238	187	239	188
rect	239	187	240	188
rect	240	187	241	188
rect	241	187	242	188
rect	242	187	243	188
rect	243	187	244	188
rect	244	187	245	188
rect	245	187	246	188
rect	246	187	247	188
rect	247	187	248	188
rect	248	187	249	188
rect	249	187	250	188
rect	250	187	251	188
rect	251	187	252	188
rect	252	187	253	188
rect	253	187	254	188
rect	254	187	255	188
rect	255	187	256	188
rect	256	187	257	188
rect	257	187	258	188
rect	258	187	259	188
rect	259	187	260	188
rect	260	187	261	188
rect	261	187	262	188
rect	262	187	263	188
rect	263	187	264	188
rect	264	187	265	188
rect	265	187	266	188
rect	266	187	267	188
rect	267	187	268	188
rect	268	187	269	188
rect	269	187	270	188
rect	270	187	271	188
rect	271	187	272	188
rect	272	187	273	188
rect	273	187	274	188
rect	274	187	275	188
rect	275	187	276	188
rect	276	187	277	188
rect	277	187	278	188
rect	278	187	279	188
rect	279	187	280	188
rect	280	187	281	188
rect	281	187	282	188
rect	282	187	283	188
rect	283	187	284	188
rect	284	187	285	188
rect	285	187	286	188
rect	286	187	287	188
rect	287	187	288	188
rect	288	187	289	188
rect	289	187	290	188
rect	290	187	291	188
rect	291	187	292	188
rect	292	187	293	188
rect	293	187	294	188
rect	294	187	295	188
rect	295	187	296	188
rect	296	187	297	188
rect	297	187	298	188
rect	298	187	299	188
rect	299	187	300	188
rect	300	187	301	188
rect	301	187	302	188
rect	302	187	303	188
rect	303	187	304	188
rect	304	187	305	188
rect	305	187	306	188
rect	306	187	307	188
rect	307	187	308	188
rect	308	187	309	188
rect	309	187	310	188
rect	310	187	311	188
rect	311	187	312	188
rect	312	187	313	188
rect	313	187	314	188
rect	314	187	315	188
rect	315	187	316	188
rect	316	187	317	188
rect	317	187	318	188
rect	318	187	319	188
rect	319	187	320	188
rect	320	187	321	188
rect	321	187	322	188
rect	322	187	323	188
rect	323	187	324	188
rect	324	187	325	188
rect	325	187	326	188
rect	326	187	327	188
rect	327	187	328	188
rect	328	187	329	188
rect	329	187	330	188
rect	330	187	331	188
rect	331	187	332	188
rect	332	187	333	188
rect	333	187	334	188
rect	334	187	335	188
rect	335	187	336	188
rect	336	187	337	188
rect	337	187	338	188
rect	338	187	339	188
rect	339	187	340	188
rect	340	187	341	188
rect	341	187	342	188
rect	342	187	343	188
rect	343	187	344	188
rect	344	187	345	188
rect	345	187	346	188
rect	346	187	347	188
rect	347	187	348	188
rect	348	187	349	188
rect	349	187	350	188
rect	350	187	351	188
rect	351	187	352	188
rect	352	187	353	188
rect	353	187	354	188
rect	354	187	355	188
rect	355	187	356	188
rect	356	187	357	188
rect	357	187	358	188
rect	358	187	359	188
rect	359	187	360	188
rect	360	187	361	188
rect	361	187	362	188
rect	362	187	363	188
rect	363	187	364	188
rect	364	187	365	188
rect	365	187	366	188
rect	366	187	367	188
rect	367	187	368	188
rect	368	187	369	188
rect	369	187	370	188
rect	370	187	371	188
rect	371	187	372	188
rect	372	187	373	188
rect	373	187	374	188
rect	374	187	375	188
rect	375	187	376	188
rect	377	187	378	188
rect	378	187	379	188
rect	379	187	380	188
rect	380	187	381	188
rect	381	187	382	188
rect	382	187	383	188
rect	384	187	385	188
rect	385	187	386	188
rect	386	187	387	188
rect	387	187	388	188
rect	388	187	389	188
rect	389	187	390	188
rect	390	187	391	188
rect	391	187	392	188
rect	392	187	393	188
rect	393	187	394	188
rect	394	187	395	188
rect	395	187	396	188
rect	396	187	397	188
rect	397	187	398	188
rect	398	187	399	188
rect	0	188	1	189
rect	1	188	2	189
rect	2	188	3	189
rect	3	188	4	189
rect	4	188	5	189
rect	5	188	6	189
rect	7	188	8	189
rect	8	188	9	189
rect	9	188	10	189
rect	10	188	11	189
rect	11	188	12	189
rect	12	188	13	189
rect	13	188	14	189
rect	14	188	15	189
rect	15	188	16	189
rect	16	188	17	189
rect	17	188	18	189
rect	18	188	19	189
rect	19	188	20	189
rect	20	188	21	189
rect	21	188	22	189
rect	23	188	24	189
rect	24	188	25	189
rect	25	188	26	189
rect	26	188	27	189
rect	27	188	28	189
rect	28	188	29	189
rect	29	188	30	189
rect	30	188	31	189
rect	31	188	32	189
rect	32	188	33	189
rect	33	188	34	189
rect	34	188	35	189
rect	35	188	36	189
rect	36	188	37	189
rect	37	188	38	189
rect	38	188	39	189
rect	39	188	40	189
rect	40	188	41	189
rect	41	188	42	189
rect	42	188	43	189
rect	43	188	44	189
rect	44	188	45	189
rect	45	188	46	189
rect	46	188	47	189
rect	47	188	48	189
rect	48	188	49	189
rect	49	188	50	189
rect	50	188	51	189
rect	51	188	52	189
rect	52	188	53	189
rect	53	188	54	189
rect	54	188	55	189
rect	55	188	56	189
rect	56	188	57	189
rect	57	188	58	189
rect	58	188	59	189
rect	60	188	61	189
rect	61	188	62	189
rect	62	188	63	189
rect	63	188	64	189
rect	64	188	65	189
rect	65	188	66	189
rect	66	188	67	189
rect	67	188	68	189
rect	68	188	69	189
rect	69	188	70	189
rect	70	188	71	189
rect	71	188	72	189
rect	72	188	73	189
rect	73	188	74	189
rect	74	188	75	189
rect	76	188	77	189
rect	77	188	78	189
rect	78	188	79	189
rect	79	188	80	189
rect	80	188	81	189
rect	81	188	82	189
rect	83	188	84	189
rect	84	188	85	189
rect	85	188	86	189
rect	86	188	87	189
rect	87	188	88	189
rect	88	188	89	189
rect	90	188	91	189
rect	91	188	92	189
rect	92	188	93	189
rect	93	188	94	189
rect	94	188	95	189
rect	95	188	96	189
rect	96	188	97	189
rect	97	188	98	189
rect	98	188	99	189
rect	99	188	100	189
rect	100	188	101	189
rect	101	188	102	189
rect	102	188	103	189
rect	103	188	104	189
rect	104	188	105	189
rect	105	188	106	189
rect	106	188	107	189
rect	107	188	108	189
rect	109	188	110	189
rect	110	188	111	189
rect	111	188	112	189
rect	112	188	113	189
rect	113	188	114	189
rect	114	188	115	189
rect	115	188	116	189
rect	116	188	117	189
rect	117	188	118	189
rect	118	188	119	189
rect	119	188	120	189
rect	120	188	121	189
rect	121	188	122	189
rect	122	188	123	189
rect	123	188	124	189
rect	124	188	125	189
rect	125	188	126	189
rect	126	188	127	189
rect	127	188	128	189
rect	128	188	129	189
rect	129	188	130	189
rect	130	188	131	189
rect	131	188	132	189
rect	132	188	133	189
rect	133	188	134	189
rect	134	188	135	189
rect	135	188	136	189
rect	136	188	137	189
rect	137	188	138	189
rect	138	188	139	189
rect	139	188	140	189
rect	140	188	141	189
rect	141	188	142	189
rect	142	188	143	189
rect	143	188	144	189
rect	144	188	145	189
rect	145	188	146	189
rect	146	188	147	189
rect	147	188	148	189
rect	148	188	149	189
rect	149	188	150	189
rect	150	188	151	189
rect	151	188	152	189
rect	152	188	153	189
rect	153	188	154	189
rect	154	188	155	189
rect	155	188	156	189
rect	156	188	157	189
rect	157	188	158	189
rect	158	188	159	189
rect	159	188	160	189
rect	161	188	162	189
rect	162	188	163	189
rect	163	188	164	189
rect	164	188	165	189
rect	165	188	166	189
rect	166	188	167	189
rect	167	188	168	189
rect	168	188	169	189
rect	169	188	170	189
rect	170	188	171	189
rect	171	188	172	189
rect	172	188	173	189
rect	173	188	174	189
rect	174	188	175	189
rect	175	188	176	189
rect	176	188	177	189
rect	177	188	178	189
rect	178	188	179	189
rect	179	188	180	189
rect	180	188	181	189
rect	181	188	182	189
rect	182	188	183	189
rect	183	188	184	189
rect	184	188	185	189
rect	185	188	186	189
rect	186	188	187	189
rect	187	188	188	189
rect	188	188	189	189
rect	189	188	190	189
rect	190	188	191	189
rect	191	188	192	189
rect	192	188	193	189
rect	193	188	194	189
rect	195	188	196	189
rect	196	188	197	189
rect	197	188	198	189
rect	198	188	199	189
rect	199	188	200	189
rect	200	188	201	189
rect	201	188	202	189
rect	202	188	203	189
rect	203	188	204	189
rect	204	188	205	189
rect	205	188	206	189
rect	206	188	207	189
rect	207	188	208	189
rect	208	188	209	189
rect	209	188	210	189
rect	210	188	211	189
rect	211	188	212	189
rect	212	188	213	189
rect	213	188	214	189
rect	214	188	215	189
rect	215	188	216	189
rect	216	188	217	189
rect	217	188	218	189
rect	218	188	219	189
rect	219	188	220	189
rect	220	188	221	189
rect	221	188	222	189
rect	223	188	224	189
rect	224	188	225	189
rect	225	188	226	189
rect	226	188	227	189
rect	227	188	228	189
rect	228	188	229	189
rect	229	188	230	189
rect	230	188	231	189
rect	231	188	232	189
rect	232	188	233	189
rect	233	188	234	189
rect	234	188	235	189
rect	235	188	236	189
rect	236	188	237	189
rect	237	188	238	189
rect	238	188	239	189
rect	239	188	240	189
rect	240	188	241	189
rect	241	188	242	189
rect	242	188	243	189
rect	243	188	244	189
rect	244	188	245	189
rect	245	188	246	189
rect	246	188	247	189
rect	247	188	248	189
rect	248	188	249	189
rect	249	188	250	189
rect	250	188	251	189
rect	251	188	252	189
rect	252	188	253	189
rect	253	188	254	189
rect	254	188	255	189
rect	255	188	256	189
rect	256	188	257	189
rect	257	188	258	189
rect	258	188	259	189
rect	259	188	260	189
rect	260	188	261	189
rect	261	188	262	189
rect	262	188	263	189
rect	263	188	264	189
rect	264	188	265	189
rect	265	188	266	189
rect	266	188	267	189
rect	267	188	268	189
rect	268	188	269	189
rect	269	188	270	189
rect	270	188	271	189
rect	271	188	272	189
rect	272	188	273	189
rect	273	188	274	189
rect	274	188	275	189
rect	275	188	276	189
rect	276	188	277	189
rect	277	188	278	189
rect	278	188	279	189
rect	279	188	280	189
rect	280	188	281	189
rect	281	188	282	189
rect	282	188	283	189
rect	283	188	284	189
rect	284	188	285	189
rect	285	188	286	189
rect	286	188	287	189
rect	287	188	288	189
rect	288	188	289	189
rect	289	188	290	189
rect	290	188	291	189
rect	291	188	292	189
rect	292	188	293	189
rect	293	188	294	189
rect	294	188	295	189
rect	295	188	296	189
rect	296	188	297	189
rect	297	188	298	189
rect	298	188	299	189
rect	299	188	300	189
rect	300	188	301	189
rect	301	188	302	189
rect	302	188	303	189
rect	303	188	304	189
rect	304	188	305	189
rect	305	188	306	189
rect	306	188	307	189
rect	307	188	308	189
rect	308	188	309	189
rect	309	188	310	189
rect	310	188	311	189
rect	311	188	312	189
rect	312	188	313	189
rect	313	188	314	189
rect	314	188	315	189
rect	315	188	316	189
rect	316	188	317	189
rect	317	188	318	189
rect	318	188	319	189
rect	319	188	320	189
rect	320	188	321	189
rect	321	188	322	189
rect	322	188	323	189
rect	323	188	324	189
rect	324	188	325	189
rect	325	188	326	189
rect	326	188	327	189
rect	327	188	328	189
rect	328	188	329	189
rect	329	188	330	189
rect	330	188	331	189
rect	331	188	332	189
rect	332	188	333	189
rect	333	188	334	189
rect	334	188	335	189
rect	335	188	336	189
rect	336	188	337	189
rect	337	188	338	189
rect	338	188	339	189
rect	339	188	340	189
rect	340	188	341	189
rect	341	188	342	189
rect	342	188	343	189
rect	343	188	344	189
rect	344	188	345	189
rect	345	188	346	189
rect	346	188	347	189
rect	347	188	348	189
rect	348	188	349	189
rect	349	188	350	189
rect	350	188	351	189
rect	351	188	352	189
rect	352	188	353	189
rect	353	188	354	189
rect	354	188	355	189
rect	355	188	356	189
rect	356	188	357	189
rect	357	188	358	189
rect	358	188	359	189
rect	359	188	360	189
rect	360	188	361	189
rect	361	188	362	189
rect	362	188	363	189
rect	363	188	364	189
rect	364	188	365	189
rect	365	188	366	189
rect	366	188	367	189
rect	367	188	368	189
rect	368	188	369	189
rect	369	188	370	189
rect	370	188	371	189
rect	371	188	372	189
rect	372	188	373	189
rect	373	188	374	189
rect	374	188	375	189
rect	375	188	376	189
rect	377	188	378	189
rect	378	188	379	189
rect	379	188	380	189
rect	380	188	381	189
rect	381	188	382	189
rect	382	188	383	189
rect	384	188	385	189
rect	385	188	386	189
rect	386	188	387	189
rect	387	188	388	189
rect	388	188	389	189
rect	389	188	390	189
rect	390	188	391	189
rect	391	188	392	189
rect	392	188	393	189
rect	393	188	394	189
rect	394	188	395	189
rect	395	188	396	189
rect	396	188	397	189
rect	397	188	398	189
rect	398	188	399	189
rect	0	189	1	190
rect	1	189	2	190
rect	2	189	3	190
rect	3	189	4	190
rect	4	189	5	190
rect	5	189	6	190
rect	7	189	8	190
rect	8	189	9	190
rect	9	189	10	190
rect	10	189	11	190
rect	11	189	12	190
rect	12	189	13	190
rect	13	189	14	190
rect	14	189	15	190
rect	15	189	16	190
rect	16	189	17	190
rect	17	189	18	190
rect	18	189	19	190
rect	19	189	20	190
rect	20	189	21	190
rect	21	189	22	190
rect	23	189	24	190
rect	24	189	25	190
rect	25	189	26	190
rect	26	189	27	190
rect	27	189	28	190
rect	28	189	29	190
rect	29	189	30	190
rect	30	189	31	190
rect	31	189	32	190
rect	32	189	33	190
rect	33	189	34	190
rect	34	189	35	190
rect	35	189	36	190
rect	36	189	37	190
rect	37	189	38	190
rect	38	189	39	190
rect	39	189	40	190
rect	40	189	41	190
rect	41	189	42	190
rect	42	189	43	190
rect	43	189	44	190
rect	44	189	45	190
rect	45	189	46	190
rect	46	189	47	190
rect	47	189	48	190
rect	48	189	49	190
rect	49	189	50	190
rect	50	189	51	190
rect	51	189	52	190
rect	52	189	53	190
rect	53	189	54	190
rect	54	189	55	190
rect	55	189	56	190
rect	56	189	57	190
rect	57	189	58	190
rect	58	189	59	190
rect	60	189	61	190
rect	61	189	62	190
rect	62	189	63	190
rect	63	189	64	190
rect	64	189	65	190
rect	65	189	66	190
rect	66	189	67	190
rect	67	189	68	190
rect	68	189	69	190
rect	69	189	70	190
rect	70	189	71	190
rect	71	189	72	190
rect	72	189	73	190
rect	73	189	74	190
rect	74	189	75	190
rect	76	189	77	190
rect	77	189	78	190
rect	78	189	79	190
rect	79	189	80	190
rect	80	189	81	190
rect	81	189	82	190
rect	83	189	84	190
rect	84	189	85	190
rect	85	189	86	190
rect	86	189	87	190
rect	87	189	88	190
rect	88	189	89	190
rect	90	189	91	190
rect	91	189	92	190
rect	92	189	93	190
rect	93	189	94	190
rect	94	189	95	190
rect	95	189	96	190
rect	96	189	97	190
rect	97	189	98	190
rect	98	189	99	190
rect	99	189	100	190
rect	100	189	101	190
rect	101	189	102	190
rect	102	189	103	190
rect	103	189	104	190
rect	104	189	105	190
rect	105	189	106	190
rect	106	189	107	190
rect	107	189	108	190
rect	109	189	110	190
rect	110	189	111	190
rect	111	189	112	190
rect	112	189	113	190
rect	113	189	114	190
rect	114	189	115	190
rect	115	189	116	190
rect	116	189	117	190
rect	117	189	118	190
rect	118	189	119	190
rect	119	189	120	190
rect	120	189	121	190
rect	121	189	122	190
rect	122	189	123	190
rect	123	189	124	190
rect	124	189	125	190
rect	125	189	126	190
rect	126	189	127	190
rect	127	189	128	190
rect	128	189	129	190
rect	129	189	130	190
rect	130	189	131	190
rect	131	189	132	190
rect	132	189	133	190
rect	133	189	134	190
rect	134	189	135	190
rect	135	189	136	190
rect	136	189	137	190
rect	137	189	138	190
rect	138	189	139	190
rect	139	189	140	190
rect	140	189	141	190
rect	141	189	142	190
rect	142	189	143	190
rect	143	189	144	190
rect	144	189	145	190
rect	145	189	146	190
rect	146	189	147	190
rect	147	189	148	190
rect	148	189	149	190
rect	149	189	150	190
rect	150	189	151	190
rect	151	189	152	190
rect	152	189	153	190
rect	153	189	154	190
rect	154	189	155	190
rect	155	189	156	190
rect	156	189	157	190
rect	157	189	158	190
rect	158	189	159	190
rect	159	189	160	190
rect	161	189	162	190
rect	162	189	163	190
rect	163	189	164	190
rect	164	189	165	190
rect	165	189	166	190
rect	166	189	167	190
rect	167	189	168	190
rect	168	189	169	190
rect	169	189	170	190
rect	170	189	171	190
rect	171	189	172	190
rect	172	189	173	190
rect	173	189	174	190
rect	174	189	175	190
rect	175	189	176	190
rect	176	189	177	190
rect	177	189	178	190
rect	178	189	179	190
rect	179	189	180	190
rect	180	189	181	190
rect	181	189	182	190
rect	182	189	183	190
rect	183	189	184	190
rect	184	189	185	190
rect	185	189	186	190
rect	186	189	187	190
rect	187	189	188	190
rect	188	189	189	190
rect	189	189	190	190
rect	190	189	191	190
rect	191	189	192	190
rect	192	189	193	190
rect	193	189	194	190
rect	195	189	196	190
rect	196	189	197	190
rect	197	189	198	190
rect	198	189	199	190
rect	199	189	200	190
rect	200	189	201	190
rect	201	189	202	190
rect	202	189	203	190
rect	203	189	204	190
rect	204	189	205	190
rect	205	189	206	190
rect	206	189	207	190
rect	207	189	208	190
rect	208	189	209	190
rect	209	189	210	190
rect	210	189	211	190
rect	211	189	212	190
rect	212	189	213	190
rect	213	189	214	190
rect	214	189	215	190
rect	215	189	216	190
rect	216	189	217	190
rect	217	189	218	190
rect	218	189	219	190
rect	219	189	220	190
rect	220	189	221	190
rect	221	189	222	190
rect	223	189	224	190
rect	224	189	225	190
rect	225	189	226	190
rect	226	189	227	190
rect	227	189	228	190
rect	228	189	229	190
rect	229	189	230	190
rect	230	189	231	190
rect	231	189	232	190
rect	232	189	233	190
rect	233	189	234	190
rect	234	189	235	190
rect	235	189	236	190
rect	236	189	237	190
rect	237	189	238	190
rect	238	189	239	190
rect	239	189	240	190
rect	240	189	241	190
rect	241	189	242	190
rect	242	189	243	190
rect	243	189	244	190
rect	244	189	245	190
rect	245	189	246	190
rect	246	189	247	190
rect	247	189	248	190
rect	248	189	249	190
rect	249	189	250	190
rect	250	189	251	190
rect	251	189	252	190
rect	252	189	253	190
rect	253	189	254	190
rect	254	189	255	190
rect	255	189	256	190
rect	256	189	257	190
rect	257	189	258	190
rect	258	189	259	190
rect	259	189	260	190
rect	260	189	261	190
rect	261	189	262	190
rect	262	189	263	190
rect	263	189	264	190
rect	264	189	265	190
rect	265	189	266	190
rect	266	189	267	190
rect	267	189	268	190
rect	268	189	269	190
rect	269	189	270	190
rect	270	189	271	190
rect	271	189	272	190
rect	272	189	273	190
rect	273	189	274	190
rect	274	189	275	190
rect	275	189	276	190
rect	276	189	277	190
rect	277	189	278	190
rect	278	189	279	190
rect	279	189	280	190
rect	280	189	281	190
rect	281	189	282	190
rect	282	189	283	190
rect	283	189	284	190
rect	284	189	285	190
rect	285	189	286	190
rect	286	189	287	190
rect	287	189	288	190
rect	288	189	289	190
rect	289	189	290	190
rect	290	189	291	190
rect	291	189	292	190
rect	292	189	293	190
rect	293	189	294	190
rect	294	189	295	190
rect	295	189	296	190
rect	296	189	297	190
rect	297	189	298	190
rect	298	189	299	190
rect	299	189	300	190
rect	300	189	301	190
rect	301	189	302	190
rect	302	189	303	190
rect	303	189	304	190
rect	304	189	305	190
rect	305	189	306	190
rect	306	189	307	190
rect	307	189	308	190
rect	308	189	309	190
rect	309	189	310	190
rect	310	189	311	190
rect	311	189	312	190
rect	312	189	313	190
rect	313	189	314	190
rect	314	189	315	190
rect	315	189	316	190
rect	316	189	317	190
rect	317	189	318	190
rect	318	189	319	190
rect	319	189	320	190
rect	320	189	321	190
rect	321	189	322	190
rect	322	189	323	190
rect	323	189	324	190
rect	324	189	325	190
rect	325	189	326	190
rect	326	189	327	190
rect	327	189	328	190
rect	328	189	329	190
rect	329	189	330	190
rect	330	189	331	190
rect	331	189	332	190
rect	332	189	333	190
rect	333	189	334	190
rect	334	189	335	190
rect	335	189	336	190
rect	336	189	337	190
rect	337	189	338	190
rect	338	189	339	190
rect	339	189	340	190
rect	340	189	341	190
rect	341	189	342	190
rect	342	189	343	190
rect	343	189	344	190
rect	344	189	345	190
rect	345	189	346	190
rect	346	189	347	190
rect	347	189	348	190
rect	348	189	349	190
rect	349	189	350	190
rect	350	189	351	190
rect	351	189	352	190
rect	352	189	353	190
rect	353	189	354	190
rect	354	189	355	190
rect	355	189	356	190
rect	356	189	357	190
rect	357	189	358	190
rect	358	189	359	190
rect	359	189	360	190
rect	360	189	361	190
rect	361	189	362	190
rect	362	189	363	190
rect	363	189	364	190
rect	364	189	365	190
rect	365	189	366	190
rect	366	189	367	190
rect	367	189	368	190
rect	368	189	369	190
rect	369	189	370	190
rect	370	189	371	190
rect	371	189	372	190
rect	372	189	373	190
rect	373	189	374	190
rect	374	189	375	190
rect	375	189	376	190
rect	377	189	378	190
rect	378	189	379	190
rect	379	189	380	190
rect	380	189	381	190
rect	381	189	382	190
rect	382	189	383	190
rect	384	189	385	190
rect	385	189	386	190
rect	386	189	387	190
rect	387	189	388	190
rect	388	189	389	190
rect	389	189	390	190
rect	390	189	391	190
rect	391	189	392	190
rect	392	189	393	190
rect	393	189	394	190
rect	394	189	395	190
rect	395	189	396	190
rect	396	189	397	190
rect	397	189	398	190
rect	398	189	399	190
rect	0	190	1	191
rect	1	190	2	191
rect	2	190	3	191
rect	3	190	4	191
rect	4	190	5	191
rect	5	190	6	191
rect	7	190	8	191
rect	8	190	9	191
rect	9	190	10	191
rect	10	190	11	191
rect	11	190	12	191
rect	12	190	13	191
rect	13	190	14	191
rect	14	190	15	191
rect	15	190	16	191
rect	16	190	17	191
rect	17	190	18	191
rect	18	190	19	191
rect	19	190	20	191
rect	20	190	21	191
rect	21	190	22	191
rect	23	190	24	191
rect	24	190	25	191
rect	25	190	26	191
rect	26	190	27	191
rect	27	190	28	191
rect	28	190	29	191
rect	29	190	30	191
rect	30	190	31	191
rect	31	190	32	191
rect	32	190	33	191
rect	33	190	34	191
rect	34	190	35	191
rect	35	190	36	191
rect	36	190	37	191
rect	37	190	38	191
rect	38	190	39	191
rect	39	190	40	191
rect	40	190	41	191
rect	41	190	42	191
rect	42	190	43	191
rect	43	190	44	191
rect	44	190	45	191
rect	45	190	46	191
rect	46	190	47	191
rect	47	190	48	191
rect	48	190	49	191
rect	49	190	50	191
rect	50	190	51	191
rect	51	190	52	191
rect	52	190	53	191
rect	53	190	54	191
rect	54	190	55	191
rect	55	190	56	191
rect	56	190	57	191
rect	57	190	58	191
rect	58	190	59	191
rect	60	190	61	191
rect	61	190	62	191
rect	62	190	63	191
rect	63	190	64	191
rect	64	190	65	191
rect	65	190	66	191
rect	66	190	67	191
rect	67	190	68	191
rect	68	190	69	191
rect	69	190	70	191
rect	70	190	71	191
rect	71	190	72	191
rect	72	190	73	191
rect	73	190	74	191
rect	74	190	75	191
rect	76	190	77	191
rect	77	190	78	191
rect	78	190	79	191
rect	79	190	80	191
rect	80	190	81	191
rect	81	190	82	191
rect	83	190	84	191
rect	84	190	85	191
rect	85	190	86	191
rect	86	190	87	191
rect	87	190	88	191
rect	88	190	89	191
rect	90	190	91	191
rect	91	190	92	191
rect	92	190	93	191
rect	93	190	94	191
rect	94	190	95	191
rect	95	190	96	191
rect	96	190	97	191
rect	97	190	98	191
rect	98	190	99	191
rect	99	190	100	191
rect	100	190	101	191
rect	101	190	102	191
rect	102	190	103	191
rect	103	190	104	191
rect	104	190	105	191
rect	105	190	106	191
rect	106	190	107	191
rect	107	190	108	191
rect	109	190	110	191
rect	110	190	111	191
rect	111	190	112	191
rect	112	190	113	191
rect	113	190	114	191
rect	114	190	115	191
rect	115	190	116	191
rect	116	190	117	191
rect	117	190	118	191
rect	118	190	119	191
rect	119	190	120	191
rect	120	190	121	191
rect	121	190	122	191
rect	122	190	123	191
rect	123	190	124	191
rect	124	190	125	191
rect	125	190	126	191
rect	126	190	127	191
rect	127	190	128	191
rect	128	190	129	191
rect	129	190	130	191
rect	130	190	131	191
rect	131	190	132	191
rect	132	190	133	191
rect	133	190	134	191
rect	134	190	135	191
rect	135	190	136	191
rect	136	190	137	191
rect	137	190	138	191
rect	138	190	139	191
rect	139	190	140	191
rect	140	190	141	191
rect	141	190	142	191
rect	142	190	143	191
rect	143	190	144	191
rect	144	190	145	191
rect	145	190	146	191
rect	146	190	147	191
rect	147	190	148	191
rect	148	190	149	191
rect	149	190	150	191
rect	150	190	151	191
rect	151	190	152	191
rect	152	190	153	191
rect	153	190	154	191
rect	154	190	155	191
rect	155	190	156	191
rect	156	190	157	191
rect	157	190	158	191
rect	158	190	159	191
rect	159	190	160	191
rect	161	190	162	191
rect	162	190	163	191
rect	163	190	164	191
rect	164	190	165	191
rect	165	190	166	191
rect	166	190	167	191
rect	167	190	168	191
rect	168	190	169	191
rect	169	190	170	191
rect	170	190	171	191
rect	171	190	172	191
rect	172	190	173	191
rect	173	190	174	191
rect	174	190	175	191
rect	175	190	176	191
rect	176	190	177	191
rect	177	190	178	191
rect	178	190	179	191
rect	179	190	180	191
rect	180	190	181	191
rect	181	190	182	191
rect	182	190	183	191
rect	183	190	184	191
rect	184	190	185	191
rect	185	190	186	191
rect	186	190	187	191
rect	187	190	188	191
rect	188	190	189	191
rect	189	190	190	191
rect	190	190	191	191
rect	191	190	192	191
rect	192	190	193	191
rect	193	190	194	191
rect	195	190	196	191
rect	196	190	197	191
rect	197	190	198	191
rect	198	190	199	191
rect	199	190	200	191
rect	200	190	201	191
rect	201	190	202	191
rect	202	190	203	191
rect	203	190	204	191
rect	204	190	205	191
rect	205	190	206	191
rect	206	190	207	191
rect	207	190	208	191
rect	208	190	209	191
rect	209	190	210	191
rect	210	190	211	191
rect	211	190	212	191
rect	212	190	213	191
rect	213	190	214	191
rect	214	190	215	191
rect	215	190	216	191
rect	216	190	217	191
rect	217	190	218	191
rect	218	190	219	191
rect	219	190	220	191
rect	220	190	221	191
rect	221	190	222	191
rect	223	190	224	191
rect	224	190	225	191
rect	225	190	226	191
rect	226	190	227	191
rect	227	190	228	191
rect	228	190	229	191
rect	229	190	230	191
rect	230	190	231	191
rect	231	190	232	191
rect	232	190	233	191
rect	233	190	234	191
rect	234	190	235	191
rect	235	190	236	191
rect	236	190	237	191
rect	237	190	238	191
rect	238	190	239	191
rect	239	190	240	191
rect	240	190	241	191
rect	241	190	242	191
rect	242	190	243	191
rect	243	190	244	191
rect	244	190	245	191
rect	245	190	246	191
rect	246	190	247	191
rect	247	190	248	191
rect	248	190	249	191
rect	249	190	250	191
rect	250	190	251	191
rect	251	190	252	191
rect	252	190	253	191
rect	253	190	254	191
rect	254	190	255	191
rect	255	190	256	191
rect	256	190	257	191
rect	257	190	258	191
rect	258	190	259	191
rect	259	190	260	191
rect	260	190	261	191
rect	261	190	262	191
rect	262	190	263	191
rect	263	190	264	191
rect	264	190	265	191
rect	265	190	266	191
rect	266	190	267	191
rect	267	190	268	191
rect	268	190	269	191
rect	269	190	270	191
rect	270	190	271	191
rect	271	190	272	191
rect	272	190	273	191
rect	273	190	274	191
rect	274	190	275	191
rect	275	190	276	191
rect	276	190	277	191
rect	277	190	278	191
rect	278	190	279	191
rect	279	190	280	191
rect	280	190	281	191
rect	281	190	282	191
rect	282	190	283	191
rect	283	190	284	191
rect	284	190	285	191
rect	285	190	286	191
rect	286	190	287	191
rect	287	190	288	191
rect	288	190	289	191
rect	289	190	290	191
rect	290	190	291	191
rect	291	190	292	191
rect	292	190	293	191
rect	293	190	294	191
rect	294	190	295	191
rect	295	190	296	191
rect	296	190	297	191
rect	297	190	298	191
rect	298	190	299	191
rect	299	190	300	191
rect	300	190	301	191
rect	301	190	302	191
rect	302	190	303	191
rect	303	190	304	191
rect	304	190	305	191
rect	305	190	306	191
rect	306	190	307	191
rect	307	190	308	191
rect	308	190	309	191
rect	309	190	310	191
rect	310	190	311	191
rect	311	190	312	191
rect	312	190	313	191
rect	313	190	314	191
rect	314	190	315	191
rect	315	190	316	191
rect	316	190	317	191
rect	317	190	318	191
rect	318	190	319	191
rect	319	190	320	191
rect	320	190	321	191
rect	321	190	322	191
rect	322	190	323	191
rect	323	190	324	191
rect	324	190	325	191
rect	325	190	326	191
rect	326	190	327	191
rect	327	190	328	191
rect	328	190	329	191
rect	329	190	330	191
rect	330	190	331	191
rect	331	190	332	191
rect	332	190	333	191
rect	333	190	334	191
rect	334	190	335	191
rect	335	190	336	191
rect	336	190	337	191
rect	337	190	338	191
rect	338	190	339	191
rect	339	190	340	191
rect	340	190	341	191
rect	341	190	342	191
rect	342	190	343	191
rect	343	190	344	191
rect	344	190	345	191
rect	345	190	346	191
rect	346	190	347	191
rect	347	190	348	191
rect	348	190	349	191
rect	349	190	350	191
rect	350	190	351	191
rect	351	190	352	191
rect	352	190	353	191
rect	353	190	354	191
rect	354	190	355	191
rect	355	190	356	191
rect	356	190	357	191
rect	357	190	358	191
rect	358	190	359	191
rect	359	190	360	191
rect	360	190	361	191
rect	361	190	362	191
rect	362	190	363	191
rect	363	190	364	191
rect	364	190	365	191
rect	365	190	366	191
rect	366	190	367	191
rect	367	190	368	191
rect	368	190	369	191
rect	369	190	370	191
rect	370	190	371	191
rect	371	190	372	191
rect	372	190	373	191
rect	373	190	374	191
rect	374	190	375	191
rect	375	190	376	191
rect	377	190	378	191
rect	378	190	379	191
rect	379	190	380	191
rect	380	190	381	191
rect	381	190	382	191
rect	382	190	383	191
rect	384	190	385	191
rect	385	190	386	191
rect	386	190	387	191
rect	387	190	388	191
rect	388	190	389	191
rect	389	190	390	191
rect	390	190	391	191
rect	391	190	392	191
rect	392	190	393	191
rect	393	190	394	191
rect	394	190	395	191
rect	395	190	396	191
rect	396	190	397	191
rect	397	190	398	191
rect	398	190	399	191
rect	0	191	1	192
rect	1	191	2	192
rect	2	191	3	192
rect	3	191	4	192
rect	4	191	5	192
rect	5	191	6	192
rect	7	191	8	192
rect	8	191	9	192
rect	9	191	10	192
rect	10	191	11	192
rect	11	191	12	192
rect	12	191	13	192
rect	13	191	14	192
rect	14	191	15	192
rect	15	191	16	192
rect	16	191	17	192
rect	17	191	18	192
rect	18	191	19	192
rect	19	191	20	192
rect	20	191	21	192
rect	21	191	22	192
rect	23	191	24	192
rect	24	191	25	192
rect	25	191	26	192
rect	26	191	27	192
rect	27	191	28	192
rect	28	191	29	192
rect	29	191	30	192
rect	30	191	31	192
rect	31	191	32	192
rect	32	191	33	192
rect	33	191	34	192
rect	34	191	35	192
rect	35	191	36	192
rect	36	191	37	192
rect	37	191	38	192
rect	38	191	39	192
rect	39	191	40	192
rect	40	191	41	192
rect	41	191	42	192
rect	42	191	43	192
rect	43	191	44	192
rect	44	191	45	192
rect	45	191	46	192
rect	46	191	47	192
rect	47	191	48	192
rect	48	191	49	192
rect	49	191	50	192
rect	50	191	51	192
rect	51	191	52	192
rect	52	191	53	192
rect	53	191	54	192
rect	54	191	55	192
rect	55	191	56	192
rect	56	191	57	192
rect	57	191	58	192
rect	58	191	59	192
rect	60	191	61	192
rect	61	191	62	192
rect	62	191	63	192
rect	63	191	64	192
rect	64	191	65	192
rect	65	191	66	192
rect	66	191	67	192
rect	67	191	68	192
rect	68	191	69	192
rect	69	191	70	192
rect	70	191	71	192
rect	71	191	72	192
rect	72	191	73	192
rect	73	191	74	192
rect	74	191	75	192
rect	76	191	77	192
rect	77	191	78	192
rect	78	191	79	192
rect	79	191	80	192
rect	80	191	81	192
rect	81	191	82	192
rect	83	191	84	192
rect	84	191	85	192
rect	85	191	86	192
rect	86	191	87	192
rect	87	191	88	192
rect	88	191	89	192
rect	90	191	91	192
rect	91	191	92	192
rect	92	191	93	192
rect	93	191	94	192
rect	94	191	95	192
rect	95	191	96	192
rect	96	191	97	192
rect	97	191	98	192
rect	98	191	99	192
rect	99	191	100	192
rect	100	191	101	192
rect	101	191	102	192
rect	102	191	103	192
rect	103	191	104	192
rect	104	191	105	192
rect	105	191	106	192
rect	106	191	107	192
rect	107	191	108	192
rect	109	191	110	192
rect	110	191	111	192
rect	111	191	112	192
rect	112	191	113	192
rect	113	191	114	192
rect	114	191	115	192
rect	115	191	116	192
rect	116	191	117	192
rect	117	191	118	192
rect	118	191	119	192
rect	119	191	120	192
rect	120	191	121	192
rect	121	191	122	192
rect	122	191	123	192
rect	123	191	124	192
rect	124	191	125	192
rect	125	191	126	192
rect	126	191	127	192
rect	127	191	128	192
rect	128	191	129	192
rect	129	191	130	192
rect	130	191	131	192
rect	131	191	132	192
rect	132	191	133	192
rect	133	191	134	192
rect	134	191	135	192
rect	135	191	136	192
rect	136	191	137	192
rect	137	191	138	192
rect	138	191	139	192
rect	139	191	140	192
rect	140	191	141	192
rect	141	191	142	192
rect	142	191	143	192
rect	143	191	144	192
rect	144	191	145	192
rect	145	191	146	192
rect	146	191	147	192
rect	147	191	148	192
rect	148	191	149	192
rect	149	191	150	192
rect	150	191	151	192
rect	151	191	152	192
rect	152	191	153	192
rect	153	191	154	192
rect	154	191	155	192
rect	155	191	156	192
rect	156	191	157	192
rect	157	191	158	192
rect	158	191	159	192
rect	159	191	160	192
rect	161	191	162	192
rect	162	191	163	192
rect	163	191	164	192
rect	164	191	165	192
rect	165	191	166	192
rect	166	191	167	192
rect	167	191	168	192
rect	168	191	169	192
rect	169	191	170	192
rect	170	191	171	192
rect	171	191	172	192
rect	172	191	173	192
rect	173	191	174	192
rect	174	191	175	192
rect	175	191	176	192
rect	176	191	177	192
rect	177	191	178	192
rect	178	191	179	192
rect	179	191	180	192
rect	180	191	181	192
rect	181	191	182	192
rect	182	191	183	192
rect	183	191	184	192
rect	184	191	185	192
rect	185	191	186	192
rect	186	191	187	192
rect	187	191	188	192
rect	188	191	189	192
rect	189	191	190	192
rect	190	191	191	192
rect	191	191	192	192
rect	192	191	193	192
rect	193	191	194	192
rect	195	191	196	192
rect	196	191	197	192
rect	197	191	198	192
rect	198	191	199	192
rect	199	191	200	192
rect	200	191	201	192
rect	201	191	202	192
rect	202	191	203	192
rect	203	191	204	192
rect	204	191	205	192
rect	205	191	206	192
rect	206	191	207	192
rect	207	191	208	192
rect	208	191	209	192
rect	209	191	210	192
rect	210	191	211	192
rect	211	191	212	192
rect	212	191	213	192
rect	213	191	214	192
rect	214	191	215	192
rect	215	191	216	192
rect	216	191	217	192
rect	217	191	218	192
rect	218	191	219	192
rect	219	191	220	192
rect	220	191	221	192
rect	221	191	222	192
rect	223	191	224	192
rect	224	191	225	192
rect	225	191	226	192
rect	226	191	227	192
rect	227	191	228	192
rect	228	191	229	192
rect	229	191	230	192
rect	230	191	231	192
rect	231	191	232	192
rect	232	191	233	192
rect	233	191	234	192
rect	234	191	235	192
rect	235	191	236	192
rect	236	191	237	192
rect	237	191	238	192
rect	238	191	239	192
rect	239	191	240	192
rect	240	191	241	192
rect	241	191	242	192
rect	242	191	243	192
rect	243	191	244	192
rect	244	191	245	192
rect	245	191	246	192
rect	246	191	247	192
rect	247	191	248	192
rect	248	191	249	192
rect	249	191	250	192
rect	250	191	251	192
rect	251	191	252	192
rect	252	191	253	192
rect	253	191	254	192
rect	254	191	255	192
rect	255	191	256	192
rect	256	191	257	192
rect	257	191	258	192
rect	258	191	259	192
rect	259	191	260	192
rect	260	191	261	192
rect	261	191	262	192
rect	262	191	263	192
rect	263	191	264	192
rect	264	191	265	192
rect	265	191	266	192
rect	266	191	267	192
rect	267	191	268	192
rect	268	191	269	192
rect	269	191	270	192
rect	270	191	271	192
rect	271	191	272	192
rect	272	191	273	192
rect	273	191	274	192
rect	274	191	275	192
rect	275	191	276	192
rect	276	191	277	192
rect	277	191	278	192
rect	278	191	279	192
rect	279	191	280	192
rect	280	191	281	192
rect	281	191	282	192
rect	282	191	283	192
rect	283	191	284	192
rect	284	191	285	192
rect	285	191	286	192
rect	286	191	287	192
rect	287	191	288	192
rect	288	191	289	192
rect	289	191	290	192
rect	290	191	291	192
rect	291	191	292	192
rect	292	191	293	192
rect	293	191	294	192
rect	294	191	295	192
rect	295	191	296	192
rect	296	191	297	192
rect	297	191	298	192
rect	298	191	299	192
rect	299	191	300	192
rect	300	191	301	192
rect	301	191	302	192
rect	302	191	303	192
rect	303	191	304	192
rect	304	191	305	192
rect	305	191	306	192
rect	306	191	307	192
rect	307	191	308	192
rect	308	191	309	192
rect	309	191	310	192
rect	310	191	311	192
rect	311	191	312	192
rect	312	191	313	192
rect	313	191	314	192
rect	314	191	315	192
rect	315	191	316	192
rect	316	191	317	192
rect	317	191	318	192
rect	318	191	319	192
rect	319	191	320	192
rect	320	191	321	192
rect	321	191	322	192
rect	322	191	323	192
rect	323	191	324	192
rect	324	191	325	192
rect	325	191	326	192
rect	326	191	327	192
rect	327	191	328	192
rect	328	191	329	192
rect	329	191	330	192
rect	330	191	331	192
rect	331	191	332	192
rect	332	191	333	192
rect	333	191	334	192
rect	334	191	335	192
rect	335	191	336	192
rect	336	191	337	192
rect	337	191	338	192
rect	338	191	339	192
rect	339	191	340	192
rect	340	191	341	192
rect	341	191	342	192
rect	342	191	343	192
rect	343	191	344	192
rect	344	191	345	192
rect	345	191	346	192
rect	346	191	347	192
rect	347	191	348	192
rect	348	191	349	192
rect	349	191	350	192
rect	350	191	351	192
rect	351	191	352	192
rect	352	191	353	192
rect	353	191	354	192
rect	354	191	355	192
rect	355	191	356	192
rect	356	191	357	192
rect	357	191	358	192
rect	358	191	359	192
rect	359	191	360	192
rect	360	191	361	192
rect	361	191	362	192
rect	362	191	363	192
rect	363	191	364	192
rect	364	191	365	192
rect	365	191	366	192
rect	366	191	367	192
rect	367	191	368	192
rect	368	191	369	192
rect	369	191	370	192
rect	370	191	371	192
rect	371	191	372	192
rect	372	191	373	192
rect	373	191	374	192
rect	374	191	375	192
rect	375	191	376	192
rect	377	191	378	192
rect	378	191	379	192
rect	379	191	380	192
rect	380	191	381	192
rect	381	191	382	192
rect	382	191	383	192
rect	384	191	385	192
rect	385	191	386	192
rect	386	191	387	192
rect	387	191	388	192
rect	388	191	389	192
rect	389	191	390	192
rect	390	191	391	192
rect	391	191	392	192
rect	392	191	393	192
rect	393	191	394	192
rect	394	191	395	192
rect	395	191	396	192
rect	396	191	397	192
rect	397	191	398	192
rect	398	191	399	192
rect	0	217	1	218
rect	1	217	2	218
rect	2	217	3	218
rect	3	217	4	218
rect	4	217	5	218
rect	5	217	6	218
rect	7	217	8	218
rect	8	217	9	218
rect	9	217	10	218
rect	10	217	11	218
rect	11	217	12	218
rect	12	217	13	218
rect	13	217	14	218
rect	14	217	15	218
rect	15	217	16	218
rect	16	217	17	218
rect	17	217	18	218
rect	18	217	19	218
rect	19	217	20	218
rect	20	217	21	218
rect	21	217	22	218
rect	22	217	23	218
rect	23	217	24	218
rect	24	217	25	218
rect	25	217	26	218
rect	26	217	27	218
rect	27	217	28	218
rect	28	217	29	218
rect	29	217	30	218
rect	30	217	31	218
rect	31	217	32	218
rect	32	217	33	218
rect	33	217	34	218
rect	34	217	35	218
rect	35	217	36	218
rect	36	217	37	218
rect	37	217	38	218
rect	38	217	39	218
rect	39	217	40	218
rect	40	217	41	218
rect	41	217	42	218
rect	42	217	43	218
rect	43	217	44	218
rect	44	217	45	218
rect	45	217	46	218
rect	46	217	47	218
rect	47	217	48	218
rect	48	217	49	218
rect	49	217	50	218
rect	50	217	51	218
rect	51	217	52	218
rect	52	217	53	218
rect	53	217	54	218
rect	54	217	55	218
rect	55	217	56	218
rect	56	217	57	218
rect	57	217	58	218
rect	58	217	59	218
rect	59	217	60	218
rect	60	217	61	218
rect	61	217	62	218
rect	62	217	63	218
rect	63	217	64	218
rect	65	217	66	218
rect	66	217	67	218
rect	67	217	68	218
rect	68	217	69	218
rect	69	217	70	218
rect	70	217	71	218
rect	71	217	72	218
rect	72	217	73	218
rect	73	217	74	218
rect	74	217	75	218
rect	75	217	76	218
rect	76	217	77	218
rect	77	217	78	218
rect	78	217	79	218
rect	79	217	80	218
rect	80	217	81	218
rect	81	217	82	218
rect	82	217	83	218
rect	84	217	85	218
rect	85	217	86	218
rect	86	217	87	218
rect	87	217	88	218
rect	88	217	89	218
rect	89	217	90	218
rect	91	217	92	218
rect	92	217	93	218
rect	93	217	94	218
rect	94	217	95	218
rect	95	217	96	218
rect	96	217	97	218
rect	97	217	98	218
rect	98	217	99	218
rect	99	217	100	218
rect	100	217	101	218
rect	101	217	102	218
rect	102	217	103	218
rect	103	217	104	218
rect	104	217	105	218
rect	105	217	106	218
rect	106	217	107	218
rect	107	217	108	218
rect	108	217	109	218
rect	110	217	111	218
rect	111	217	112	218
rect	112	217	113	218
rect	113	217	114	218
rect	114	217	115	218
rect	115	217	116	218
rect	116	217	117	218
rect	117	217	118	218
rect	118	217	119	218
rect	119	217	120	218
rect	120	217	121	218
rect	121	217	122	218
rect	122	217	123	218
rect	123	217	124	218
rect	124	217	125	218
rect	125	217	126	218
rect	126	217	127	218
rect	127	217	128	218
rect	128	217	129	218
rect	129	217	130	218
rect	130	217	131	218
rect	131	217	132	218
rect	132	217	133	218
rect	133	217	134	218
rect	134	217	135	218
rect	135	217	136	218
rect	136	217	137	218
rect	137	217	138	218
rect	138	217	139	218
rect	139	217	140	218
rect	140	217	141	218
rect	141	217	142	218
rect	142	217	143	218
rect	143	217	144	218
rect	144	217	145	218
rect	145	217	146	218
rect	146	217	147	218
rect	147	217	148	218
rect	148	217	149	218
rect	149	217	150	218
rect	150	217	151	218
rect	151	217	152	218
rect	152	217	153	218
rect	153	217	154	218
rect	154	217	155	218
rect	155	217	156	218
rect	156	217	157	218
rect	157	217	158	218
rect	158	217	159	218
rect	159	217	160	218
rect	160	217	161	218
rect	161	217	162	218
rect	162	217	163	218
rect	163	217	164	218
rect	164	217	165	218
rect	165	217	166	218
rect	166	217	167	218
rect	167	217	168	218
rect	168	217	169	218
rect	169	217	170	218
rect	170	217	171	218
rect	171	217	172	218
rect	172	217	173	218
rect	173	217	174	218
rect	174	217	175	218
rect	175	217	176	218
rect	176	217	177	218
rect	177	217	178	218
rect	178	217	179	218
rect	179	217	180	218
rect	180	217	181	218
rect	181	217	182	218
rect	182	217	183	218
rect	183	217	184	218
rect	184	217	185	218
rect	185	217	186	218
rect	186	217	187	218
rect	187	217	188	218
rect	189	217	190	218
rect	190	217	191	218
rect	191	217	192	218
rect	192	217	193	218
rect	193	217	194	218
rect	194	217	195	218
rect	196	217	197	218
rect	197	217	198	218
rect	198	217	199	218
rect	199	217	200	218
rect	200	217	201	218
rect	201	217	202	218
rect	202	217	203	218
rect	203	217	204	218
rect	204	217	205	218
rect	205	217	206	218
rect	206	217	207	218
rect	207	217	208	218
rect	208	217	209	218
rect	209	217	210	218
rect	210	217	211	218
rect	211	217	212	218
rect	212	217	213	218
rect	213	217	214	218
rect	214	217	215	218
rect	215	217	216	218
rect	216	217	217	218
rect	217	217	218	218
rect	218	217	219	218
rect	219	217	220	218
rect	220	217	221	218
rect	221	217	222	218
rect	222	217	223	218
rect	223	217	224	218
rect	224	217	225	218
rect	225	217	226	218
rect	226	217	227	218
rect	227	217	228	218
rect	228	217	229	218
rect	229	217	230	218
rect	230	217	231	218
rect	231	217	232	218
rect	232	217	233	218
rect	233	217	234	218
rect	234	217	235	218
rect	236	217	237	218
rect	237	217	238	218
rect	238	217	239	218
rect	239	217	240	218
rect	240	217	241	218
rect	241	217	242	218
rect	242	217	243	218
rect	243	217	244	218
rect	244	217	245	218
rect	245	217	246	218
rect	246	217	247	218
rect	247	217	248	218
rect	248	217	249	218
rect	249	217	250	218
rect	250	217	251	218
rect	251	217	252	218
rect	252	217	253	218
rect	253	217	254	218
rect	254	217	255	218
rect	255	217	256	218
rect	256	217	257	218
rect	257	217	258	218
rect	258	217	259	218
rect	259	217	260	218
rect	260	217	261	218
rect	261	217	262	218
rect	262	217	263	218
rect	263	217	264	218
rect	264	217	265	218
rect	265	217	266	218
rect	266	217	267	218
rect	267	217	268	218
rect	268	217	269	218
rect	269	217	270	218
rect	270	217	271	218
rect	271	217	272	218
rect	272	217	273	218
rect	273	217	274	218
rect	274	217	275	218
rect	275	217	276	218
rect	276	217	277	218
rect	277	217	278	218
rect	278	217	279	218
rect	279	217	280	218
rect	280	217	281	218
rect	281	217	282	218
rect	282	217	283	218
rect	283	217	284	218
rect	284	217	285	218
rect	285	217	286	218
rect	286	217	287	218
rect	287	217	288	218
rect	288	217	289	218
rect	289	217	290	218
rect	290	217	291	218
rect	291	217	292	218
rect	292	217	293	218
rect	294	217	295	218
rect	295	217	296	218
rect	296	217	297	218
rect	297	217	298	218
rect	298	217	299	218
rect	299	217	300	218
rect	300	217	301	218
rect	301	217	302	218
rect	302	217	303	218
rect	303	217	304	218
rect	304	217	305	218
rect	305	217	306	218
rect	306	217	307	218
rect	307	217	308	218
rect	308	217	309	218
rect	309	217	310	218
rect	310	217	311	218
rect	311	217	312	218
rect	312	217	313	218
rect	313	217	314	218
rect	314	217	315	218
rect	315	217	316	218
rect	316	217	317	218
rect	317	217	318	218
rect	318	217	319	218
rect	319	217	320	218
rect	320	217	321	218
rect	321	217	322	218
rect	322	217	323	218
rect	323	217	324	218
rect	324	217	325	218
rect	325	217	326	218
rect	326	217	327	218
rect	327	217	328	218
rect	328	217	329	218
rect	329	217	330	218
rect	330	217	331	218
rect	331	217	332	218
rect	332	217	333	218
rect	333	217	334	218
rect	334	217	335	218
rect	335	217	336	218
rect	336	217	337	218
rect	337	217	338	218
rect	338	217	339	218
rect	339	217	340	218
rect	340	217	341	218
rect	341	217	342	218
rect	342	217	343	218
rect	343	217	344	218
rect	344	217	345	218
rect	345	217	346	218
rect	346	217	347	218
rect	347	217	348	218
rect	348	217	349	218
rect	349	217	350	218
rect	350	217	351	218
rect	351	217	352	218
rect	352	217	353	218
rect	353	217	354	218
rect	354	217	355	218
rect	355	217	356	218
rect	356	217	357	218
rect	357	217	358	218
rect	358	217	359	218
rect	359	217	360	218
rect	361	217	362	218
rect	362	217	363	218
rect	363	217	364	218
rect	364	217	365	218
rect	365	217	366	218
rect	366	217	367	218
rect	367	217	368	218
rect	368	217	369	218
rect	369	217	370	218
rect	370	217	371	218
rect	371	217	372	218
rect	372	217	373	218
rect	373	217	374	218
rect	374	217	375	218
rect	375	217	376	218
rect	376	217	377	218
rect	377	217	378	218
rect	378	217	379	218
rect	380	217	381	218
rect	381	217	382	218
rect	382	217	383	218
rect	383	217	384	218
rect	384	217	385	218
rect	385	217	386	218
rect	386	217	387	218
rect	387	217	388	218
rect	388	217	389	218
rect	0	218	1	219
rect	1	218	2	219
rect	2	218	3	219
rect	3	218	4	219
rect	4	218	5	219
rect	5	218	6	219
rect	7	218	8	219
rect	8	218	9	219
rect	9	218	10	219
rect	10	218	11	219
rect	11	218	12	219
rect	12	218	13	219
rect	13	218	14	219
rect	14	218	15	219
rect	15	218	16	219
rect	16	218	17	219
rect	17	218	18	219
rect	18	218	19	219
rect	19	218	20	219
rect	20	218	21	219
rect	21	218	22	219
rect	22	218	23	219
rect	23	218	24	219
rect	24	218	25	219
rect	25	218	26	219
rect	26	218	27	219
rect	27	218	28	219
rect	28	218	29	219
rect	29	218	30	219
rect	30	218	31	219
rect	31	218	32	219
rect	32	218	33	219
rect	33	218	34	219
rect	34	218	35	219
rect	35	218	36	219
rect	36	218	37	219
rect	37	218	38	219
rect	38	218	39	219
rect	39	218	40	219
rect	40	218	41	219
rect	41	218	42	219
rect	42	218	43	219
rect	43	218	44	219
rect	44	218	45	219
rect	45	218	46	219
rect	46	218	47	219
rect	47	218	48	219
rect	48	218	49	219
rect	49	218	50	219
rect	50	218	51	219
rect	51	218	52	219
rect	52	218	53	219
rect	53	218	54	219
rect	54	218	55	219
rect	55	218	56	219
rect	56	218	57	219
rect	57	218	58	219
rect	58	218	59	219
rect	59	218	60	219
rect	60	218	61	219
rect	61	218	62	219
rect	62	218	63	219
rect	63	218	64	219
rect	65	218	66	219
rect	66	218	67	219
rect	67	218	68	219
rect	68	218	69	219
rect	69	218	70	219
rect	70	218	71	219
rect	71	218	72	219
rect	72	218	73	219
rect	73	218	74	219
rect	74	218	75	219
rect	75	218	76	219
rect	76	218	77	219
rect	77	218	78	219
rect	78	218	79	219
rect	79	218	80	219
rect	80	218	81	219
rect	81	218	82	219
rect	82	218	83	219
rect	84	218	85	219
rect	85	218	86	219
rect	86	218	87	219
rect	87	218	88	219
rect	88	218	89	219
rect	89	218	90	219
rect	91	218	92	219
rect	92	218	93	219
rect	93	218	94	219
rect	94	218	95	219
rect	95	218	96	219
rect	96	218	97	219
rect	97	218	98	219
rect	98	218	99	219
rect	99	218	100	219
rect	100	218	101	219
rect	101	218	102	219
rect	102	218	103	219
rect	103	218	104	219
rect	104	218	105	219
rect	105	218	106	219
rect	106	218	107	219
rect	107	218	108	219
rect	108	218	109	219
rect	110	218	111	219
rect	111	218	112	219
rect	112	218	113	219
rect	113	218	114	219
rect	114	218	115	219
rect	115	218	116	219
rect	116	218	117	219
rect	117	218	118	219
rect	118	218	119	219
rect	119	218	120	219
rect	120	218	121	219
rect	121	218	122	219
rect	122	218	123	219
rect	123	218	124	219
rect	124	218	125	219
rect	125	218	126	219
rect	126	218	127	219
rect	127	218	128	219
rect	128	218	129	219
rect	129	218	130	219
rect	130	218	131	219
rect	131	218	132	219
rect	132	218	133	219
rect	133	218	134	219
rect	134	218	135	219
rect	135	218	136	219
rect	136	218	137	219
rect	137	218	138	219
rect	138	218	139	219
rect	139	218	140	219
rect	140	218	141	219
rect	141	218	142	219
rect	142	218	143	219
rect	143	218	144	219
rect	144	218	145	219
rect	145	218	146	219
rect	146	218	147	219
rect	147	218	148	219
rect	148	218	149	219
rect	149	218	150	219
rect	150	218	151	219
rect	151	218	152	219
rect	152	218	153	219
rect	153	218	154	219
rect	154	218	155	219
rect	155	218	156	219
rect	156	218	157	219
rect	157	218	158	219
rect	158	218	159	219
rect	159	218	160	219
rect	160	218	161	219
rect	161	218	162	219
rect	162	218	163	219
rect	163	218	164	219
rect	164	218	165	219
rect	165	218	166	219
rect	166	218	167	219
rect	167	218	168	219
rect	168	218	169	219
rect	169	218	170	219
rect	170	218	171	219
rect	171	218	172	219
rect	172	218	173	219
rect	173	218	174	219
rect	174	218	175	219
rect	175	218	176	219
rect	176	218	177	219
rect	177	218	178	219
rect	178	218	179	219
rect	179	218	180	219
rect	180	218	181	219
rect	181	218	182	219
rect	182	218	183	219
rect	183	218	184	219
rect	184	218	185	219
rect	185	218	186	219
rect	186	218	187	219
rect	187	218	188	219
rect	189	218	190	219
rect	190	218	191	219
rect	191	218	192	219
rect	192	218	193	219
rect	193	218	194	219
rect	194	218	195	219
rect	196	218	197	219
rect	197	218	198	219
rect	198	218	199	219
rect	199	218	200	219
rect	200	218	201	219
rect	201	218	202	219
rect	202	218	203	219
rect	203	218	204	219
rect	204	218	205	219
rect	205	218	206	219
rect	206	218	207	219
rect	207	218	208	219
rect	208	218	209	219
rect	209	218	210	219
rect	210	218	211	219
rect	211	218	212	219
rect	212	218	213	219
rect	213	218	214	219
rect	214	218	215	219
rect	215	218	216	219
rect	216	218	217	219
rect	217	218	218	219
rect	218	218	219	219
rect	219	218	220	219
rect	220	218	221	219
rect	221	218	222	219
rect	222	218	223	219
rect	223	218	224	219
rect	224	218	225	219
rect	225	218	226	219
rect	226	218	227	219
rect	227	218	228	219
rect	228	218	229	219
rect	229	218	230	219
rect	230	218	231	219
rect	231	218	232	219
rect	232	218	233	219
rect	233	218	234	219
rect	234	218	235	219
rect	236	218	237	219
rect	237	218	238	219
rect	238	218	239	219
rect	239	218	240	219
rect	240	218	241	219
rect	241	218	242	219
rect	242	218	243	219
rect	243	218	244	219
rect	244	218	245	219
rect	245	218	246	219
rect	246	218	247	219
rect	247	218	248	219
rect	248	218	249	219
rect	249	218	250	219
rect	250	218	251	219
rect	251	218	252	219
rect	252	218	253	219
rect	253	218	254	219
rect	254	218	255	219
rect	255	218	256	219
rect	256	218	257	219
rect	257	218	258	219
rect	258	218	259	219
rect	259	218	260	219
rect	260	218	261	219
rect	261	218	262	219
rect	262	218	263	219
rect	263	218	264	219
rect	264	218	265	219
rect	265	218	266	219
rect	266	218	267	219
rect	267	218	268	219
rect	268	218	269	219
rect	269	218	270	219
rect	270	218	271	219
rect	271	218	272	219
rect	272	218	273	219
rect	273	218	274	219
rect	274	218	275	219
rect	275	218	276	219
rect	276	218	277	219
rect	277	218	278	219
rect	278	218	279	219
rect	279	218	280	219
rect	280	218	281	219
rect	281	218	282	219
rect	282	218	283	219
rect	283	218	284	219
rect	284	218	285	219
rect	285	218	286	219
rect	286	218	287	219
rect	287	218	288	219
rect	288	218	289	219
rect	289	218	290	219
rect	290	218	291	219
rect	291	218	292	219
rect	292	218	293	219
rect	294	218	295	219
rect	295	218	296	219
rect	296	218	297	219
rect	297	218	298	219
rect	298	218	299	219
rect	299	218	300	219
rect	300	218	301	219
rect	301	218	302	219
rect	302	218	303	219
rect	303	218	304	219
rect	304	218	305	219
rect	305	218	306	219
rect	306	218	307	219
rect	307	218	308	219
rect	308	218	309	219
rect	309	218	310	219
rect	310	218	311	219
rect	311	218	312	219
rect	312	218	313	219
rect	313	218	314	219
rect	314	218	315	219
rect	315	218	316	219
rect	316	218	317	219
rect	317	218	318	219
rect	318	218	319	219
rect	319	218	320	219
rect	320	218	321	219
rect	321	218	322	219
rect	322	218	323	219
rect	323	218	324	219
rect	324	218	325	219
rect	325	218	326	219
rect	326	218	327	219
rect	327	218	328	219
rect	328	218	329	219
rect	329	218	330	219
rect	330	218	331	219
rect	331	218	332	219
rect	332	218	333	219
rect	333	218	334	219
rect	334	218	335	219
rect	335	218	336	219
rect	336	218	337	219
rect	337	218	338	219
rect	338	218	339	219
rect	339	218	340	219
rect	340	218	341	219
rect	341	218	342	219
rect	342	218	343	219
rect	343	218	344	219
rect	344	218	345	219
rect	345	218	346	219
rect	346	218	347	219
rect	347	218	348	219
rect	348	218	349	219
rect	349	218	350	219
rect	350	218	351	219
rect	351	218	352	219
rect	352	218	353	219
rect	353	218	354	219
rect	354	218	355	219
rect	355	218	356	219
rect	356	218	357	219
rect	357	218	358	219
rect	358	218	359	219
rect	359	218	360	219
rect	361	218	362	219
rect	362	218	363	219
rect	363	218	364	219
rect	364	218	365	219
rect	365	218	366	219
rect	366	218	367	219
rect	367	218	368	219
rect	368	218	369	219
rect	369	218	370	219
rect	370	218	371	219
rect	371	218	372	219
rect	372	218	373	219
rect	373	218	374	219
rect	374	218	375	219
rect	375	218	376	219
rect	376	218	377	219
rect	377	218	378	219
rect	378	218	379	219
rect	380	218	381	219
rect	381	218	382	219
rect	382	218	383	219
rect	383	218	384	219
rect	384	218	385	219
rect	385	218	386	219
rect	386	218	387	219
rect	387	218	388	219
rect	388	218	389	219
rect	0	219	1	220
rect	1	219	2	220
rect	2	219	3	220
rect	3	219	4	220
rect	4	219	5	220
rect	5	219	6	220
rect	7	219	8	220
rect	8	219	9	220
rect	9	219	10	220
rect	10	219	11	220
rect	11	219	12	220
rect	12	219	13	220
rect	13	219	14	220
rect	14	219	15	220
rect	15	219	16	220
rect	16	219	17	220
rect	17	219	18	220
rect	18	219	19	220
rect	19	219	20	220
rect	20	219	21	220
rect	21	219	22	220
rect	22	219	23	220
rect	23	219	24	220
rect	24	219	25	220
rect	25	219	26	220
rect	26	219	27	220
rect	27	219	28	220
rect	28	219	29	220
rect	29	219	30	220
rect	30	219	31	220
rect	31	219	32	220
rect	32	219	33	220
rect	33	219	34	220
rect	34	219	35	220
rect	35	219	36	220
rect	36	219	37	220
rect	37	219	38	220
rect	38	219	39	220
rect	39	219	40	220
rect	40	219	41	220
rect	41	219	42	220
rect	42	219	43	220
rect	43	219	44	220
rect	44	219	45	220
rect	45	219	46	220
rect	46	219	47	220
rect	47	219	48	220
rect	48	219	49	220
rect	49	219	50	220
rect	50	219	51	220
rect	51	219	52	220
rect	52	219	53	220
rect	53	219	54	220
rect	54	219	55	220
rect	55	219	56	220
rect	56	219	57	220
rect	57	219	58	220
rect	58	219	59	220
rect	59	219	60	220
rect	60	219	61	220
rect	61	219	62	220
rect	62	219	63	220
rect	63	219	64	220
rect	65	219	66	220
rect	66	219	67	220
rect	67	219	68	220
rect	68	219	69	220
rect	69	219	70	220
rect	70	219	71	220
rect	71	219	72	220
rect	72	219	73	220
rect	73	219	74	220
rect	74	219	75	220
rect	75	219	76	220
rect	76	219	77	220
rect	77	219	78	220
rect	78	219	79	220
rect	79	219	80	220
rect	80	219	81	220
rect	81	219	82	220
rect	82	219	83	220
rect	84	219	85	220
rect	85	219	86	220
rect	86	219	87	220
rect	87	219	88	220
rect	88	219	89	220
rect	89	219	90	220
rect	91	219	92	220
rect	92	219	93	220
rect	93	219	94	220
rect	94	219	95	220
rect	95	219	96	220
rect	96	219	97	220
rect	97	219	98	220
rect	98	219	99	220
rect	99	219	100	220
rect	100	219	101	220
rect	101	219	102	220
rect	102	219	103	220
rect	103	219	104	220
rect	104	219	105	220
rect	105	219	106	220
rect	106	219	107	220
rect	107	219	108	220
rect	108	219	109	220
rect	110	219	111	220
rect	111	219	112	220
rect	112	219	113	220
rect	113	219	114	220
rect	114	219	115	220
rect	115	219	116	220
rect	116	219	117	220
rect	117	219	118	220
rect	118	219	119	220
rect	119	219	120	220
rect	120	219	121	220
rect	121	219	122	220
rect	122	219	123	220
rect	123	219	124	220
rect	124	219	125	220
rect	125	219	126	220
rect	126	219	127	220
rect	127	219	128	220
rect	128	219	129	220
rect	129	219	130	220
rect	130	219	131	220
rect	131	219	132	220
rect	132	219	133	220
rect	133	219	134	220
rect	134	219	135	220
rect	135	219	136	220
rect	136	219	137	220
rect	137	219	138	220
rect	138	219	139	220
rect	139	219	140	220
rect	140	219	141	220
rect	141	219	142	220
rect	142	219	143	220
rect	143	219	144	220
rect	144	219	145	220
rect	145	219	146	220
rect	146	219	147	220
rect	147	219	148	220
rect	148	219	149	220
rect	149	219	150	220
rect	150	219	151	220
rect	151	219	152	220
rect	152	219	153	220
rect	153	219	154	220
rect	154	219	155	220
rect	155	219	156	220
rect	156	219	157	220
rect	157	219	158	220
rect	158	219	159	220
rect	159	219	160	220
rect	160	219	161	220
rect	161	219	162	220
rect	162	219	163	220
rect	163	219	164	220
rect	164	219	165	220
rect	165	219	166	220
rect	166	219	167	220
rect	167	219	168	220
rect	168	219	169	220
rect	169	219	170	220
rect	170	219	171	220
rect	171	219	172	220
rect	172	219	173	220
rect	173	219	174	220
rect	174	219	175	220
rect	175	219	176	220
rect	176	219	177	220
rect	177	219	178	220
rect	178	219	179	220
rect	179	219	180	220
rect	180	219	181	220
rect	181	219	182	220
rect	182	219	183	220
rect	183	219	184	220
rect	184	219	185	220
rect	185	219	186	220
rect	186	219	187	220
rect	187	219	188	220
rect	189	219	190	220
rect	190	219	191	220
rect	191	219	192	220
rect	192	219	193	220
rect	193	219	194	220
rect	194	219	195	220
rect	196	219	197	220
rect	197	219	198	220
rect	198	219	199	220
rect	199	219	200	220
rect	200	219	201	220
rect	201	219	202	220
rect	202	219	203	220
rect	203	219	204	220
rect	204	219	205	220
rect	205	219	206	220
rect	206	219	207	220
rect	207	219	208	220
rect	208	219	209	220
rect	209	219	210	220
rect	210	219	211	220
rect	211	219	212	220
rect	212	219	213	220
rect	213	219	214	220
rect	214	219	215	220
rect	215	219	216	220
rect	216	219	217	220
rect	217	219	218	220
rect	218	219	219	220
rect	219	219	220	220
rect	220	219	221	220
rect	221	219	222	220
rect	222	219	223	220
rect	223	219	224	220
rect	224	219	225	220
rect	225	219	226	220
rect	226	219	227	220
rect	227	219	228	220
rect	228	219	229	220
rect	229	219	230	220
rect	230	219	231	220
rect	231	219	232	220
rect	232	219	233	220
rect	233	219	234	220
rect	234	219	235	220
rect	236	219	237	220
rect	237	219	238	220
rect	238	219	239	220
rect	239	219	240	220
rect	240	219	241	220
rect	241	219	242	220
rect	242	219	243	220
rect	243	219	244	220
rect	244	219	245	220
rect	245	219	246	220
rect	246	219	247	220
rect	247	219	248	220
rect	248	219	249	220
rect	249	219	250	220
rect	250	219	251	220
rect	251	219	252	220
rect	252	219	253	220
rect	253	219	254	220
rect	254	219	255	220
rect	255	219	256	220
rect	256	219	257	220
rect	257	219	258	220
rect	258	219	259	220
rect	259	219	260	220
rect	260	219	261	220
rect	261	219	262	220
rect	262	219	263	220
rect	263	219	264	220
rect	264	219	265	220
rect	265	219	266	220
rect	266	219	267	220
rect	267	219	268	220
rect	268	219	269	220
rect	269	219	270	220
rect	270	219	271	220
rect	271	219	272	220
rect	272	219	273	220
rect	273	219	274	220
rect	274	219	275	220
rect	275	219	276	220
rect	276	219	277	220
rect	277	219	278	220
rect	278	219	279	220
rect	279	219	280	220
rect	280	219	281	220
rect	281	219	282	220
rect	282	219	283	220
rect	283	219	284	220
rect	284	219	285	220
rect	285	219	286	220
rect	286	219	287	220
rect	287	219	288	220
rect	288	219	289	220
rect	289	219	290	220
rect	290	219	291	220
rect	291	219	292	220
rect	292	219	293	220
rect	294	219	295	220
rect	295	219	296	220
rect	296	219	297	220
rect	297	219	298	220
rect	298	219	299	220
rect	299	219	300	220
rect	300	219	301	220
rect	301	219	302	220
rect	302	219	303	220
rect	303	219	304	220
rect	304	219	305	220
rect	305	219	306	220
rect	306	219	307	220
rect	307	219	308	220
rect	308	219	309	220
rect	309	219	310	220
rect	310	219	311	220
rect	311	219	312	220
rect	312	219	313	220
rect	313	219	314	220
rect	314	219	315	220
rect	315	219	316	220
rect	316	219	317	220
rect	317	219	318	220
rect	318	219	319	220
rect	319	219	320	220
rect	320	219	321	220
rect	321	219	322	220
rect	322	219	323	220
rect	323	219	324	220
rect	324	219	325	220
rect	325	219	326	220
rect	326	219	327	220
rect	327	219	328	220
rect	328	219	329	220
rect	329	219	330	220
rect	330	219	331	220
rect	331	219	332	220
rect	332	219	333	220
rect	333	219	334	220
rect	334	219	335	220
rect	335	219	336	220
rect	336	219	337	220
rect	337	219	338	220
rect	338	219	339	220
rect	339	219	340	220
rect	340	219	341	220
rect	341	219	342	220
rect	342	219	343	220
rect	343	219	344	220
rect	344	219	345	220
rect	345	219	346	220
rect	346	219	347	220
rect	347	219	348	220
rect	348	219	349	220
rect	349	219	350	220
rect	350	219	351	220
rect	351	219	352	220
rect	352	219	353	220
rect	353	219	354	220
rect	354	219	355	220
rect	355	219	356	220
rect	356	219	357	220
rect	357	219	358	220
rect	358	219	359	220
rect	359	219	360	220
rect	361	219	362	220
rect	362	219	363	220
rect	363	219	364	220
rect	364	219	365	220
rect	365	219	366	220
rect	366	219	367	220
rect	367	219	368	220
rect	368	219	369	220
rect	369	219	370	220
rect	370	219	371	220
rect	371	219	372	220
rect	372	219	373	220
rect	373	219	374	220
rect	374	219	375	220
rect	375	219	376	220
rect	376	219	377	220
rect	377	219	378	220
rect	378	219	379	220
rect	380	219	381	220
rect	381	219	382	220
rect	382	219	383	220
rect	383	219	384	220
rect	384	219	385	220
rect	385	219	386	220
rect	386	219	387	220
rect	387	219	388	220
rect	388	219	389	220
rect	0	220	1	221
rect	1	220	2	221
rect	2	220	3	221
rect	3	220	4	221
rect	4	220	5	221
rect	5	220	6	221
rect	7	220	8	221
rect	8	220	9	221
rect	9	220	10	221
rect	10	220	11	221
rect	11	220	12	221
rect	12	220	13	221
rect	13	220	14	221
rect	14	220	15	221
rect	15	220	16	221
rect	16	220	17	221
rect	17	220	18	221
rect	18	220	19	221
rect	19	220	20	221
rect	20	220	21	221
rect	21	220	22	221
rect	22	220	23	221
rect	23	220	24	221
rect	24	220	25	221
rect	25	220	26	221
rect	26	220	27	221
rect	27	220	28	221
rect	28	220	29	221
rect	29	220	30	221
rect	30	220	31	221
rect	31	220	32	221
rect	32	220	33	221
rect	33	220	34	221
rect	34	220	35	221
rect	35	220	36	221
rect	36	220	37	221
rect	37	220	38	221
rect	38	220	39	221
rect	39	220	40	221
rect	40	220	41	221
rect	41	220	42	221
rect	42	220	43	221
rect	43	220	44	221
rect	44	220	45	221
rect	45	220	46	221
rect	46	220	47	221
rect	47	220	48	221
rect	48	220	49	221
rect	49	220	50	221
rect	50	220	51	221
rect	51	220	52	221
rect	52	220	53	221
rect	53	220	54	221
rect	54	220	55	221
rect	55	220	56	221
rect	56	220	57	221
rect	57	220	58	221
rect	58	220	59	221
rect	59	220	60	221
rect	60	220	61	221
rect	61	220	62	221
rect	62	220	63	221
rect	63	220	64	221
rect	65	220	66	221
rect	66	220	67	221
rect	67	220	68	221
rect	68	220	69	221
rect	69	220	70	221
rect	70	220	71	221
rect	71	220	72	221
rect	72	220	73	221
rect	73	220	74	221
rect	74	220	75	221
rect	75	220	76	221
rect	76	220	77	221
rect	77	220	78	221
rect	78	220	79	221
rect	79	220	80	221
rect	80	220	81	221
rect	81	220	82	221
rect	82	220	83	221
rect	84	220	85	221
rect	85	220	86	221
rect	86	220	87	221
rect	87	220	88	221
rect	88	220	89	221
rect	89	220	90	221
rect	91	220	92	221
rect	92	220	93	221
rect	93	220	94	221
rect	94	220	95	221
rect	95	220	96	221
rect	96	220	97	221
rect	97	220	98	221
rect	98	220	99	221
rect	99	220	100	221
rect	100	220	101	221
rect	101	220	102	221
rect	102	220	103	221
rect	103	220	104	221
rect	104	220	105	221
rect	105	220	106	221
rect	106	220	107	221
rect	107	220	108	221
rect	108	220	109	221
rect	110	220	111	221
rect	111	220	112	221
rect	112	220	113	221
rect	113	220	114	221
rect	114	220	115	221
rect	115	220	116	221
rect	116	220	117	221
rect	117	220	118	221
rect	118	220	119	221
rect	119	220	120	221
rect	120	220	121	221
rect	121	220	122	221
rect	122	220	123	221
rect	123	220	124	221
rect	124	220	125	221
rect	125	220	126	221
rect	126	220	127	221
rect	127	220	128	221
rect	128	220	129	221
rect	129	220	130	221
rect	130	220	131	221
rect	131	220	132	221
rect	132	220	133	221
rect	133	220	134	221
rect	134	220	135	221
rect	135	220	136	221
rect	136	220	137	221
rect	137	220	138	221
rect	138	220	139	221
rect	139	220	140	221
rect	140	220	141	221
rect	141	220	142	221
rect	142	220	143	221
rect	143	220	144	221
rect	144	220	145	221
rect	145	220	146	221
rect	146	220	147	221
rect	147	220	148	221
rect	148	220	149	221
rect	149	220	150	221
rect	150	220	151	221
rect	151	220	152	221
rect	152	220	153	221
rect	153	220	154	221
rect	154	220	155	221
rect	155	220	156	221
rect	156	220	157	221
rect	157	220	158	221
rect	158	220	159	221
rect	159	220	160	221
rect	160	220	161	221
rect	161	220	162	221
rect	162	220	163	221
rect	163	220	164	221
rect	164	220	165	221
rect	165	220	166	221
rect	166	220	167	221
rect	167	220	168	221
rect	168	220	169	221
rect	169	220	170	221
rect	170	220	171	221
rect	171	220	172	221
rect	172	220	173	221
rect	173	220	174	221
rect	174	220	175	221
rect	175	220	176	221
rect	176	220	177	221
rect	177	220	178	221
rect	178	220	179	221
rect	179	220	180	221
rect	180	220	181	221
rect	181	220	182	221
rect	182	220	183	221
rect	183	220	184	221
rect	184	220	185	221
rect	185	220	186	221
rect	186	220	187	221
rect	187	220	188	221
rect	189	220	190	221
rect	190	220	191	221
rect	191	220	192	221
rect	192	220	193	221
rect	193	220	194	221
rect	194	220	195	221
rect	196	220	197	221
rect	197	220	198	221
rect	198	220	199	221
rect	199	220	200	221
rect	200	220	201	221
rect	201	220	202	221
rect	202	220	203	221
rect	203	220	204	221
rect	204	220	205	221
rect	205	220	206	221
rect	206	220	207	221
rect	207	220	208	221
rect	208	220	209	221
rect	209	220	210	221
rect	210	220	211	221
rect	211	220	212	221
rect	212	220	213	221
rect	213	220	214	221
rect	214	220	215	221
rect	215	220	216	221
rect	216	220	217	221
rect	217	220	218	221
rect	218	220	219	221
rect	219	220	220	221
rect	220	220	221	221
rect	221	220	222	221
rect	222	220	223	221
rect	223	220	224	221
rect	224	220	225	221
rect	225	220	226	221
rect	226	220	227	221
rect	227	220	228	221
rect	228	220	229	221
rect	229	220	230	221
rect	230	220	231	221
rect	231	220	232	221
rect	232	220	233	221
rect	233	220	234	221
rect	234	220	235	221
rect	236	220	237	221
rect	237	220	238	221
rect	238	220	239	221
rect	239	220	240	221
rect	240	220	241	221
rect	241	220	242	221
rect	242	220	243	221
rect	243	220	244	221
rect	244	220	245	221
rect	245	220	246	221
rect	246	220	247	221
rect	247	220	248	221
rect	248	220	249	221
rect	249	220	250	221
rect	250	220	251	221
rect	251	220	252	221
rect	252	220	253	221
rect	253	220	254	221
rect	254	220	255	221
rect	255	220	256	221
rect	256	220	257	221
rect	257	220	258	221
rect	258	220	259	221
rect	259	220	260	221
rect	260	220	261	221
rect	261	220	262	221
rect	262	220	263	221
rect	263	220	264	221
rect	264	220	265	221
rect	265	220	266	221
rect	266	220	267	221
rect	267	220	268	221
rect	268	220	269	221
rect	269	220	270	221
rect	270	220	271	221
rect	271	220	272	221
rect	272	220	273	221
rect	273	220	274	221
rect	274	220	275	221
rect	275	220	276	221
rect	276	220	277	221
rect	277	220	278	221
rect	278	220	279	221
rect	279	220	280	221
rect	280	220	281	221
rect	281	220	282	221
rect	282	220	283	221
rect	283	220	284	221
rect	284	220	285	221
rect	285	220	286	221
rect	286	220	287	221
rect	287	220	288	221
rect	288	220	289	221
rect	289	220	290	221
rect	290	220	291	221
rect	291	220	292	221
rect	292	220	293	221
rect	294	220	295	221
rect	295	220	296	221
rect	296	220	297	221
rect	297	220	298	221
rect	298	220	299	221
rect	299	220	300	221
rect	300	220	301	221
rect	301	220	302	221
rect	302	220	303	221
rect	303	220	304	221
rect	304	220	305	221
rect	305	220	306	221
rect	306	220	307	221
rect	307	220	308	221
rect	308	220	309	221
rect	309	220	310	221
rect	310	220	311	221
rect	311	220	312	221
rect	312	220	313	221
rect	313	220	314	221
rect	314	220	315	221
rect	315	220	316	221
rect	316	220	317	221
rect	317	220	318	221
rect	318	220	319	221
rect	319	220	320	221
rect	320	220	321	221
rect	321	220	322	221
rect	322	220	323	221
rect	323	220	324	221
rect	324	220	325	221
rect	325	220	326	221
rect	326	220	327	221
rect	327	220	328	221
rect	328	220	329	221
rect	329	220	330	221
rect	330	220	331	221
rect	331	220	332	221
rect	332	220	333	221
rect	333	220	334	221
rect	334	220	335	221
rect	335	220	336	221
rect	336	220	337	221
rect	337	220	338	221
rect	338	220	339	221
rect	339	220	340	221
rect	340	220	341	221
rect	341	220	342	221
rect	342	220	343	221
rect	343	220	344	221
rect	344	220	345	221
rect	345	220	346	221
rect	346	220	347	221
rect	347	220	348	221
rect	348	220	349	221
rect	349	220	350	221
rect	350	220	351	221
rect	351	220	352	221
rect	352	220	353	221
rect	353	220	354	221
rect	354	220	355	221
rect	355	220	356	221
rect	356	220	357	221
rect	357	220	358	221
rect	358	220	359	221
rect	359	220	360	221
rect	361	220	362	221
rect	362	220	363	221
rect	363	220	364	221
rect	364	220	365	221
rect	365	220	366	221
rect	366	220	367	221
rect	367	220	368	221
rect	368	220	369	221
rect	369	220	370	221
rect	370	220	371	221
rect	371	220	372	221
rect	372	220	373	221
rect	373	220	374	221
rect	374	220	375	221
rect	375	220	376	221
rect	376	220	377	221
rect	377	220	378	221
rect	378	220	379	221
rect	380	220	381	221
rect	381	220	382	221
rect	382	220	383	221
rect	383	220	384	221
rect	384	220	385	221
rect	385	220	386	221
rect	386	220	387	221
rect	387	220	388	221
rect	388	220	389	221
rect	0	221	1	222
rect	1	221	2	222
rect	2	221	3	222
rect	3	221	4	222
rect	4	221	5	222
rect	5	221	6	222
rect	7	221	8	222
rect	8	221	9	222
rect	9	221	10	222
rect	10	221	11	222
rect	11	221	12	222
rect	12	221	13	222
rect	13	221	14	222
rect	14	221	15	222
rect	15	221	16	222
rect	16	221	17	222
rect	17	221	18	222
rect	18	221	19	222
rect	19	221	20	222
rect	20	221	21	222
rect	21	221	22	222
rect	22	221	23	222
rect	23	221	24	222
rect	24	221	25	222
rect	25	221	26	222
rect	26	221	27	222
rect	27	221	28	222
rect	28	221	29	222
rect	29	221	30	222
rect	30	221	31	222
rect	31	221	32	222
rect	32	221	33	222
rect	33	221	34	222
rect	34	221	35	222
rect	35	221	36	222
rect	36	221	37	222
rect	37	221	38	222
rect	38	221	39	222
rect	39	221	40	222
rect	40	221	41	222
rect	41	221	42	222
rect	42	221	43	222
rect	43	221	44	222
rect	44	221	45	222
rect	45	221	46	222
rect	46	221	47	222
rect	47	221	48	222
rect	48	221	49	222
rect	49	221	50	222
rect	50	221	51	222
rect	51	221	52	222
rect	52	221	53	222
rect	53	221	54	222
rect	54	221	55	222
rect	55	221	56	222
rect	56	221	57	222
rect	57	221	58	222
rect	58	221	59	222
rect	59	221	60	222
rect	60	221	61	222
rect	61	221	62	222
rect	62	221	63	222
rect	63	221	64	222
rect	65	221	66	222
rect	66	221	67	222
rect	67	221	68	222
rect	68	221	69	222
rect	69	221	70	222
rect	70	221	71	222
rect	71	221	72	222
rect	72	221	73	222
rect	73	221	74	222
rect	74	221	75	222
rect	75	221	76	222
rect	76	221	77	222
rect	77	221	78	222
rect	78	221	79	222
rect	79	221	80	222
rect	80	221	81	222
rect	81	221	82	222
rect	82	221	83	222
rect	84	221	85	222
rect	85	221	86	222
rect	86	221	87	222
rect	87	221	88	222
rect	88	221	89	222
rect	89	221	90	222
rect	91	221	92	222
rect	92	221	93	222
rect	93	221	94	222
rect	94	221	95	222
rect	95	221	96	222
rect	96	221	97	222
rect	97	221	98	222
rect	98	221	99	222
rect	99	221	100	222
rect	100	221	101	222
rect	101	221	102	222
rect	102	221	103	222
rect	103	221	104	222
rect	104	221	105	222
rect	105	221	106	222
rect	106	221	107	222
rect	107	221	108	222
rect	108	221	109	222
rect	110	221	111	222
rect	111	221	112	222
rect	112	221	113	222
rect	113	221	114	222
rect	114	221	115	222
rect	115	221	116	222
rect	116	221	117	222
rect	117	221	118	222
rect	118	221	119	222
rect	119	221	120	222
rect	120	221	121	222
rect	121	221	122	222
rect	122	221	123	222
rect	123	221	124	222
rect	124	221	125	222
rect	125	221	126	222
rect	126	221	127	222
rect	127	221	128	222
rect	128	221	129	222
rect	129	221	130	222
rect	130	221	131	222
rect	131	221	132	222
rect	132	221	133	222
rect	133	221	134	222
rect	134	221	135	222
rect	135	221	136	222
rect	136	221	137	222
rect	137	221	138	222
rect	138	221	139	222
rect	139	221	140	222
rect	140	221	141	222
rect	141	221	142	222
rect	142	221	143	222
rect	143	221	144	222
rect	144	221	145	222
rect	145	221	146	222
rect	146	221	147	222
rect	147	221	148	222
rect	148	221	149	222
rect	149	221	150	222
rect	150	221	151	222
rect	151	221	152	222
rect	152	221	153	222
rect	153	221	154	222
rect	154	221	155	222
rect	155	221	156	222
rect	156	221	157	222
rect	157	221	158	222
rect	158	221	159	222
rect	159	221	160	222
rect	160	221	161	222
rect	161	221	162	222
rect	162	221	163	222
rect	163	221	164	222
rect	164	221	165	222
rect	165	221	166	222
rect	166	221	167	222
rect	167	221	168	222
rect	168	221	169	222
rect	169	221	170	222
rect	170	221	171	222
rect	171	221	172	222
rect	172	221	173	222
rect	173	221	174	222
rect	174	221	175	222
rect	175	221	176	222
rect	176	221	177	222
rect	177	221	178	222
rect	178	221	179	222
rect	179	221	180	222
rect	180	221	181	222
rect	181	221	182	222
rect	182	221	183	222
rect	183	221	184	222
rect	184	221	185	222
rect	185	221	186	222
rect	186	221	187	222
rect	187	221	188	222
rect	189	221	190	222
rect	190	221	191	222
rect	191	221	192	222
rect	192	221	193	222
rect	193	221	194	222
rect	194	221	195	222
rect	196	221	197	222
rect	197	221	198	222
rect	198	221	199	222
rect	199	221	200	222
rect	200	221	201	222
rect	201	221	202	222
rect	202	221	203	222
rect	203	221	204	222
rect	204	221	205	222
rect	205	221	206	222
rect	206	221	207	222
rect	207	221	208	222
rect	208	221	209	222
rect	209	221	210	222
rect	210	221	211	222
rect	211	221	212	222
rect	212	221	213	222
rect	213	221	214	222
rect	214	221	215	222
rect	215	221	216	222
rect	216	221	217	222
rect	217	221	218	222
rect	218	221	219	222
rect	219	221	220	222
rect	220	221	221	222
rect	221	221	222	222
rect	222	221	223	222
rect	223	221	224	222
rect	224	221	225	222
rect	225	221	226	222
rect	226	221	227	222
rect	227	221	228	222
rect	228	221	229	222
rect	229	221	230	222
rect	230	221	231	222
rect	231	221	232	222
rect	232	221	233	222
rect	233	221	234	222
rect	234	221	235	222
rect	236	221	237	222
rect	237	221	238	222
rect	238	221	239	222
rect	239	221	240	222
rect	240	221	241	222
rect	241	221	242	222
rect	242	221	243	222
rect	243	221	244	222
rect	244	221	245	222
rect	245	221	246	222
rect	246	221	247	222
rect	247	221	248	222
rect	248	221	249	222
rect	249	221	250	222
rect	250	221	251	222
rect	251	221	252	222
rect	252	221	253	222
rect	253	221	254	222
rect	254	221	255	222
rect	255	221	256	222
rect	256	221	257	222
rect	257	221	258	222
rect	258	221	259	222
rect	259	221	260	222
rect	260	221	261	222
rect	261	221	262	222
rect	262	221	263	222
rect	263	221	264	222
rect	264	221	265	222
rect	265	221	266	222
rect	266	221	267	222
rect	267	221	268	222
rect	268	221	269	222
rect	269	221	270	222
rect	270	221	271	222
rect	271	221	272	222
rect	272	221	273	222
rect	273	221	274	222
rect	274	221	275	222
rect	275	221	276	222
rect	276	221	277	222
rect	277	221	278	222
rect	278	221	279	222
rect	279	221	280	222
rect	280	221	281	222
rect	281	221	282	222
rect	282	221	283	222
rect	283	221	284	222
rect	284	221	285	222
rect	285	221	286	222
rect	286	221	287	222
rect	287	221	288	222
rect	288	221	289	222
rect	289	221	290	222
rect	290	221	291	222
rect	291	221	292	222
rect	292	221	293	222
rect	294	221	295	222
rect	295	221	296	222
rect	296	221	297	222
rect	297	221	298	222
rect	298	221	299	222
rect	299	221	300	222
rect	300	221	301	222
rect	301	221	302	222
rect	302	221	303	222
rect	303	221	304	222
rect	304	221	305	222
rect	305	221	306	222
rect	306	221	307	222
rect	307	221	308	222
rect	308	221	309	222
rect	309	221	310	222
rect	310	221	311	222
rect	311	221	312	222
rect	312	221	313	222
rect	313	221	314	222
rect	314	221	315	222
rect	315	221	316	222
rect	316	221	317	222
rect	317	221	318	222
rect	318	221	319	222
rect	319	221	320	222
rect	320	221	321	222
rect	321	221	322	222
rect	322	221	323	222
rect	323	221	324	222
rect	324	221	325	222
rect	325	221	326	222
rect	326	221	327	222
rect	327	221	328	222
rect	328	221	329	222
rect	329	221	330	222
rect	330	221	331	222
rect	331	221	332	222
rect	332	221	333	222
rect	333	221	334	222
rect	334	221	335	222
rect	335	221	336	222
rect	336	221	337	222
rect	337	221	338	222
rect	338	221	339	222
rect	339	221	340	222
rect	340	221	341	222
rect	341	221	342	222
rect	342	221	343	222
rect	343	221	344	222
rect	344	221	345	222
rect	345	221	346	222
rect	346	221	347	222
rect	347	221	348	222
rect	348	221	349	222
rect	349	221	350	222
rect	350	221	351	222
rect	351	221	352	222
rect	352	221	353	222
rect	353	221	354	222
rect	354	221	355	222
rect	355	221	356	222
rect	356	221	357	222
rect	357	221	358	222
rect	358	221	359	222
rect	359	221	360	222
rect	361	221	362	222
rect	362	221	363	222
rect	363	221	364	222
rect	364	221	365	222
rect	365	221	366	222
rect	366	221	367	222
rect	367	221	368	222
rect	368	221	369	222
rect	369	221	370	222
rect	370	221	371	222
rect	371	221	372	222
rect	372	221	373	222
rect	373	221	374	222
rect	374	221	375	222
rect	375	221	376	222
rect	376	221	377	222
rect	377	221	378	222
rect	378	221	379	222
rect	380	221	381	222
rect	381	221	382	222
rect	382	221	383	222
rect	383	221	384	222
rect	384	221	385	222
rect	385	221	386	222
rect	386	221	387	222
rect	387	221	388	222
rect	388	221	389	222
rect	0	222	1	223
rect	1	222	2	223
rect	2	222	3	223
rect	3	222	4	223
rect	4	222	5	223
rect	5	222	6	223
rect	7	222	8	223
rect	8	222	9	223
rect	9	222	10	223
rect	10	222	11	223
rect	11	222	12	223
rect	12	222	13	223
rect	13	222	14	223
rect	14	222	15	223
rect	15	222	16	223
rect	16	222	17	223
rect	17	222	18	223
rect	18	222	19	223
rect	19	222	20	223
rect	20	222	21	223
rect	21	222	22	223
rect	22	222	23	223
rect	23	222	24	223
rect	24	222	25	223
rect	25	222	26	223
rect	26	222	27	223
rect	27	222	28	223
rect	28	222	29	223
rect	29	222	30	223
rect	30	222	31	223
rect	31	222	32	223
rect	32	222	33	223
rect	33	222	34	223
rect	34	222	35	223
rect	35	222	36	223
rect	36	222	37	223
rect	37	222	38	223
rect	38	222	39	223
rect	39	222	40	223
rect	40	222	41	223
rect	41	222	42	223
rect	42	222	43	223
rect	43	222	44	223
rect	44	222	45	223
rect	45	222	46	223
rect	46	222	47	223
rect	47	222	48	223
rect	48	222	49	223
rect	49	222	50	223
rect	50	222	51	223
rect	51	222	52	223
rect	52	222	53	223
rect	53	222	54	223
rect	54	222	55	223
rect	55	222	56	223
rect	56	222	57	223
rect	57	222	58	223
rect	58	222	59	223
rect	59	222	60	223
rect	60	222	61	223
rect	61	222	62	223
rect	62	222	63	223
rect	63	222	64	223
rect	65	222	66	223
rect	66	222	67	223
rect	67	222	68	223
rect	68	222	69	223
rect	69	222	70	223
rect	70	222	71	223
rect	71	222	72	223
rect	72	222	73	223
rect	73	222	74	223
rect	74	222	75	223
rect	75	222	76	223
rect	76	222	77	223
rect	77	222	78	223
rect	78	222	79	223
rect	79	222	80	223
rect	80	222	81	223
rect	81	222	82	223
rect	82	222	83	223
rect	84	222	85	223
rect	85	222	86	223
rect	86	222	87	223
rect	87	222	88	223
rect	88	222	89	223
rect	89	222	90	223
rect	91	222	92	223
rect	92	222	93	223
rect	93	222	94	223
rect	94	222	95	223
rect	95	222	96	223
rect	96	222	97	223
rect	97	222	98	223
rect	98	222	99	223
rect	99	222	100	223
rect	100	222	101	223
rect	101	222	102	223
rect	102	222	103	223
rect	103	222	104	223
rect	104	222	105	223
rect	105	222	106	223
rect	106	222	107	223
rect	107	222	108	223
rect	108	222	109	223
rect	110	222	111	223
rect	111	222	112	223
rect	112	222	113	223
rect	113	222	114	223
rect	114	222	115	223
rect	115	222	116	223
rect	116	222	117	223
rect	117	222	118	223
rect	118	222	119	223
rect	119	222	120	223
rect	120	222	121	223
rect	121	222	122	223
rect	122	222	123	223
rect	123	222	124	223
rect	124	222	125	223
rect	125	222	126	223
rect	126	222	127	223
rect	127	222	128	223
rect	128	222	129	223
rect	129	222	130	223
rect	130	222	131	223
rect	131	222	132	223
rect	132	222	133	223
rect	133	222	134	223
rect	134	222	135	223
rect	135	222	136	223
rect	136	222	137	223
rect	137	222	138	223
rect	138	222	139	223
rect	139	222	140	223
rect	140	222	141	223
rect	141	222	142	223
rect	142	222	143	223
rect	143	222	144	223
rect	144	222	145	223
rect	145	222	146	223
rect	146	222	147	223
rect	147	222	148	223
rect	148	222	149	223
rect	149	222	150	223
rect	150	222	151	223
rect	151	222	152	223
rect	152	222	153	223
rect	153	222	154	223
rect	154	222	155	223
rect	155	222	156	223
rect	156	222	157	223
rect	157	222	158	223
rect	158	222	159	223
rect	159	222	160	223
rect	160	222	161	223
rect	161	222	162	223
rect	162	222	163	223
rect	163	222	164	223
rect	164	222	165	223
rect	165	222	166	223
rect	166	222	167	223
rect	167	222	168	223
rect	168	222	169	223
rect	169	222	170	223
rect	170	222	171	223
rect	171	222	172	223
rect	172	222	173	223
rect	173	222	174	223
rect	174	222	175	223
rect	175	222	176	223
rect	176	222	177	223
rect	177	222	178	223
rect	178	222	179	223
rect	179	222	180	223
rect	180	222	181	223
rect	181	222	182	223
rect	182	222	183	223
rect	183	222	184	223
rect	184	222	185	223
rect	185	222	186	223
rect	186	222	187	223
rect	187	222	188	223
rect	189	222	190	223
rect	190	222	191	223
rect	191	222	192	223
rect	192	222	193	223
rect	193	222	194	223
rect	194	222	195	223
rect	196	222	197	223
rect	197	222	198	223
rect	198	222	199	223
rect	199	222	200	223
rect	200	222	201	223
rect	201	222	202	223
rect	202	222	203	223
rect	203	222	204	223
rect	204	222	205	223
rect	205	222	206	223
rect	206	222	207	223
rect	207	222	208	223
rect	208	222	209	223
rect	209	222	210	223
rect	210	222	211	223
rect	211	222	212	223
rect	212	222	213	223
rect	213	222	214	223
rect	214	222	215	223
rect	215	222	216	223
rect	216	222	217	223
rect	217	222	218	223
rect	218	222	219	223
rect	219	222	220	223
rect	220	222	221	223
rect	221	222	222	223
rect	222	222	223	223
rect	223	222	224	223
rect	224	222	225	223
rect	225	222	226	223
rect	226	222	227	223
rect	227	222	228	223
rect	228	222	229	223
rect	229	222	230	223
rect	230	222	231	223
rect	231	222	232	223
rect	232	222	233	223
rect	233	222	234	223
rect	234	222	235	223
rect	236	222	237	223
rect	237	222	238	223
rect	238	222	239	223
rect	239	222	240	223
rect	240	222	241	223
rect	241	222	242	223
rect	242	222	243	223
rect	243	222	244	223
rect	244	222	245	223
rect	245	222	246	223
rect	246	222	247	223
rect	247	222	248	223
rect	248	222	249	223
rect	249	222	250	223
rect	250	222	251	223
rect	251	222	252	223
rect	252	222	253	223
rect	253	222	254	223
rect	254	222	255	223
rect	255	222	256	223
rect	256	222	257	223
rect	257	222	258	223
rect	258	222	259	223
rect	259	222	260	223
rect	260	222	261	223
rect	261	222	262	223
rect	262	222	263	223
rect	263	222	264	223
rect	264	222	265	223
rect	265	222	266	223
rect	266	222	267	223
rect	267	222	268	223
rect	268	222	269	223
rect	269	222	270	223
rect	270	222	271	223
rect	271	222	272	223
rect	272	222	273	223
rect	273	222	274	223
rect	274	222	275	223
rect	275	222	276	223
rect	276	222	277	223
rect	277	222	278	223
rect	278	222	279	223
rect	279	222	280	223
rect	280	222	281	223
rect	281	222	282	223
rect	282	222	283	223
rect	283	222	284	223
rect	284	222	285	223
rect	285	222	286	223
rect	286	222	287	223
rect	287	222	288	223
rect	288	222	289	223
rect	289	222	290	223
rect	290	222	291	223
rect	291	222	292	223
rect	292	222	293	223
rect	294	222	295	223
rect	295	222	296	223
rect	296	222	297	223
rect	297	222	298	223
rect	298	222	299	223
rect	299	222	300	223
rect	300	222	301	223
rect	301	222	302	223
rect	302	222	303	223
rect	303	222	304	223
rect	304	222	305	223
rect	305	222	306	223
rect	306	222	307	223
rect	307	222	308	223
rect	308	222	309	223
rect	309	222	310	223
rect	310	222	311	223
rect	311	222	312	223
rect	312	222	313	223
rect	313	222	314	223
rect	314	222	315	223
rect	315	222	316	223
rect	316	222	317	223
rect	317	222	318	223
rect	318	222	319	223
rect	319	222	320	223
rect	320	222	321	223
rect	321	222	322	223
rect	322	222	323	223
rect	323	222	324	223
rect	324	222	325	223
rect	325	222	326	223
rect	326	222	327	223
rect	327	222	328	223
rect	328	222	329	223
rect	329	222	330	223
rect	330	222	331	223
rect	331	222	332	223
rect	332	222	333	223
rect	333	222	334	223
rect	334	222	335	223
rect	335	222	336	223
rect	336	222	337	223
rect	337	222	338	223
rect	338	222	339	223
rect	339	222	340	223
rect	340	222	341	223
rect	341	222	342	223
rect	342	222	343	223
rect	343	222	344	223
rect	344	222	345	223
rect	345	222	346	223
rect	346	222	347	223
rect	347	222	348	223
rect	348	222	349	223
rect	349	222	350	223
rect	350	222	351	223
rect	351	222	352	223
rect	352	222	353	223
rect	353	222	354	223
rect	354	222	355	223
rect	355	222	356	223
rect	356	222	357	223
rect	357	222	358	223
rect	358	222	359	223
rect	359	222	360	223
rect	361	222	362	223
rect	362	222	363	223
rect	363	222	364	223
rect	364	222	365	223
rect	365	222	366	223
rect	366	222	367	223
rect	367	222	368	223
rect	368	222	369	223
rect	369	222	370	223
rect	370	222	371	223
rect	371	222	372	223
rect	372	222	373	223
rect	373	222	374	223
rect	374	222	375	223
rect	375	222	376	223
rect	376	222	377	223
rect	377	222	378	223
rect	378	222	379	223
rect	380	222	381	223
rect	381	222	382	223
rect	382	222	383	223
rect	383	222	384	223
rect	384	222	385	223
rect	385	222	386	223
rect	386	222	387	223
rect	387	222	388	223
rect	388	222	389	223
rect	0	248	1	249
rect	1	248	2	249
rect	2	248	3	249
rect	3	248	4	249
rect	4	248	5	249
rect	5	248	6	249
rect	7	248	8	249
rect	8	248	9	249
rect	9	248	10	249
rect	10	248	11	249
rect	11	248	12	249
rect	12	248	13	249
rect	14	248	15	249
rect	15	248	16	249
rect	16	248	17	249
rect	17	248	18	249
rect	18	248	19	249
rect	19	248	20	249
rect	20	248	21	249
rect	21	248	22	249
rect	22	248	23	249
rect	23	248	24	249
rect	24	248	25	249
rect	25	248	26	249
rect	26	248	27	249
rect	27	248	28	249
rect	28	248	29	249
rect	29	248	30	249
rect	30	248	31	249
rect	31	248	32	249
rect	32	248	33	249
rect	33	248	34	249
rect	34	248	35	249
rect	35	248	36	249
rect	36	248	37	249
rect	37	248	38	249
rect	38	248	39	249
rect	39	248	40	249
rect	40	248	41	249
rect	41	248	42	249
rect	42	248	43	249
rect	43	248	44	249
rect	44	248	45	249
rect	45	248	46	249
rect	46	248	47	249
rect	47	248	48	249
rect	48	248	49	249
rect	49	248	50	249
rect	50	248	51	249
rect	51	248	52	249
rect	52	248	53	249
rect	53	248	54	249
rect	54	248	55	249
rect	55	248	56	249
rect	56	248	57	249
rect	57	248	58	249
rect	58	248	59	249
rect	59	248	60	249
rect	60	248	61	249
rect	61	248	62	249
rect	62	248	63	249
rect	63	248	64	249
rect	64	248	65	249
rect	65	248	66	249
rect	66	248	67	249
rect	67	248	68	249
rect	69	248	70	249
rect	70	248	71	249
rect	71	248	72	249
rect	72	248	73	249
rect	73	248	74	249
rect	74	248	75	249
rect	76	248	77	249
rect	77	248	78	249
rect	78	248	79	249
rect	79	248	80	249
rect	80	248	81	249
rect	81	248	82	249
rect	82	248	83	249
rect	83	248	84	249
rect	84	248	85	249
rect	85	248	86	249
rect	86	248	87	249
rect	87	248	88	249
rect	88	248	89	249
rect	89	248	90	249
rect	90	248	91	249
rect	92	248	93	249
rect	93	248	94	249
rect	94	248	95	249
rect	95	248	96	249
rect	96	248	97	249
rect	97	248	98	249
rect	99	248	100	249
rect	100	248	101	249
rect	101	248	102	249
rect	102	248	103	249
rect	103	248	104	249
rect	104	248	105	249
rect	105	248	106	249
rect	106	248	107	249
rect	107	248	108	249
rect	108	248	109	249
rect	109	248	110	249
rect	110	248	111	249
rect	111	248	112	249
rect	112	248	113	249
rect	113	248	114	249
rect	114	248	115	249
rect	115	248	116	249
rect	116	248	117	249
rect	117	248	118	249
rect	118	248	119	249
rect	119	248	120	249
rect	120	248	121	249
rect	121	248	122	249
rect	122	248	123	249
rect	123	248	124	249
rect	124	248	125	249
rect	125	248	126	249
rect	127	248	128	249
rect	128	248	129	249
rect	129	248	130	249
rect	130	248	131	249
rect	131	248	132	249
rect	132	248	133	249
rect	133	248	134	249
rect	134	248	135	249
rect	135	248	136	249
rect	136	248	137	249
rect	137	248	138	249
rect	138	248	139	249
rect	139	248	140	249
rect	140	248	141	249
rect	141	248	142	249
rect	142	248	143	249
rect	143	248	144	249
rect	144	248	145	249
rect	145	248	146	249
rect	146	248	147	249
rect	147	248	148	249
rect	148	248	149	249
rect	149	248	150	249
rect	150	248	151	249
rect	151	248	152	249
rect	152	248	153	249
rect	153	248	154	249
rect	154	248	155	249
rect	155	248	156	249
rect	156	248	157	249
rect	157	248	158	249
rect	158	248	159	249
rect	159	248	160	249
rect	160	248	161	249
rect	161	248	162	249
rect	162	248	163	249
rect	163	248	164	249
rect	164	248	165	249
rect	165	248	166	249
rect	166	248	167	249
rect	167	248	168	249
rect	168	248	169	249
rect	169	248	170	249
rect	170	248	171	249
rect	171	248	172	249
rect	172	248	173	249
rect	173	248	174	249
rect	174	248	175	249
rect	175	248	176	249
rect	176	248	177	249
rect	177	248	178	249
rect	178	248	179	249
rect	179	248	180	249
rect	180	248	181	249
rect	181	248	182	249
rect	182	248	183	249
rect	183	248	184	249
rect	184	248	185	249
rect	185	248	186	249
rect	186	248	187	249
rect	187	248	188	249
rect	188	248	189	249
rect	189	248	190	249
rect	190	248	191	249
rect	191	248	192	249
rect	192	248	193	249
rect	193	248	194	249
rect	194	248	195	249
rect	195	248	196	249
rect	196	248	197	249
rect	197	248	198	249
rect	198	248	199	249
rect	199	248	200	249
rect	200	248	201	249
rect	201	248	202	249
rect	202	248	203	249
rect	203	248	204	249
rect	204	248	205	249
rect	206	248	207	249
rect	207	248	208	249
rect	208	248	209	249
rect	209	248	210	249
rect	210	248	211	249
rect	211	248	212	249
rect	213	248	214	249
rect	214	248	215	249
rect	215	248	216	249
rect	216	248	217	249
rect	217	248	218	249
rect	218	248	219	249
rect	219	248	220	249
rect	220	248	221	249
rect	221	248	222	249
rect	222	248	223	249
rect	223	248	224	249
rect	224	248	225	249
rect	225	248	226	249
rect	226	248	227	249
rect	227	248	228	249
rect	228	248	229	249
rect	229	248	230	249
rect	230	248	231	249
rect	231	248	232	249
rect	232	248	233	249
rect	233	248	234	249
rect	234	248	235	249
rect	235	248	236	249
rect	236	248	237	249
rect	237	248	238	249
rect	238	248	239	249
rect	239	248	240	249
rect	241	248	242	249
rect	242	248	243	249
rect	243	248	244	249
rect	244	248	245	249
rect	245	248	246	249
rect	246	248	247	249
rect	247	248	248	249
rect	248	248	249	249
rect	249	248	250	249
rect	250	248	251	249
rect	251	248	252	249
rect	252	248	253	249
rect	253	248	254	249
rect	254	248	255	249
rect	255	248	256	249
rect	256	248	257	249
rect	257	248	258	249
rect	258	248	259	249
rect	259	248	260	249
rect	260	248	261	249
rect	261	248	262	249
rect	262	248	263	249
rect	263	248	264	249
rect	264	248	265	249
rect	265	248	266	249
rect	266	248	267	249
rect	267	248	268	249
rect	268	248	269	249
rect	269	248	270	249
rect	270	248	271	249
rect	271	248	272	249
rect	272	248	273	249
rect	273	248	274	249
rect	274	248	275	249
rect	275	248	276	249
rect	276	248	277	249
rect	277	248	278	249
rect	278	248	279	249
rect	279	248	280	249
rect	280	248	281	249
rect	281	248	282	249
rect	282	248	283	249
rect	283	248	284	249
rect	284	248	285	249
rect	285	248	286	249
rect	286	248	287	249
rect	287	248	288	249
rect	288	248	289	249
rect	289	248	290	249
rect	290	248	291	249
rect	291	248	292	249
rect	292	248	293	249
rect	293	248	294	249
rect	294	248	295	249
rect	295	248	296	249
rect	296	248	297	249
rect	297	248	298	249
rect	298	248	299	249
rect	299	248	300	249
rect	300	248	301	249
rect	301	248	302	249
rect	302	248	303	249
rect	303	248	304	249
rect	304	248	305	249
rect	305	248	306	249
rect	306	248	307	249
rect	307	248	308	249
rect	308	248	309	249
rect	309	248	310	249
rect	310	248	311	249
rect	311	248	312	249
rect	312	248	313	249
rect	313	248	314	249
rect	314	248	315	249
rect	315	248	316	249
rect	317	248	318	249
rect	318	248	319	249
rect	319	248	320	249
rect	320	248	321	249
rect	321	248	322	249
rect	322	248	323	249
rect	323	248	324	249
rect	324	248	325	249
rect	325	248	326	249
rect	326	248	327	249
rect	327	248	328	249
rect	328	248	329	249
rect	329	248	330	249
rect	330	248	331	249
rect	331	248	332	249
rect	332	248	333	249
rect	333	248	334	249
rect	334	248	335	249
rect	335	248	336	249
rect	336	248	337	249
rect	337	248	338	249
rect	338	248	339	249
rect	339	248	340	249
rect	340	248	341	249
rect	341	248	342	249
rect	342	248	343	249
rect	343	248	344	249
rect	344	248	345	249
rect	345	248	346	249
rect	346	248	347	249
rect	347	248	348	249
rect	348	248	349	249
rect	349	248	350	249
rect	350	248	351	249
rect	351	248	352	249
rect	352	248	353	249
rect	353	248	354	249
rect	354	248	355	249
rect	355	248	356	249
rect	356	248	357	249
rect	357	248	358	249
rect	358	248	359	249
rect	359	248	360	249
rect	360	248	361	249
rect	361	248	362	249
rect	362	248	363	249
rect	363	248	364	249
rect	364	248	365	249
rect	366	248	367	249
rect	367	248	368	249
rect	368	248	369	249
rect	369	248	370	249
rect	370	248	371	249
rect	371	248	372	249
rect	372	248	373	249
rect	373	248	374	249
rect	374	248	375	249
rect	375	248	376	249
rect	376	248	377	249
rect	377	248	378	249
rect	378	248	379	249
rect	379	248	380	249
rect	380	248	381	249
rect	0	249	1	250
rect	1	249	2	250
rect	2	249	3	250
rect	3	249	4	250
rect	4	249	5	250
rect	5	249	6	250
rect	7	249	8	250
rect	8	249	9	250
rect	9	249	10	250
rect	10	249	11	250
rect	11	249	12	250
rect	12	249	13	250
rect	14	249	15	250
rect	15	249	16	250
rect	16	249	17	250
rect	17	249	18	250
rect	18	249	19	250
rect	19	249	20	250
rect	20	249	21	250
rect	21	249	22	250
rect	22	249	23	250
rect	23	249	24	250
rect	24	249	25	250
rect	25	249	26	250
rect	26	249	27	250
rect	27	249	28	250
rect	28	249	29	250
rect	29	249	30	250
rect	30	249	31	250
rect	31	249	32	250
rect	32	249	33	250
rect	33	249	34	250
rect	34	249	35	250
rect	35	249	36	250
rect	36	249	37	250
rect	37	249	38	250
rect	38	249	39	250
rect	39	249	40	250
rect	40	249	41	250
rect	41	249	42	250
rect	42	249	43	250
rect	43	249	44	250
rect	44	249	45	250
rect	45	249	46	250
rect	46	249	47	250
rect	47	249	48	250
rect	48	249	49	250
rect	49	249	50	250
rect	50	249	51	250
rect	51	249	52	250
rect	52	249	53	250
rect	53	249	54	250
rect	54	249	55	250
rect	55	249	56	250
rect	56	249	57	250
rect	57	249	58	250
rect	58	249	59	250
rect	59	249	60	250
rect	60	249	61	250
rect	61	249	62	250
rect	62	249	63	250
rect	63	249	64	250
rect	64	249	65	250
rect	65	249	66	250
rect	66	249	67	250
rect	67	249	68	250
rect	69	249	70	250
rect	70	249	71	250
rect	71	249	72	250
rect	72	249	73	250
rect	73	249	74	250
rect	74	249	75	250
rect	76	249	77	250
rect	77	249	78	250
rect	78	249	79	250
rect	79	249	80	250
rect	80	249	81	250
rect	81	249	82	250
rect	82	249	83	250
rect	83	249	84	250
rect	84	249	85	250
rect	85	249	86	250
rect	86	249	87	250
rect	87	249	88	250
rect	88	249	89	250
rect	89	249	90	250
rect	90	249	91	250
rect	92	249	93	250
rect	93	249	94	250
rect	94	249	95	250
rect	95	249	96	250
rect	96	249	97	250
rect	97	249	98	250
rect	99	249	100	250
rect	100	249	101	250
rect	101	249	102	250
rect	102	249	103	250
rect	103	249	104	250
rect	104	249	105	250
rect	105	249	106	250
rect	106	249	107	250
rect	107	249	108	250
rect	108	249	109	250
rect	109	249	110	250
rect	110	249	111	250
rect	111	249	112	250
rect	112	249	113	250
rect	113	249	114	250
rect	114	249	115	250
rect	115	249	116	250
rect	116	249	117	250
rect	117	249	118	250
rect	118	249	119	250
rect	119	249	120	250
rect	120	249	121	250
rect	121	249	122	250
rect	122	249	123	250
rect	123	249	124	250
rect	124	249	125	250
rect	125	249	126	250
rect	127	249	128	250
rect	128	249	129	250
rect	129	249	130	250
rect	130	249	131	250
rect	131	249	132	250
rect	132	249	133	250
rect	133	249	134	250
rect	134	249	135	250
rect	135	249	136	250
rect	136	249	137	250
rect	137	249	138	250
rect	138	249	139	250
rect	139	249	140	250
rect	140	249	141	250
rect	141	249	142	250
rect	142	249	143	250
rect	143	249	144	250
rect	144	249	145	250
rect	145	249	146	250
rect	146	249	147	250
rect	147	249	148	250
rect	148	249	149	250
rect	149	249	150	250
rect	150	249	151	250
rect	151	249	152	250
rect	152	249	153	250
rect	153	249	154	250
rect	154	249	155	250
rect	155	249	156	250
rect	156	249	157	250
rect	157	249	158	250
rect	158	249	159	250
rect	159	249	160	250
rect	160	249	161	250
rect	161	249	162	250
rect	162	249	163	250
rect	163	249	164	250
rect	164	249	165	250
rect	165	249	166	250
rect	166	249	167	250
rect	167	249	168	250
rect	168	249	169	250
rect	169	249	170	250
rect	170	249	171	250
rect	171	249	172	250
rect	172	249	173	250
rect	173	249	174	250
rect	174	249	175	250
rect	175	249	176	250
rect	176	249	177	250
rect	177	249	178	250
rect	178	249	179	250
rect	179	249	180	250
rect	180	249	181	250
rect	181	249	182	250
rect	182	249	183	250
rect	183	249	184	250
rect	184	249	185	250
rect	185	249	186	250
rect	186	249	187	250
rect	187	249	188	250
rect	188	249	189	250
rect	189	249	190	250
rect	190	249	191	250
rect	191	249	192	250
rect	192	249	193	250
rect	193	249	194	250
rect	194	249	195	250
rect	195	249	196	250
rect	196	249	197	250
rect	197	249	198	250
rect	198	249	199	250
rect	199	249	200	250
rect	200	249	201	250
rect	201	249	202	250
rect	202	249	203	250
rect	203	249	204	250
rect	204	249	205	250
rect	206	249	207	250
rect	207	249	208	250
rect	208	249	209	250
rect	209	249	210	250
rect	210	249	211	250
rect	211	249	212	250
rect	213	249	214	250
rect	214	249	215	250
rect	215	249	216	250
rect	216	249	217	250
rect	217	249	218	250
rect	218	249	219	250
rect	219	249	220	250
rect	220	249	221	250
rect	221	249	222	250
rect	222	249	223	250
rect	223	249	224	250
rect	224	249	225	250
rect	225	249	226	250
rect	226	249	227	250
rect	227	249	228	250
rect	228	249	229	250
rect	229	249	230	250
rect	230	249	231	250
rect	231	249	232	250
rect	232	249	233	250
rect	233	249	234	250
rect	234	249	235	250
rect	235	249	236	250
rect	236	249	237	250
rect	237	249	238	250
rect	238	249	239	250
rect	239	249	240	250
rect	241	249	242	250
rect	242	249	243	250
rect	243	249	244	250
rect	244	249	245	250
rect	245	249	246	250
rect	246	249	247	250
rect	247	249	248	250
rect	248	249	249	250
rect	249	249	250	250
rect	250	249	251	250
rect	251	249	252	250
rect	252	249	253	250
rect	253	249	254	250
rect	254	249	255	250
rect	255	249	256	250
rect	256	249	257	250
rect	257	249	258	250
rect	258	249	259	250
rect	259	249	260	250
rect	260	249	261	250
rect	261	249	262	250
rect	262	249	263	250
rect	263	249	264	250
rect	264	249	265	250
rect	265	249	266	250
rect	266	249	267	250
rect	267	249	268	250
rect	268	249	269	250
rect	269	249	270	250
rect	270	249	271	250
rect	271	249	272	250
rect	272	249	273	250
rect	273	249	274	250
rect	274	249	275	250
rect	275	249	276	250
rect	276	249	277	250
rect	277	249	278	250
rect	278	249	279	250
rect	279	249	280	250
rect	280	249	281	250
rect	281	249	282	250
rect	282	249	283	250
rect	283	249	284	250
rect	284	249	285	250
rect	285	249	286	250
rect	286	249	287	250
rect	287	249	288	250
rect	288	249	289	250
rect	289	249	290	250
rect	290	249	291	250
rect	291	249	292	250
rect	292	249	293	250
rect	293	249	294	250
rect	294	249	295	250
rect	295	249	296	250
rect	296	249	297	250
rect	297	249	298	250
rect	298	249	299	250
rect	299	249	300	250
rect	300	249	301	250
rect	301	249	302	250
rect	302	249	303	250
rect	303	249	304	250
rect	304	249	305	250
rect	305	249	306	250
rect	306	249	307	250
rect	307	249	308	250
rect	308	249	309	250
rect	309	249	310	250
rect	310	249	311	250
rect	311	249	312	250
rect	312	249	313	250
rect	313	249	314	250
rect	314	249	315	250
rect	315	249	316	250
rect	317	249	318	250
rect	318	249	319	250
rect	319	249	320	250
rect	320	249	321	250
rect	321	249	322	250
rect	322	249	323	250
rect	323	249	324	250
rect	324	249	325	250
rect	325	249	326	250
rect	326	249	327	250
rect	327	249	328	250
rect	328	249	329	250
rect	329	249	330	250
rect	330	249	331	250
rect	331	249	332	250
rect	332	249	333	250
rect	333	249	334	250
rect	334	249	335	250
rect	335	249	336	250
rect	336	249	337	250
rect	337	249	338	250
rect	338	249	339	250
rect	339	249	340	250
rect	340	249	341	250
rect	341	249	342	250
rect	342	249	343	250
rect	343	249	344	250
rect	344	249	345	250
rect	345	249	346	250
rect	346	249	347	250
rect	347	249	348	250
rect	348	249	349	250
rect	349	249	350	250
rect	350	249	351	250
rect	351	249	352	250
rect	352	249	353	250
rect	353	249	354	250
rect	354	249	355	250
rect	355	249	356	250
rect	356	249	357	250
rect	357	249	358	250
rect	358	249	359	250
rect	359	249	360	250
rect	360	249	361	250
rect	361	249	362	250
rect	362	249	363	250
rect	363	249	364	250
rect	364	249	365	250
rect	366	249	367	250
rect	367	249	368	250
rect	368	249	369	250
rect	369	249	370	250
rect	370	249	371	250
rect	371	249	372	250
rect	372	249	373	250
rect	373	249	374	250
rect	374	249	375	250
rect	375	249	376	250
rect	376	249	377	250
rect	377	249	378	250
rect	378	249	379	250
rect	379	249	380	250
rect	380	249	381	250
rect	0	250	1	251
rect	1	250	2	251
rect	2	250	3	251
rect	3	250	4	251
rect	4	250	5	251
rect	5	250	6	251
rect	7	250	8	251
rect	8	250	9	251
rect	9	250	10	251
rect	10	250	11	251
rect	11	250	12	251
rect	12	250	13	251
rect	14	250	15	251
rect	15	250	16	251
rect	16	250	17	251
rect	17	250	18	251
rect	18	250	19	251
rect	19	250	20	251
rect	20	250	21	251
rect	21	250	22	251
rect	22	250	23	251
rect	23	250	24	251
rect	24	250	25	251
rect	25	250	26	251
rect	26	250	27	251
rect	27	250	28	251
rect	28	250	29	251
rect	29	250	30	251
rect	30	250	31	251
rect	31	250	32	251
rect	32	250	33	251
rect	33	250	34	251
rect	34	250	35	251
rect	35	250	36	251
rect	36	250	37	251
rect	37	250	38	251
rect	38	250	39	251
rect	39	250	40	251
rect	40	250	41	251
rect	41	250	42	251
rect	42	250	43	251
rect	43	250	44	251
rect	44	250	45	251
rect	45	250	46	251
rect	46	250	47	251
rect	47	250	48	251
rect	48	250	49	251
rect	49	250	50	251
rect	50	250	51	251
rect	51	250	52	251
rect	52	250	53	251
rect	53	250	54	251
rect	54	250	55	251
rect	55	250	56	251
rect	56	250	57	251
rect	57	250	58	251
rect	58	250	59	251
rect	59	250	60	251
rect	60	250	61	251
rect	61	250	62	251
rect	62	250	63	251
rect	63	250	64	251
rect	64	250	65	251
rect	65	250	66	251
rect	66	250	67	251
rect	67	250	68	251
rect	69	250	70	251
rect	70	250	71	251
rect	71	250	72	251
rect	72	250	73	251
rect	73	250	74	251
rect	74	250	75	251
rect	76	250	77	251
rect	77	250	78	251
rect	78	250	79	251
rect	79	250	80	251
rect	80	250	81	251
rect	81	250	82	251
rect	82	250	83	251
rect	83	250	84	251
rect	84	250	85	251
rect	85	250	86	251
rect	86	250	87	251
rect	87	250	88	251
rect	88	250	89	251
rect	89	250	90	251
rect	90	250	91	251
rect	92	250	93	251
rect	93	250	94	251
rect	94	250	95	251
rect	95	250	96	251
rect	96	250	97	251
rect	97	250	98	251
rect	99	250	100	251
rect	100	250	101	251
rect	101	250	102	251
rect	102	250	103	251
rect	103	250	104	251
rect	104	250	105	251
rect	105	250	106	251
rect	106	250	107	251
rect	107	250	108	251
rect	108	250	109	251
rect	109	250	110	251
rect	110	250	111	251
rect	111	250	112	251
rect	112	250	113	251
rect	113	250	114	251
rect	114	250	115	251
rect	115	250	116	251
rect	116	250	117	251
rect	117	250	118	251
rect	118	250	119	251
rect	119	250	120	251
rect	120	250	121	251
rect	121	250	122	251
rect	122	250	123	251
rect	123	250	124	251
rect	124	250	125	251
rect	125	250	126	251
rect	127	250	128	251
rect	128	250	129	251
rect	129	250	130	251
rect	130	250	131	251
rect	131	250	132	251
rect	132	250	133	251
rect	133	250	134	251
rect	134	250	135	251
rect	135	250	136	251
rect	136	250	137	251
rect	137	250	138	251
rect	138	250	139	251
rect	139	250	140	251
rect	140	250	141	251
rect	141	250	142	251
rect	142	250	143	251
rect	143	250	144	251
rect	144	250	145	251
rect	145	250	146	251
rect	146	250	147	251
rect	147	250	148	251
rect	148	250	149	251
rect	149	250	150	251
rect	150	250	151	251
rect	151	250	152	251
rect	152	250	153	251
rect	153	250	154	251
rect	154	250	155	251
rect	155	250	156	251
rect	156	250	157	251
rect	157	250	158	251
rect	158	250	159	251
rect	159	250	160	251
rect	160	250	161	251
rect	161	250	162	251
rect	162	250	163	251
rect	163	250	164	251
rect	164	250	165	251
rect	165	250	166	251
rect	166	250	167	251
rect	167	250	168	251
rect	168	250	169	251
rect	169	250	170	251
rect	170	250	171	251
rect	171	250	172	251
rect	172	250	173	251
rect	173	250	174	251
rect	174	250	175	251
rect	175	250	176	251
rect	176	250	177	251
rect	177	250	178	251
rect	178	250	179	251
rect	179	250	180	251
rect	180	250	181	251
rect	181	250	182	251
rect	182	250	183	251
rect	183	250	184	251
rect	184	250	185	251
rect	185	250	186	251
rect	186	250	187	251
rect	187	250	188	251
rect	188	250	189	251
rect	189	250	190	251
rect	190	250	191	251
rect	191	250	192	251
rect	192	250	193	251
rect	193	250	194	251
rect	194	250	195	251
rect	195	250	196	251
rect	196	250	197	251
rect	197	250	198	251
rect	198	250	199	251
rect	199	250	200	251
rect	200	250	201	251
rect	201	250	202	251
rect	202	250	203	251
rect	203	250	204	251
rect	204	250	205	251
rect	206	250	207	251
rect	207	250	208	251
rect	208	250	209	251
rect	209	250	210	251
rect	210	250	211	251
rect	211	250	212	251
rect	213	250	214	251
rect	214	250	215	251
rect	215	250	216	251
rect	216	250	217	251
rect	217	250	218	251
rect	218	250	219	251
rect	219	250	220	251
rect	220	250	221	251
rect	221	250	222	251
rect	222	250	223	251
rect	223	250	224	251
rect	224	250	225	251
rect	225	250	226	251
rect	226	250	227	251
rect	227	250	228	251
rect	228	250	229	251
rect	229	250	230	251
rect	230	250	231	251
rect	231	250	232	251
rect	232	250	233	251
rect	233	250	234	251
rect	234	250	235	251
rect	235	250	236	251
rect	236	250	237	251
rect	237	250	238	251
rect	238	250	239	251
rect	239	250	240	251
rect	241	250	242	251
rect	242	250	243	251
rect	243	250	244	251
rect	244	250	245	251
rect	245	250	246	251
rect	246	250	247	251
rect	247	250	248	251
rect	248	250	249	251
rect	249	250	250	251
rect	250	250	251	251
rect	251	250	252	251
rect	252	250	253	251
rect	253	250	254	251
rect	254	250	255	251
rect	255	250	256	251
rect	256	250	257	251
rect	257	250	258	251
rect	258	250	259	251
rect	259	250	260	251
rect	260	250	261	251
rect	261	250	262	251
rect	262	250	263	251
rect	263	250	264	251
rect	264	250	265	251
rect	265	250	266	251
rect	266	250	267	251
rect	267	250	268	251
rect	268	250	269	251
rect	269	250	270	251
rect	270	250	271	251
rect	271	250	272	251
rect	272	250	273	251
rect	273	250	274	251
rect	274	250	275	251
rect	275	250	276	251
rect	276	250	277	251
rect	277	250	278	251
rect	278	250	279	251
rect	279	250	280	251
rect	280	250	281	251
rect	281	250	282	251
rect	282	250	283	251
rect	283	250	284	251
rect	284	250	285	251
rect	285	250	286	251
rect	286	250	287	251
rect	287	250	288	251
rect	288	250	289	251
rect	289	250	290	251
rect	290	250	291	251
rect	291	250	292	251
rect	292	250	293	251
rect	293	250	294	251
rect	294	250	295	251
rect	295	250	296	251
rect	296	250	297	251
rect	297	250	298	251
rect	298	250	299	251
rect	299	250	300	251
rect	300	250	301	251
rect	301	250	302	251
rect	302	250	303	251
rect	303	250	304	251
rect	304	250	305	251
rect	305	250	306	251
rect	306	250	307	251
rect	307	250	308	251
rect	308	250	309	251
rect	309	250	310	251
rect	310	250	311	251
rect	311	250	312	251
rect	312	250	313	251
rect	313	250	314	251
rect	314	250	315	251
rect	315	250	316	251
rect	317	250	318	251
rect	318	250	319	251
rect	319	250	320	251
rect	320	250	321	251
rect	321	250	322	251
rect	322	250	323	251
rect	323	250	324	251
rect	324	250	325	251
rect	325	250	326	251
rect	326	250	327	251
rect	327	250	328	251
rect	328	250	329	251
rect	329	250	330	251
rect	330	250	331	251
rect	331	250	332	251
rect	332	250	333	251
rect	333	250	334	251
rect	334	250	335	251
rect	335	250	336	251
rect	336	250	337	251
rect	337	250	338	251
rect	338	250	339	251
rect	339	250	340	251
rect	340	250	341	251
rect	341	250	342	251
rect	342	250	343	251
rect	343	250	344	251
rect	344	250	345	251
rect	345	250	346	251
rect	346	250	347	251
rect	347	250	348	251
rect	348	250	349	251
rect	349	250	350	251
rect	350	250	351	251
rect	351	250	352	251
rect	352	250	353	251
rect	353	250	354	251
rect	354	250	355	251
rect	355	250	356	251
rect	356	250	357	251
rect	357	250	358	251
rect	358	250	359	251
rect	359	250	360	251
rect	360	250	361	251
rect	361	250	362	251
rect	362	250	363	251
rect	363	250	364	251
rect	364	250	365	251
rect	366	250	367	251
rect	367	250	368	251
rect	368	250	369	251
rect	369	250	370	251
rect	370	250	371	251
rect	371	250	372	251
rect	372	250	373	251
rect	373	250	374	251
rect	374	250	375	251
rect	375	250	376	251
rect	376	250	377	251
rect	377	250	378	251
rect	378	250	379	251
rect	379	250	380	251
rect	380	250	381	251
rect	0	251	1	252
rect	1	251	2	252
rect	2	251	3	252
rect	3	251	4	252
rect	4	251	5	252
rect	5	251	6	252
rect	7	251	8	252
rect	8	251	9	252
rect	9	251	10	252
rect	10	251	11	252
rect	11	251	12	252
rect	12	251	13	252
rect	14	251	15	252
rect	15	251	16	252
rect	16	251	17	252
rect	17	251	18	252
rect	18	251	19	252
rect	19	251	20	252
rect	20	251	21	252
rect	21	251	22	252
rect	22	251	23	252
rect	23	251	24	252
rect	24	251	25	252
rect	25	251	26	252
rect	26	251	27	252
rect	27	251	28	252
rect	28	251	29	252
rect	29	251	30	252
rect	30	251	31	252
rect	31	251	32	252
rect	32	251	33	252
rect	33	251	34	252
rect	34	251	35	252
rect	35	251	36	252
rect	36	251	37	252
rect	37	251	38	252
rect	38	251	39	252
rect	39	251	40	252
rect	40	251	41	252
rect	41	251	42	252
rect	42	251	43	252
rect	43	251	44	252
rect	44	251	45	252
rect	45	251	46	252
rect	46	251	47	252
rect	47	251	48	252
rect	48	251	49	252
rect	49	251	50	252
rect	50	251	51	252
rect	51	251	52	252
rect	52	251	53	252
rect	53	251	54	252
rect	54	251	55	252
rect	55	251	56	252
rect	56	251	57	252
rect	57	251	58	252
rect	58	251	59	252
rect	59	251	60	252
rect	60	251	61	252
rect	61	251	62	252
rect	62	251	63	252
rect	63	251	64	252
rect	64	251	65	252
rect	65	251	66	252
rect	66	251	67	252
rect	67	251	68	252
rect	69	251	70	252
rect	70	251	71	252
rect	71	251	72	252
rect	72	251	73	252
rect	73	251	74	252
rect	74	251	75	252
rect	76	251	77	252
rect	77	251	78	252
rect	78	251	79	252
rect	79	251	80	252
rect	80	251	81	252
rect	81	251	82	252
rect	82	251	83	252
rect	83	251	84	252
rect	84	251	85	252
rect	85	251	86	252
rect	86	251	87	252
rect	87	251	88	252
rect	88	251	89	252
rect	89	251	90	252
rect	90	251	91	252
rect	92	251	93	252
rect	93	251	94	252
rect	94	251	95	252
rect	95	251	96	252
rect	96	251	97	252
rect	97	251	98	252
rect	99	251	100	252
rect	100	251	101	252
rect	101	251	102	252
rect	102	251	103	252
rect	103	251	104	252
rect	104	251	105	252
rect	105	251	106	252
rect	106	251	107	252
rect	107	251	108	252
rect	108	251	109	252
rect	109	251	110	252
rect	110	251	111	252
rect	111	251	112	252
rect	112	251	113	252
rect	113	251	114	252
rect	114	251	115	252
rect	115	251	116	252
rect	116	251	117	252
rect	117	251	118	252
rect	118	251	119	252
rect	119	251	120	252
rect	120	251	121	252
rect	121	251	122	252
rect	122	251	123	252
rect	123	251	124	252
rect	124	251	125	252
rect	125	251	126	252
rect	127	251	128	252
rect	128	251	129	252
rect	129	251	130	252
rect	130	251	131	252
rect	131	251	132	252
rect	132	251	133	252
rect	133	251	134	252
rect	134	251	135	252
rect	135	251	136	252
rect	136	251	137	252
rect	137	251	138	252
rect	138	251	139	252
rect	139	251	140	252
rect	140	251	141	252
rect	141	251	142	252
rect	142	251	143	252
rect	143	251	144	252
rect	144	251	145	252
rect	145	251	146	252
rect	146	251	147	252
rect	147	251	148	252
rect	148	251	149	252
rect	149	251	150	252
rect	150	251	151	252
rect	151	251	152	252
rect	152	251	153	252
rect	153	251	154	252
rect	154	251	155	252
rect	155	251	156	252
rect	156	251	157	252
rect	157	251	158	252
rect	158	251	159	252
rect	159	251	160	252
rect	160	251	161	252
rect	161	251	162	252
rect	162	251	163	252
rect	163	251	164	252
rect	164	251	165	252
rect	165	251	166	252
rect	166	251	167	252
rect	167	251	168	252
rect	168	251	169	252
rect	169	251	170	252
rect	170	251	171	252
rect	171	251	172	252
rect	172	251	173	252
rect	173	251	174	252
rect	174	251	175	252
rect	175	251	176	252
rect	176	251	177	252
rect	177	251	178	252
rect	178	251	179	252
rect	179	251	180	252
rect	180	251	181	252
rect	181	251	182	252
rect	182	251	183	252
rect	183	251	184	252
rect	184	251	185	252
rect	185	251	186	252
rect	186	251	187	252
rect	187	251	188	252
rect	188	251	189	252
rect	189	251	190	252
rect	190	251	191	252
rect	191	251	192	252
rect	192	251	193	252
rect	193	251	194	252
rect	194	251	195	252
rect	195	251	196	252
rect	196	251	197	252
rect	197	251	198	252
rect	198	251	199	252
rect	199	251	200	252
rect	200	251	201	252
rect	201	251	202	252
rect	202	251	203	252
rect	203	251	204	252
rect	204	251	205	252
rect	206	251	207	252
rect	207	251	208	252
rect	208	251	209	252
rect	209	251	210	252
rect	210	251	211	252
rect	211	251	212	252
rect	213	251	214	252
rect	214	251	215	252
rect	215	251	216	252
rect	216	251	217	252
rect	217	251	218	252
rect	218	251	219	252
rect	219	251	220	252
rect	220	251	221	252
rect	221	251	222	252
rect	222	251	223	252
rect	223	251	224	252
rect	224	251	225	252
rect	225	251	226	252
rect	226	251	227	252
rect	227	251	228	252
rect	228	251	229	252
rect	229	251	230	252
rect	230	251	231	252
rect	231	251	232	252
rect	232	251	233	252
rect	233	251	234	252
rect	234	251	235	252
rect	235	251	236	252
rect	236	251	237	252
rect	237	251	238	252
rect	238	251	239	252
rect	239	251	240	252
rect	241	251	242	252
rect	242	251	243	252
rect	243	251	244	252
rect	244	251	245	252
rect	245	251	246	252
rect	246	251	247	252
rect	247	251	248	252
rect	248	251	249	252
rect	249	251	250	252
rect	250	251	251	252
rect	251	251	252	252
rect	252	251	253	252
rect	253	251	254	252
rect	254	251	255	252
rect	255	251	256	252
rect	256	251	257	252
rect	257	251	258	252
rect	258	251	259	252
rect	259	251	260	252
rect	260	251	261	252
rect	261	251	262	252
rect	262	251	263	252
rect	263	251	264	252
rect	264	251	265	252
rect	265	251	266	252
rect	266	251	267	252
rect	267	251	268	252
rect	268	251	269	252
rect	269	251	270	252
rect	270	251	271	252
rect	271	251	272	252
rect	272	251	273	252
rect	273	251	274	252
rect	274	251	275	252
rect	275	251	276	252
rect	276	251	277	252
rect	277	251	278	252
rect	278	251	279	252
rect	279	251	280	252
rect	280	251	281	252
rect	281	251	282	252
rect	282	251	283	252
rect	283	251	284	252
rect	284	251	285	252
rect	285	251	286	252
rect	286	251	287	252
rect	287	251	288	252
rect	288	251	289	252
rect	289	251	290	252
rect	290	251	291	252
rect	291	251	292	252
rect	292	251	293	252
rect	293	251	294	252
rect	294	251	295	252
rect	295	251	296	252
rect	296	251	297	252
rect	297	251	298	252
rect	298	251	299	252
rect	299	251	300	252
rect	300	251	301	252
rect	301	251	302	252
rect	302	251	303	252
rect	303	251	304	252
rect	304	251	305	252
rect	305	251	306	252
rect	306	251	307	252
rect	307	251	308	252
rect	308	251	309	252
rect	309	251	310	252
rect	310	251	311	252
rect	311	251	312	252
rect	312	251	313	252
rect	313	251	314	252
rect	314	251	315	252
rect	315	251	316	252
rect	317	251	318	252
rect	318	251	319	252
rect	319	251	320	252
rect	320	251	321	252
rect	321	251	322	252
rect	322	251	323	252
rect	323	251	324	252
rect	324	251	325	252
rect	325	251	326	252
rect	326	251	327	252
rect	327	251	328	252
rect	328	251	329	252
rect	329	251	330	252
rect	330	251	331	252
rect	331	251	332	252
rect	332	251	333	252
rect	333	251	334	252
rect	334	251	335	252
rect	335	251	336	252
rect	336	251	337	252
rect	337	251	338	252
rect	338	251	339	252
rect	339	251	340	252
rect	340	251	341	252
rect	341	251	342	252
rect	342	251	343	252
rect	343	251	344	252
rect	344	251	345	252
rect	345	251	346	252
rect	346	251	347	252
rect	347	251	348	252
rect	348	251	349	252
rect	349	251	350	252
rect	350	251	351	252
rect	351	251	352	252
rect	352	251	353	252
rect	353	251	354	252
rect	354	251	355	252
rect	355	251	356	252
rect	356	251	357	252
rect	357	251	358	252
rect	358	251	359	252
rect	359	251	360	252
rect	360	251	361	252
rect	361	251	362	252
rect	362	251	363	252
rect	363	251	364	252
rect	364	251	365	252
rect	366	251	367	252
rect	367	251	368	252
rect	368	251	369	252
rect	369	251	370	252
rect	370	251	371	252
rect	371	251	372	252
rect	372	251	373	252
rect	373	251	374	252
rect	374	251	375	252
rect	375	251	376	252
rect	376	251	377	252
rect	377	251	378	252
rect	378	251	379	252
rect	379	251	380	252
rect	380	251	381	252
rect	0	252	1	253
rect	1	252	2	253
rect	2	252	3	253
rect	3	252	4	253
rect	4	252	5	253
rect	5	252	6	253
rect	7	252	8	253
rect	8	252	9	253
rect	9	252	10	253
rect	10	252	11	253
rect	11	252	12	253
rect	12	252	13	253
rect	14	252	15	253
rect	15	252	16	253
rect	16	252	17	253
rect	17	252	18	253
rect	18	252	19	253
rect	19	252	20	253
rect	20	252	21	253
rect	21	252	22	253
rect	22	252	23	253
rect	23	252	24	253
rect	24	252	25	253
rect	25	252	26	253
rect	26	252	27	253
rect	27	252	28	253
rect	28	252	29	253
rect	29	252	30	253
rect	30	252	31	253
rect	31	252	32	253
rect	32	252	33	253
rect	33	252	34	253
rect	34	252	35	253
rect	35	252	36	253
rect	36	252	37	253
rect	37	252	38	253
rect	38	252	39	253
rect	39	252	40	253
rect	40	252	41	253
rect	41	252	42	253
rect	42	252	43	253
rect	43	252	44	253
rect	44	252	45	253
rect	45	252	46	253
rect	46	252	47	253
rect	47	252	48	253
rect	48	252	49	253
rect	49	252	50	253
rect	50	252	51	253
rect	51	252	52	253
rect	52	252	53	253
rect	53	252	54	253
rect	54	252	55	253
rect	55	252	56	253
rect	56	252	57	253
rect	57	252	58	253
rect	58	252	59	253
rect	59	252	60	253
rect	60	252	61	253
rect	61	252	62	253
rect	62	252	63	253
rect	63	252	64	253
rect	64	252	65	253
rect	65	252	66	253
rect	66	252	67	253
rect	67	252	68	253
rect	69	252	70	253
rect	70	252	71	253
rect	71	252	72	253
rect	72	252	73	253
rect	73	252	74	253
rect	74	252	75	253
rect	76	252	77	253
rect	77	252	78	253
rect	78	252	79	253
rect	79	252	80	253
rect	80	252	81	253
rect	81	252	82	253
rect	82	252	83	253
rect	83	252	84	253
rect	84	252	85	253
rect	85	252	86	253
rect	86	252	87	253
rect	87	252	88	253
rect	88	252	89	253
rect	89	252	90	253
rect	90	252	91	253
rect	92	252	93	253
rect	93	252	94	253
rect	94	252	95	253
rect	95	252	96	253
rect	96	252	97	253
rect	97	252	98	253
rect	99	252	100	253
rect	100	252	101	253
rect	101	252	102	253
rect	102	252	103	253
rect	103	252	104	253
rect	104	252	105	253
rect	105	252	106	253
rect	106	252	107	253
rect	107	252	108	253
rect	108	252	109	253
rect	109	252	110	253
rect	110	252	111	253
rect	111	252	112	253
rect	112	252	113	253
rect	113	252	114	253
rect	114	252	115	253
rect	115	252	116	253
rect	116	252	117	253
rect	117	252	118	253
rect	118	252	119	253
rect	119	252	120	253
rect	120	252	121	253
rect	121	252	122	253
rect	122	252	123	253
rect	123	252	124	253
rect	124	252	125	253
rect	125	252	126	253
rect	127	252	128	253
rect	128	252	129	253
rect	129	252	130	253
rect	130	252	131	253
rect	131	252	132	253
rect	132	252	133	253
rect	133	252	134	253
rect	134	252	135	253
rect	135	252	136	253
rect	136	252	137	253
rect	137	252	138	253
rect	138	252	139	253
rect	139	252	140	253
rect	140	252	141	253
rect	141	252	142	253
rect	142	252	143	253
rect	143	252	144	253
rect	144	252	145	253
rect	145	252	146	253
rect	146	252	147	253
rect	147	252	148	253
rect	148	252	149	253
rect	149	252	150	253
rect	150	252	151	253
rect	151	252	152	253
rect	152	252	153	253
rect	153	252	154	253
rect	154	252	155	253
rect	155	252	156	253
rect	156	252	157	253
rect	157	252	158	253
rect	158	252	159	253
rect	159	252	160	253
rect	160	252	161	253
rect	161	252	162	253
rect	162	252	163	253
rect	163	252	164	253
rect	164	252	165	253
rect	165	252	166	253
rect	166	252	167	253
rect	167	252	168	253
rect	168	252	169	253
rect	169	252	170	253
rect	170	252	171	253
rect	171	252	172	253
rect	172	252	173	253
rect	173	252	174	253
rect	174	252	175	253
rect	175	252	176	253
rect	176	252	177	253
rect	177	252	178	253
rect	178	252	179	253
rect	179	252	180	253
rect	180	252	181	253
rect	181	252	182	253
rect	182	252	183	253
rect	183	252	184	253
rect	184	252	185	253
rect	185	252	186	253
rect	186	252	187	253
rect	187	252	188	253
rect	188	252	189	253
rect	189	252	190	253
rect	190	252	191	253
rect	191	252	192	253
rect	192	252	193	253
rect	193	252	194	253
rect	194	252	195	253
rect	195	252	196	253
rect	196	252	197	253
rect	197	252	198	253
rect	198	252	199	253
rect	199	252	200	253
rect	200	252	201	253
rect	201	252	202	253
rect	202	252	203	253
rect	203	252	204	253
rect	204	252	205	253
rect	206	252	207	253
rect	207	252	208	253
rect	208	252	209	253
rect	209	252	210	253
rect	210	252	211	253
rect	211	252	212	253
rect	213	252	214	253
rect	214	252	215	253
rect	215	252	216	253
rect	216	252	217	253
rect	217	252	218	253
rect	218	252	219	253
rect	219	252	220	253
rect	220	252	221	253
rect	221	252	222	253
rect	222	252	223	253
rect	223	252	224	253
rect	224	252	225	253
rect	225	252	226	253
rect	226	252	227	253
rect	227	252	228	253
rect	228	252	229	253
rect	229	252	230	253
rect	230	252	231	253
rect	231	252	232	253
rect	232	252	233	253
rect	233	252	234	253
rect	234	252	235	253
rect	235	252	236	253
rect	236	252	237	253
rect	237	252	238	253
rect	238	252	239	253
rect	239	252	240	253
rect	241	252	242	253
rect	242	252	243	253
rect	243	252	244	253
rect	244	252	245	253
rect	245	252	246	253
rect	246	252	247	253
rect	247	252	248	253
rect	248	252	249	253
rect	249	252	250	253
rect	250	252	251	253
rect	251	252	252	253
rect	252	252	253	253
rect	253	252	254	253
rect	254	252	255	253
rect	255	252	256	253
rect	256	252	257	253
rect	257	252	258	253
rect	258	252	259	253
rect	259	252	260	253
rect	260	252	261	253
rect	261	252	262	253
rect	262	252	263	253
rect	263	252	264	253
rect	264	252	265	253
rect	265	252	266	253
rect	266	252	267	253
rect	267	252	268	253
rect	268	252	269	253
rect	269	252	270	253
rect	270	252	271	253
rect	271	252	272	253
rect	272	252	273	253
rect	273	252	274	253
rect	274	252	275	253
rect	275	252	276	253
rect	276	252	277	253
rect	277	252	278	253
rect	278	252	279	253
rect	279	252	280	253
rect	280	252	281	253
rect	281	252	282	253
rect	282	252	283	253
rect	283	252	284	253
rect	284	252	285	253
rect	285	252	286	253
rect	286	252	287	253
rect	287	252	288	253
rect	288	252	289	253
rect	289	252	290	253
rect	290	252	291	253
rect	291	252	292	253
rect	292	252	293	253
rect	293	252	294	253
rect	294	252	295	253
rect	295	252	296	253
rect	296	252	297	253
rect	297	252	298	253
rect	298	252	299	253
rect	299	252	300	253
rect	300	252	301	253
rect	301	252	302	253
rect	302	252	303	253
rect	303	252	304	253
rect	304	252	305	253
rect	305	252	306	253
rect	306	252	307	253
rect	307	252	308	253
rect	308	252	309	253
rect	309	252	310	253
rect	310	252	311	253
rect	311	252	312	253
rect	312	252	313	253
rect	313	252	314	253
rect	314	252	315	253
rect	315	252	316	253
rect	317	252	318	253
rect	318	252	319	253
rect	319	252	320	253
rect	320	252	321	253
rect	321	252	322	253
rect	322	252	323	253
rect	323	252	324	253
rect	324	252	325	253
rect	325	252	326	253
rect	326	252	327	253
rect	327	252	328	253
rect	328	252	329	253
rect	329	252	330	253
rect	330	252	331	253
rect	331	252	332	253
rect	332	252	333	253
rect	333	252	334	253
rect	334	252	335	253
rect	335	252	336	253
rect	336	252	337	253
rect	337	252	338	253
rect	338	252	339	253
rect	339	252	340	253
rect	340	252	341	253
rect	341	252	342	253
rect	342	252	343	253
rect	343	252	344	253
rect	344	252	345	253
rect	345	252	346	253
rect	346	252	347	253
rect	347	252	348	253
rect	348	252	349	253
rect	349	252	350	253
rect	350	252	351	253
rect	351	252	352	253
rect	352	252	353	253
rect	353	252	354	253
rect	354	252	355	253
rect	355	252	356	253
rect	356	252	357	253
rect	357	252	358	253
rect	358	252	359	253
rect	359	252	360	253
rect	360	252	361	253
rect	361	252	362	253
rect	362	252	363	253
rect	363	252	364	253
rect	364	252	365	253
rect	366	252	367	253
rect	367	252	368	253
rect	368	252	369	253
rect	369	252	370	253
rect	370	252	371	253
rect	371	252	372	253
rect	372	252	373	253
rect	373	252	374	253
rect	374	252	375	253
rect	375	252	376	253
rect	376	252	377	253
rect	377	252	378	253
rect	378	252	379	253
rect	379	252	380	253
rect	380	252	381	253
rect	0	253	1	254
rect	1	253	2	254
rect	2	253	3	254
rect	3	253	4	254
rect	4	253	5	254
rect	5	253	6	254
rect	7	253	8	254
rect	8	253	9	254
rect	9	253	10	254
rect	10	253	11	254
rect	11	253	12	254
rect	12	253	13	254
rect	14	253	15	254
rect	15	253	16	254
rect	16	253	17	254
rect	17	253	18	254
rect	18	253	19	254
rect	19	253	20	254
rect	20	253	21	254
rect	21	253	22	254
rect	22	253	23	254
rect	23	253	24	254
rect	24	253	25	254
rect	25	253	26	254
rect	26	253	27	254
rect	27	253	28	254
rect	28	253	29	254
rect	29	253	30	254
rect	30	253	31	254
rect	31	253	32	254
rect	32	253	33	254
rect	33	253	34	254
rect	34	253	35	254
rect	35	253	36	254
rect	36	253	37	254
rect	37	253	38	254
rect	38	253	39	254
rect	39	253	40	254
rect	40	253	41	254
rect	41	253	42	254
rect	42	253	43	254
rect	43	253	44	254
rect	44	253	45	254
rect	45	253	46	254
rect	46	253	47	254
rect	47	253	48	254
rect	48	253	49	254
rect	49	253	50	254
rect	50	253	51	254
rect	51	253	52	254
rect	52	253	53	254
rect	53	253	54	254
rect	54	253	55	254
rect	55	253	56	254
rect	56	253	57	254
rect	57	253	58	254
rect	58	253	59	254
rect	59	253	60	254
rect	60	253	61	254
rect	61	253	62	254
rect	62	253	63	254
rect	63	253	64	254
rect	64	253	65	254
rect	65	253	66	254
rect	66	253	67	254
rect	67	253	68	254
rect	69	253	70	254
rect	70	253	71	254
rect	71	253	72	254
rect	72	253	73	254
rect	73	253	74	254
rect	74	253	75	254
rect	76	253	77	254
rect	77	253	78	254
rect	78	253	79	254
rect	79	253	80	254
rect	80	253	81	254
rect	81	253	82	254
rect	82	253	83	254
rect	83	253	84	254
rect	84	253	85	254
rect	85	253	86	254
rect	86	253	87	254
rect	87	253	88	254
rect	88	253	89	254
rect	89	253	90	254
rect	90	253	91	254
rect	92	253	93	254
rect	93	253	94	254
rect	94	253	95	254
rect	95	253	96	254
rect	96	253	97	254
rect	97	253	98	254
rect	99	253	100	254
rect	100	253	101	254
rect	101	253	102	254
rect	102	253	103	254
rect	103	253	104	254
rect	104	253	105	254
rect	105	253	106	254
rect	106	253	107	254
rect	107	253	108	254
rect	108	253	109	254
rect	109	253	110	254
rect	110	253	111	254
rect	111	253	112	254
rect	112	253	113	254
rect	113	253	114	254
rect	114	253	115	254
rect	115	253	116	254
rect	116	253	117	254
rect	117	253	118	254
rect	118	253	119	254
rect	119	253	120	254
rect	120	253	121	254
rect	121	253	122	254
rect	122	253	123	254
rect	123	253	124	254
rect	124	253	125	254
rect	125	253	126	254
rect	127	253	128	254
rect	128	253	129	254
rect	129	253	130	254
rect	130	253	131	254
rect	131	253	132	254
rect	132	253	133	254
rect	133	253	134	254
rect	134	253	135	254
rect	135	253	136	254
rect	136	253	137	254
rect	137	253	138	254
rect	138	253	139	254
rect	139	253	140	254
rect	140	253	141	254
rect	141	253	142	254
rect	142	253	143	254
rect	143	253	144	254
rect	144	253	145	254
rect	145	253	146	254
rect	146	253	147	254
rect	147	253	148	254
rect	148	253	149	254
rect	149	253	150	254
rect	150	253	151	254
rect	151	253	152	254
rect	152	253	153	254
rect	153	253	154	254
rect	154	253	155	254
rect	155	253	156	254
rect	156	253	157	254
rect	157	253	158	254
rect	158	253	159	254
rect	159	253	160	254
rect	160	253	161	254
rect	161	253	162	254
rect	162	253	163	254
rect	163	253	164	254
rect	164	253	165	254
rect	165	253	166	254
rect	166	253	167	254
rect	167	253	168	254
rect	168	253	169	254
rect	169	253	170	254
rect	170	253	171	254
rect	171	253	172	254
rect	172	253	173	254
rect	173	253	174	254
rect	174	253	175	254
rect	175	253	176	254
rect	176	253	177	254
rect	177	253	178	254
rect	178	253	179	254
rect	179	253	180	254
rect	180	253	181	254
rect	181	253	182	254
rect	182	253	183	254
rect	183	253	184	254
rect	184	253	185	254
rect	185	253	186	254
rect	186	253	187	254
rect	187	253	188	254
rect	188	253	189	254
rect	189	253	190	254
rect	190	253	191	254
rect	191	253	192	254
rect	192	253	193	254
rect	193	253	194	254
rect	194	253	195	254
rect	195	253	196	254
rect	196	253	197	254
rect	197	253	198	254
rect	198	253	199	254
rect	199	253	200	254
rect	200	253	201	254
rect	201	253	202	254
rect	202	253	203	254
rect	203	253	204	254
rect	204	253	205	254
rect	206	253	207	254
rect	207	253	208	254
rect	208	253	209	254
rect	209	253	210	254
rect	210	253	211	254
rect	211	253	212	254
rect	213	253	214	254
rect	214	253	215	254
rect	215	253	216	254
rect	216	253	217	254
rect	217	253	218	254
rect	218	253	219	254
rect	219	253	220	254
rect	220	253	221	254
rect	221	253	222	254
rect	222	253	223	254
rect	223	253	224	254
rect	224	253	225	254
rect	225	253	226	254
rect	226	253	227	254
rect	227	253	228	254
rect	228	253	229	254
rect	229	253	230	254
rect	230	253	231	254
rect	231	253	232	254
rect	232	253	233	254
rect	233	253	234	254
rect	234	253	235	254
rect	235	253	236	254
rect	236	253	237	254
rect	237	253	238	254
rect	238	253	239	254
rect	239	253	240	254
rect	241	253	242	254
rect	242	253	243	254
rect	243	253	244	254
rect	244	253	245	254
rect	245	253	246	254
rect	246	253	247	254
rect	247	253	248	254
rect	248	253	249	254
rect	249	253	250	254
rect	250	253	251	254
rect	251	253	252	254
rect	252	253	253	254
rect	253	253	254	254
rect	254	253	255	254
rect	255	253	256	254
rect	256	253	257	254
rect	257	253	258	254
rect	258	253	259	254
rect	259	253	260	254
rect	260	253	261	254
rect	261	253	262	254
rect	262	253	263	254
rect	263	253	264	254
rect	264	253	265	254
rect	265	253	266	254
rect	266	253	267	254
rect	267	253	268	254
rect	268	253	269	254
rect	269	253	270	254
rect	270	253	271	254
rect	271	253	272	254
rect	272	253	273	254
rect	273	253	274	254
rect	274	253	275	254
rect	275	253	276	254
rect	276	253	277	254
rect	277	253	278	254
rect	278	253	279	254
rect	279	253	280	254
rect	280	253	281	254
rect	281	253	282	254
rect	282	253	283	254
rect	283	253	284	254
rect	284	253	285	254
rect	285	253	286	254
rect	286	253	287	254
rect	287	253	288	254
rect	288	253	289	254
rect	289	253	290	254
rect	290	253	291	254
rect	291	253	292	254
rect	292	253	293	254
rect	293	253	294	254
rect	294	253	295	254
rect	295	253	296	254
rect	296	253	297	254
rect	297	253	298	254
rect	298	253	299	254
rect	299	253	300	254
rect	300	253	301	254
rect	301	253	302	254
rect	302	253	303	254
rect	303	253	304	254
rect	304	253	305	254
rect	305	253	306	254
rect	306	253	307	254
rect	307	253	308	254
rect	308	253	309	254
rect	309	253	310	254
rect	310	253	311	254
rect	311	253	312	254
rect	312	253	313	254
rect	313	253	314	254
rect	314	253	315	254
rect	315	253	316	254
rect	317	253	318	254
rect	318	253	319	254
rect	319	253	320	254
rect	320	253	321	254
rect	321	253	322	254
rect	322	253	323	254
rect	323	253	324	254
rect	324	253	325	254
rect	325	253	326	254
rect	326	253	327	254
rect	327	253	328	254
rect	328	253	329	254
rect	329	253	330	254
rect	330	253	331	254
rect	331	253	332	254
rect	332	253	333	254
rect	333	253	334	254
rect	334	253	335	254
rect	335	253	336	254
rect	336	253	337	254
rect	337	253	338	254
rect	338	253	339	254
rect	339	253	340	254
rect	340	253	341	254
rect	341	253	342	254
rect	342	253	343	254
rect	343	253	344	254
rect	344	253	345	254
rect	345	253	346	254
rect	346	253	347	254
rect	347	253	348	254
rect	348	253	349	254
rect	349	253	350	254
rect	350	253	351	254
rect	351	253	352	254
rect	352	253	353	254
rect	353	253	354	254
rect	354	253	355	254
rect	355	253	356	254
rect	356	253	357	254
rect	357	253	358	254
rect	358	253	359	254
rect	359	253	360	254
rect	360	253	361	254
rect	361	253	362	254
rect	362	253	363	254
rect	363	253	364	254
rect	364	253	365	254
rect	366	253	367	254
rect	367	253	368	254
rect	368	253	369	254
rect	369	253	370	254
rect	370	253	371	254
rect	371	253	372	254
rect	372	253	373	254
rect	373	253	374	254
rect	374	253	375	254
rect	375	253	376	254
rect	376	253	377	254
rect	377	253	378	254
rect	378	253	379	254
rect	379	253	380	254
rect	380	253	381	254
rect	0	269	1	270
rect	1	269	2	270
rect	2	269	3	270
rect	3	269	4	270
rect	4	269	5	270
rect	5	269	6	270
rect	7	269	8	270
rect	8	269	9	270
rect	9	269	10	270
rect	10	269	11	270
rect	11	269	12	270
rect	12	269	13	270
rect	14	269	15	270
rect	15	269	16	270
rect	16	269	17	270
rect	17	269	18	270
rect	18	269	19	270
rect	19	269	20	270
rect	20	269	21	270
rect	21	269	22	270
rect	22	269	23	270
rect	23	269	24	270
rect	24	269	25	270
rect	25	269	26	270
rect	26	269	27	270
rect	27	269	28	270
rect	28	269	29	270
rect	29	269	30	270
rect	30	269	31	270
rect	31	269	32	270
rect	32	269	33	270
rect	33	269	34	270
rect	34	269	35	270
rect	35	269	36	270
rect	36	269	37	270
rect	37	269	38	270
rect	38	269	39	270
rect	39	269	40	270
rect	40	269	41	270
rect	41	269	42	270
rect	42	269	43	270
rect	43	269	44	270
rect	44	269	45	270
rect	45	269	46	270
rect	46	269	47	270
rect	47	269	48	270
rect	48	269	49	270
rect	49	269	50	270
rect	50	269	51	270
rect	51	269	52	270
rect	52	269	53	270
rect	53	269	54	270
rect	54	269	55	270
rect	55	269	56	270
rect	56	269	57	270
rect	57	269	58	270
rect	58	269	59	270
rect	59	269	60	270
rect	60	269	61	270
rect	61	269	62	270
rect	62	269	63	270
rect	63	269	64	270
rect	64	269	65	270
rect	65	269	66	270
rect	66	269	67	270
rect	67	269	68	270
rect	68	269	69	270
rect	69	269	70	270
rect	70	269	71	270
rect	71	269	72	270
rect	72	269	73	270
rect	73	269	74	270
rect	74	269	75	270
rect	75	269	76	270
rect	76	269	77	270
rect	77	269	78	270
rect	78	269	79	270
rect	79	269	80	270
rect	80	269	81	270
rect	81	269	82	270
rect	82	269	83	270
rect	84	269	85	270
rect	85	269	86	270
rect	86	269	87	270
rect	87	269	88	270
rect	88	269	89	270
rect	89	269	90	270
rect	90	269	91	270
rect	91	269	92	270
rect	92	269	93	270
rect	93	269	94	270
rect	94	269	95	270
rect	95	269	96	270
rect	96	269	97	270
rect	97	269	98	270
rect	98	269	99	270
rect	99	269	100	270
rect	100	269	101	270
rect	101	269	102	270
rect	102	269	103	270
rect	103	269	104	270
rect	104	269	105	270
rect	105	269	106	270
rect	106	269	107	270
rect	107	269	108	270
rect	108	269	109	270
rect	109	269	110	270
rect	110	269	111	270
rect	111	269	112	270
rect	112	269	113	270
rect	113	269	114	270
rect	114	269	115	270
rect	115	269	116	270
rect	116	269	117	270
rect	117	269	118	270
rect	118	269	119	270
rect	119	269	120	270
rect	120	269	121	270
rect	121	269	122	270
rect	122	269	123	270
rect	123	269	124	270
rect	124	269	125	270
rect	125	269	126	270
rect	126	269	127	270
rect	127	269	128	270
rect	128	269	129	270
rect	129	269	130	270
rect	130	269	131	270
rect	131	269	132	270
rect	132	269	133	270
rect	133	269	134	270
rect	134	269	135	270
rect	135	269	136	270
rect	136	269	137	270
rect	137	269	138	270
rect	138	269	139	270
rect	139	269	140	270
rect	140	269	141	270
rect	141	269	142	270
rect	142	269	143	270
rect	143	269	144	270
rect	144	269	145	270
rect	145	269	146	270
rect	146	269	147	270
rect	147	269	148	270
rect	148	269	149	270
rect	149	269	150	270
rect	150	269	151	270
rect	151	269	152	270
rect	152	269	153	270
rect	153	269	154	270
rect	154	269	155	270
rect	155	269	156	270
rect	156	269	157	270
rect	157	269	158	270
rect	158	269	159	270
rect	159	269	160	270
rect	160	269	161	270
rect	161	269	162	270
rect	162	269	163	270
rect	163	269	164	270
rect	164	269	165	270
rect	165	269	166	270
rect	166	269	167	270
rect	167	269	168	270
rect	168	269	169	270
rect	169	269	170	270
rect	170	269	171	270
rect	171	269	172	270
rect	172	269	173	270
rect	173	269	174	270
rect	174	269	175	270
rect	175	269	176	270
rect	176	269	177	270
rect	177	269	178	270
rect	178	269	179	270
rect	179	269	180	270
rect	180	269	181	270
rect	181	269	182	270
rect	182	269	183	270
rect	184	269	185	270
rect	185	269	186	270
rect	186	269	187	270
rect	187	269	188	270
rect	188	269	189	270
rect	189	269	190	270
rect	190	269	191	270
rect	191	269	192	270
rect	192	269	193	270
rect	193	269	194	270
rect	194	269	195	270
rect	195	269	196	270
rect	196	269	197	270
rect	197	269	198	270
rect	198	269	199	270
rect	199	269	200	270
rect	200	269	201	270
rect	201	269	202	270
rect	203	269	204	270
rect	204	269	205	270
rect	205	269	206	270
rect	206	269	207	270
rect	207	269	208	270
rect	208	269	209	270
rect	210	269	211	270
rect	211	269	212	270
rect	212	269	213	270
rect	213	269	214	270
rect	214	269	215	270
rect	215	269	216	270
rect	217	269	218	270
rect	218	269	219	270
rect	219	269	220	270
rect	220	269	221	270
rect	221	269	222	270
rect	222	269	223	270
rect	223	269	224	270
rect	224	269	225	270
rect	225	269	226	270
rect	226	269	227	270
rect	227	269	228	270
rect	228	269	229	270
rect	229	269	230	270
rect	230	269	231	270
rect	231	269	232	270
rect	232	269	233	270
rect	233	269	234	270
rect	234	269	235	270
rect	235	269	236	270
rect	236	269	237	270
rect	237	269	238	270
rect	238	269	239	270
rect	239	269	240	270
rect	240	269	241	270
rect	241	269	242	270
rect	242	269	243	270
rect	243	269	244	270
rect	245	269	246	270
rect	246	269	247	270
rect	247	269	248	270
rect	248	269	249	270
rect	249	269	250	270
rect	250	269	251	270
rect	252	269	253	270
rect	253	269	254	270
rect	254	269	255	270
rect	255	269	256	270
rect	256	269	257	270
rect	257	269	258	270
rect	258	269	259	270
rect	259	269	260	270
rect	260	269	261	270
rect	261	269	262	270
rect	262	269	263	270
rect	263	269	264	270
rect	264	269	265	270
rect	265	269	266	270
rect	266	269	267	270
rect	267	269	268	270
rect	268	269	269	270
rect	269	269	270	270
rect	270	269	271	270
rect	271	269	272	270
rect	272	269	273	270
rect	273	269	274	270
rect	274	269	275	270
rect	275	269	276	270
rect	276	269	277	270
rect	277	269	278	270
rect	278	269	279	270
rect	279	269	280	270
rect	280	269	281	270
rect	281	269	282	270
rect	282	269	283	270
rect	283	269	284	270
rect	284	269	285	270
rect	285	269	286	270
rect	286	269	287	270
rect	287	269	288	270
rect	288	269	289	270
rect	289	269	290	270
rect	290	269	291	270
rect	291	269	292	270
rect	292	269	293	270
rect	293	269	294	270
rect	294	269	295	270
rect	295	269	296	270
rect	296	269	297	270
rect	297	269	298	270
rect	298	269	299	270
rect	299	269	300	270
rect	301	269	302	270
rect	302	269	303	270
rect	303	269	304	270
rect	304	269	305	270
rect	305	269	306	270
rect	306	269	307	270
rect	307	269	308	270
rect	308	269	309	270
rect	309	269	310	270
rect	310	269	311	270
rect	311	269	312	270
rect	312	269	313	270
rect	313	269	314	270
rect	314	269	315	270
rect	315	269	316	270
rect	316	269	317	270
rect	317	269	318	270
rect	318	269	319	270
rect	319	269	320	270
rect	320	269	321	270
rect	321	269	322	270
rect	322	269	323	270
rect	323	269	324	270
rect	324	269	325	270
rect	325	269	326	270
rect	326	269	327	270
rect	327	269	328	270
rect	328	269	329	270
rect	329	269	330	270
rect	330	269	331	270
rect	331	269	332	270
rect	332	269	333	270
rect	333	269	334	270
rect	334	269	335	270
rect	335	269	336	270
rect	336	269	337	270
rect	337	269	338	270
rect	338	269	339	270
rect	339	269	340	270
rect	340	269	341	270
rect	341	269	342	270
rect	342	269	343	270
rect	343	269	344	270
rect	344	269	345	270
rect	345	269	346	270
rect	346	269	347	270
rect	347	269	348	270
rect	348	269	349	270
rect	349	269	350	270
rect	350	269	351	270
rect	351	269	352	270
rect	353	269	354	270
rect	354	269	355	270
rect	355	269	356	270
rect	356	269	357	270
rect	357	269	358	270
rect	358	269	359	270
rect	359	269	360	270
rect	360	269	361	270
rect	361	269	362	270
rect	362	269	363	270
rect	363	269	364	270
rect	364	269	365	270
rect	365	269	366	270
rect	366	269	367	270
rect	367	269	368	270
rect	368	269	369	270
rect	369	269	370	270
rect	370	269	371	270
rect	371	269	372	270
rect	372	269	373	270
rect	373	269	374	270
rect	374	269	375	270
rect	375	269	376	270
rect	376	269	377	270
rect	377	269	378	270
rect	378	269	379	270
rect	379	269	380	270
rect	380	269	381	270
rect	381	269	382	270
rect	382	269	383	270
rect	383	269	384	270
rect	384	269	385	270
rect	385	269	386	270
rect	386	269	387	270
rect	387	269	388	270
rect	388	269	389	270
rect	0	270	1	271
rect	1	270	2	271
rect	2	270	3	271
rect	3	270	4	271
rect	4	270	5	271
rect	5	270	6	271
rect	7	270	8	271
rect	8	270	9	271
rect	9	270	10	271
rect	10	270	11	271
rect	11	270	12	271
rect	12	270	13	271
rect	14	270	15	271
rect	15	270	16	271
rect	16	270	17	271
rect	17	270	18	271
rect	18	270	19	271
rect	19	270	20	271
rect	20	270	21	271
rect	21	270	22	271
rect	22	270	23	271
rect	23	270	24	271
rect	24	270	25	271
rect	25	270	26	271
rect	26	270	27	271
rect	27	270	28	271
rect	28	270	29	271
rect	29	270	30	271
rect	30	270	31	271
rect	31	270	32	271
rect	32	270	33	271
rect	33	270	34	271
rect	34	270	35	271
rect	35	270	36	271
rect	36	270	37	271
rect	37	270	38	271
rect	38	270	39	271
rect	39	270	40	271
rect	40	270	41	271
rect	41	270	42	271
rect	42	270	43	271
rect	43	270	44	271
rect	44	270	45	271
rect	45	270	46	271
rect	46	270	47	271
rect	47	270	48	271
rect	48	270	49	271
rect	49	270	50	271
rect	50	270	51	271
rect	51	270	52	271
rect	52	270	53	271
rect	53	270	54	271
rect	54	270	55	271
rect	55	270	56	271
rect	56	270	57	271
rect	57	270	58	271
rect	58	270	59	271
rect	59	270	60	271
rect	60	270	61	271
rect	61	270	62	271
rect	62	270	63	271
rect	63	270	64	271
rect	64	270	65	271
rect	65	270	66	271
rect	66	270	67	271
rect	67	270	68	271
rect	68	270	69	271
rect	69	270	70	271
rect	70	270	71	271
rect	71	270	72	271
rect	72	270	73	271
rect	73	270	74	271
rect	74	270	75	271
rect	75	270	76	271
rect	76	270	77	271
rect	77	270	78	271
rect	78	270	79	271
rect	79	270	80	271
rect	80	270	81	271
rect	81	270	82	271
rect	82	270	83	271
rect	84	270	85	271
rect	85	270	86	271
rect	86	270	87	271
rect	87	270	88	271
rect	88	270	89	271
rect	89	270	90	271
rect	90	270	91	271
rect	91	270	92	271
rect	92	270	93	271
rect	93	270	94	271
rect	94	270	95	271
rect	95	270	96	271
rect	96	270	97	271
rect	97	270	98	271
rect	98	270	99	271
rect	99	270	100	271
rect	100	270	101	271
rect	101	270	102	271
rect	102	270	103	271
rect	103	270	104	271
rect	104	270	105	271
rect	105	270	106	271
rect	106	270	107	271
rect	107	270	108	271
rect	108	270	109	271
rect	109	270	110	271
rect	110	270	111	271
rect	111	270	112	271
rect	112	270	113	271
rect	113	270	114	271
rect	114	270	115	271
rect	115	270	116	271
rect	116	270	117	271
rect	117	270	118	271
rect	118	270	119	271
rect	119	270	120	271
rect	120	270	121	271
rect	121	270	122	271
rect	122	270	123	271
rect	123	270	124	271
rect	124	270	125	271
rect	125	270	126	271
rect	126	270	127	271
rect	127	270	128	271
rect	128	270	129	271
rect	129	270	130	271
rect	130	270	131	271
rect	131	270	132	271
rect	132	270	133	271
rect	133	270	134	271
rect	134	270	135	271
rect	135	270	136	271
rect	136	270	137	271
rect	137	270	138	271
rect	138	270	139	271
rect	139	270	140	271
rect	140	270	141	271
rect	141	270	142	271
rect	142	270	143	271
rect	143	270	144	271
rect	144	270	145	271
rect	145	270	146	271
rect	146	270	147	271
rect	147	270	148	271
rect	148	270	149	271
rect	149	270	150	271
rect	150	270	151	271
rect	151	270	152	271
rect	152	270	153	271
rect	153	270	154	271
rect	154	270	155	271
rect	155	270	156	271
rect	156	270	157	271
rect	157	270	158	271
rect	158	270	159	271
rect	159	270	160	271
rect	160	270	161	271
rect	161	270	162	271
rect	162	270	163	271
rect	163	270	164	271
rect	164	270	165	271
rect	165	270	166	271
rect	166	270	167	271
rect	167	270	168	271
rect	168	270	169	271
rect	169	270	170	271
rect	170	270	171	271
rect	171	270	172	271
rect	172	270	173	271
rect	173	270	174	271
rect	174	270	175	271
rect	175	270	176	271
rect	176	270	177	271
rect	177	270	178	271
rect	178	270	179	271
rect	179	270	180	271
rect	180	270	181	271
rect	181	270	182	271
rect	182	270	183	271
rect	184	270	185	271
rect	185	270	186	271
rect	186	270	187	271
rect	187	270	188	271
rect	188	270	189	271
rect	189	270	190	271
rect	190	270	191	271
rect	191	270	192	271
rect	192	270	193	271
rect	193	270	194	271
rect	194	270	195	271
rect	195	270	196	271
rect	196	270	197	271
rect	197	270	198	271
rect	198	270	199	271
rect	199	270	200	271
rect	200	270	201	271
rect	201	270	202	271
rect	203	270	204	271
rect	204	270	205	271
rect	205	270	206	271
rect	206	270	207	271
rect	207	270	208	271
rect	208	270	209	271
rect	210	270	211	271
rect	211	270	212	271
rect	212	270	213	271
rect	213	270	214	271
rect	214	270	215	271
rect	215	270	216	271
rect	217	270	218	271
rect	218	270	219	271
rect	219	270	220	271
rect	220	270	221	271
rect	221	270	222	271
rect	222	270	223	271
rect	223	270	224	271
rect	224	270	225	271
rect	225	270	226	271
rect	226	270	227	271
rect	227	270	228	271
rect	228	270	229	271
rect	229	270	230	271
rect	230	270	231	271
rect	231	270	232	271
rect	232	270	233	271
rect	233	270	234	271
rect	234	270	235	271
rect	235	270	236	271
rect	236	270	237	271
rect	237	270	238	271
rect	238	270	239	271
rect	239	270	240	271
rect	240	270	241	271
rect	241	270	242	271
rect	242	270	243	271
rect	243	270	244	271
rect	245	270	246	271
rect	246	270	247	271
rect	247	270	248	271
rect	248	270	249	271
rect	249	270	250	271
rect	250	270	251	271
rect	252	270	253	271
rect	253	270	254	271
rect	254	270	255	271
rect	255	270	256	271
rect	256	270	257	271
rect	257	270	258	271
rect	258	270	259	271
rect	259	270	260	271
rect	260	270	261	271
rect	261	270	262	271
rect	262	270	263	271
rect	263	270	264	271
rect	264	270	265	271
rect	265	270	266	271
rect	266	270	267	271
rect	267	270	268	271
rect	268	270	269	271
rect	269	270	270	271
rect	270	270	271	271
rect	271	270	272	271
rect	272	270	273	271
rect	273	270	274	271
rect	274	270	275	271
rect	275	270	276	271
rect	276	270	277	271
rect	277	270	278	271
rect	278	270	279	271
rect	279	270	280	271
rect	280	270	281	271
rect	281	270	282	271
rect	282	270	283	271
rect	283	270	284	271
rect	284	270	285	271
rect	285	270	286	271
rect	286	270	287	271
rect	287	270	288	271
rect	288	270	289	271
rect	289	270	290	271
rect	290	270	291	271
rect	291	270	292	271
rect	292	270	293	271
rect	293	270	294	271
rect	294	270	295	271
rect	295	270	296	271
rect	296	270	297	271
rect	297	270	298	271
rect	298	270	299	271
rect	299	270	300	271
rect	301	270	302	271
rect	302	270	303	271
rect	303	270	304	271
rect	304	270	305	271
rect	305	270	306	271
rect	306	270	307	271
rect	307	270	308	271
rect	308	270	309	271
rect	309	270	310	271
rect	310	270	311	271
rect	311	270	312	271
rect	312	270	313	271
rect	313	270	314	271
rect	314	270	315	271
rect	315	270	316	271
rect	316	270	317	271
rect	317	270	318	271
rect	318	270	319	271
rect	319	270	320	271
rect	320	270	321	271
rect	321	270	322	271
rect	322	270	323	271
rect	323	270	324	271
rect	324	270	325	271
rect	325	270	326	271
rect	326	270	327	271
rect	327	270	328	271
rect	328	270	329	271
rect	329	270	330	271
rect	330	270	331	271
rect	331	270	332	271
rect	332	270	333	271
rect	333	270	334	271
rect	334	270	335	271
rect	335	270	336	271
rect	336	270	337	271
rect	337	270	338	271
rect	338	270	339	271
rect	339	270	340	271
rect	340	270	341	271
rect	341	270	342	271
rect	342	270	343	271
rect	343	270	344	271
rect	344	270	345	271
rect	345	270	346	271
rect	346	270	347	271
rect	347	270	348	271
rect	348	270	349	271
rect	349	270	350	271
rect	350	270	351	271
rect	351	270	352	271
rect	353	270	354	271
rect	354	270	355	271
rect	355	270	356	271
rect	356	270	357	271
rect	357	270	358	271
rect	358	270	359	271
rect	359	270	360	271
rect	360	270	361	271
rect	361	270	362	271
rect	362	270	363	271
rect	363	270	364	271
rect	364	270	365	271
rect	365	270	366	271
rect	366	270	367	271
rect	367	270	368	271
rect	368	270	369	271
rect	369	270	370	271
rect	370	270	371	271
rect	371	270	372	271
rect	372	270	373	271
rect	373	270	374	271
rect	374	270	375	271
rect	375	270	376	271
rect	376	270	377	271
rect	377	270	378	271
rect	378	270	379	271
rect	379	270	380	271
rect	380	270	381	271
rect	381	270	382	271
rect	382	270	383	271
rect	383	270	384	271
rect	384	270	385	271
rect	385	270	386	271
rect	386	270	387	271
rect	387	270	388	271
rect	388	270	389	271
rect	0	271	1	272
rect	1	271	2	272
rect	2	271	3	272
rect	3	271	4	272
rect	4	271	5	272
rect	5	271	6	272
rect	7	271	8	272
rect	8	271	9	272
rect	9	271	10	272
rect	10	271	11	272
rect	11	271	12	272
rect	12	271	13	272
rect	14	271	15	272
rect	15	271	16	272
rect	16	271	17	272
rect	17	271	18	272
rect	18	271	19	272
rect	19	271	20	272
rect	20	271	21	272
rect	21	271	22	272
rect	22	271	23	272
rect	23	271	24	272
rect	24	271	25	272
rect	25	271	26	272
rect	26	271	27	272
rect	27	271	28	272
rect	28	271	29	272
rect	29	271	30	272
rect	30	271	31	272
rect	31	271	32	272
rect	32	271	33	272
rect	33	271	34	272
rect	34	271	35	272
rect	35	271	36	272
rect	36	271	37	272
rect	37	271	38	272
rect	38	271	39	272
rect	39	271	40	272
rect	40	271	41	272
rect	41	271	42	272
rect	42	271	43	272
rect	43	271	44	272
rect	44	271	45	272
rect	45	271	46	272
rect	46	271	47	272
rect	47	271	48	272
rect	48	271	49	272
rect	49	271	50	272
rect	50	271	51	272
rect	51	271	52	272
rect	52	271	53	272
rect	53	271	54	272
rect	54	271	55	272
rect	55	271	56	272
rect	56	271	57	272
rect	57	271	58	272
rect	58	271	59	272
rect	59	271	60	272
rect	60	271	61	272
rect	61	271	62	272
rect	62	271	63	272
rect	63	271	64	272
rect	64	271	65	272
rect	65	271	66	272
rect	66	271	67	272
rect	67	271	68	272
rect	68	271	69	272
rect	69	271	70	272
rect	70	271	71	272
rect	71	271	72	272
rect	72	271	73	272
rect	73	271	74	272
rect	74	271	75	272
rect	75	271	76	272
rect	76	271	77	272
rect	77	271	78	272
rect	78	271	79	272
rect	79	271	80	272
rect	80	271	81	272
rect	81	271	82	272
rect	82	271	83	272
rect	84	271	85	272
rect	85	271	86	272
rect	86	271	87	272
rect	87	271	88	272
rect	88	271	89	272
rect	89	271	90	272
rect	90	271	91	272
rect	91	271	92	272
rect	92	271	93	272
rect	93	271	94	272
rect	94	271	95	272
rect	95	271	96	272
rect	96	271	97	272
rect	97	271	98	272
rect	98	271	99	272
rect	99	271	100	272
rect	100	271	101	272
rect	101	271	102	272
rect	102	271	103	272
rect	103	271	104	272
rect	104	271	105	272
rect	105	271	106	272
rect	106	271	107	272
rect	107	271	108	272
rect	108	271	109	272
rect	109	271	110	272
rect	110	271	111	272
rect	111	271	112	272
rect	112	271	113	272
rect	113	271	114	272
rect	114	271	115	272
rect	115	271	116	272
rect	116	271	117	272
rect	117	271	118	272
rect	118	271	119	272
rect	119	271	120	272
rect	120	271	121	272
rect	121	271	122	272
rect	122	271	123	272
rect	123	271	124	272
rect	124	271	125	272
rect	125	271	126	272
rect	126	271	127	272
rect	127	271	128	272
rect	128	271	129	272
rect	129	271	130	272
rect	130	271	131	272
rect	131	271	132	272
rect	132	271	133	272
rect	133	271	134	272
rect	134	271	135	272
rect	135	271	136	272
rect	136	271	137	272
rect	137	271	138	272
rect	138	271	139	272
rect	139	271	140	272
rect	140	271	141	272
rect	141	271	142	272
rect	142	271	143	272
rect	143	271	144	272
rect	144	271	145	272
rect	145	271	146	272
rect	146	271	147	272
rect	147	271	148	272
rect	148	271	149	272
rect	149	271	150	272
rect	150	271	151	272
rect	151	271	152	272
rect	152	271	153	272
rect	153	271	154	272
rect	154	271	155	272
rect	155	271	156	272
rect	156	271	157	272
rect	157	271	158	272
rect	158	271	159	272
rect	159	271	160	272
rect	160	271	161	272
rect	161	271	162	272
rect	162	271	163	272
rect	163	271	164	272
rect	164	271	165	272
rect	165	271	166	272
rect	166	271	167	272
rect	167	271	168	272
rect	168	271	169	272
rect	169	271	170	272
rect	170	271	171	272
rect	171	271	172	272
rect	172	271	173	272
rect	173	271	174	272
rect	174	271	175	272
rect	175	271	176	272
rect	176	271	177	272
rect	177	271	178	272
rect	178	271	179	272
rect	179	271	180	272
rect	180	271	181	272
rect	181	271	182	272
rect	182	271	183	272
rect	184	271	185	272
rect	185	271	186	272
rect	186	271	187	272
rect	187	271	188	272
rect	188	271	189	272
rect	189	271	190	272
rect	190	271	191	272
rect	191	271	192	272
rect	192	271	193	272
rect	193	271	194	272
rect	194	271	195	272
rect	195	271	196	272
rect	196	271	197	272
rect	197	271	198	272
rect	198	271	199	272
rect	199	271	200	272
rect	200	271	201	272
rect	201	271	202	272
rect	203	271	204	272
rect	204	271	205	272
rect	205	271	206	272
rect	206	271	207	272
rect	207	271	208	272
rect	208	271	209	272
rect	210	271	211	272
rect	211	271	212	272
rect	212	271	213	272
rect	213	271	214	272
rect	214	271	215	272
rect	215	271	216	272
rect	217	271	218	272
rect	218	271	219	272
rect	219	271	220	272
rect	220	271	221	272
rect	221	271	222	272
rect	222	271	223	272
rect	223	271	224	272
rect	224	271	225	272
rect	225	271	226	272
rect	226	271	227	272
rect	227	271	228	272
rect	228	271	229	272
rect	229	271	230	272
rect	230	271	231	272
rect	231	271	232	272
rect	232	271	233	272
rect	233	271	234	272
rect	234	271	235	272
rect	235	271	236	272
rect	236	271	237	272
rect	237	271	238	272
rect	238	271	239	272
rect	239	271	240	272
rect	240	271	241	272
rect	241	271	242	272
rect	242	271	243	272
rect	243	271	244	272
rect	245	271	246	272
rect	246	271	247	272
rect	247	271	248	272
rect	248	271	249	272
rect	249	271	250	272
rect	250	271	251	272
rect	252	271	253	272
rect	253	271	254	272
rect	254	271	255	272
rect	255	271	256	272
rect	256	271	257	272
rect	257	271	258	272
rect	258	271	259	272
rect	259	271	260	272
rect	260	271	261	272
rect	261	271	262	272
rect	262	271	263	272
rect	263	271	264	272
rect	264	271	265	272
rect	265	271	266	272
rect	266	271	267	272
rect	267	271	268	272
rect	268	271	269	272
rect	269	271	270	272
rect	270	271	271	272
rect	271	271	272	272
rect	272	271	273	272
rect	273	271	274	272
rect	274	271	275	272
rect	275	271	276	272
rect	276	271	277	272
rect	277	271	278	272
rect	278	271	279	272
rect	279	271	280	272
rect	280	271	281	272
rect	281	271	282	272
rect	282	271	283	272
rect	283	271	284	272
rect	284	271	285	272
rect	285	271	286	272
rect	286	271	287	272
rect	287	271	288	272
rect	288	271	289	272
rect	289	271	290	272
rect	290	271	291	272
rect	291	271	292	272
rect	292	271	293	272
rect	293	271	294	272
rect	294	271	295	272
rect	295	271	296	272
rect	296	271	297	272
rect	297	271	298	272
rect	298	271	299	272
rect	299	271	300	272
rect	301	271	302	272
rect	302	271	303	272
rect	303	271	304	272
rect	304	271	305	272
rect	305	271	306	272
rect	306	271	307	272
rect	307	271	308	272
rect	308	271	309	272
rect	309	271	310	272
rect	310	271	311	272
rect	311	271	312	272
rect	312	271	313	272
rect	313	271	314	272
rect	314	271	315	272
rect	315	271	316	272
rect	316	271	317	272
rect	317	271	318	272
rect	318	271	319	272
rect	319	271	320	272
rect	320	271	321	272
rect	321	271	322	272
rect	322	271	323	272
rect	323	271	324	272
rect	324	271	325	272
rect	325	271	326	272
rect	326	271	327	272
rect	327	271	328	272
rect	328	271	329	272
rect	329	271	330	272
rect	330	271	331	272
rect	331	271	332	272
rect	332	271	333	272
rect	333	271	334	272
rect	334	271	335	272
rect	335	271	336	272
rect	336	271	337	272
rect	337	271	338	272
rect	338	271	339	272
rect	339	271	340	272
rect	340	271	341	272
rect	341	271	342	272
rect	342	271	343	272
rect	343	271	344	272
rect	344	271	345	272
rect	345	271	346	272
rect	346	271	347	272
rect	347	271	348	272
rect	348	271	349	272
rect	349	271	350	272
rect	350	271	351	272
rect	351	271	352	272
rect	353	271	354	272
rect	354	271	355	272
rect	355	271	356	272
rect	356	271	357	272
rect	357	271	358	272
rect	358	271	359	272
rect	359	271	360	272
rect	360	271	361	272
rect	361	271	362	272
rect	362	271	363	272
rect	363	271	364	272
rect	364	271	365	272
rect	365	271	366	272
rect	366	271	367	272
rect	367	271	368	272
rect	368	271	369	272
rect	369	271	370	272
rect	370	271	371	272
rect	371	271	372	272
rect	372	271	373	272
rect	373	271	374	272
rect	374	271	375	272
rect	375	271	376	272
rect	376	271	377	272
rect	377	271	378	272
rect	378	271	379	272
rect	379	271	380	272
rect	380	271	381	272
rect	381	271	382	272
rect	382	271	383	272
rect	383	271	384	272
rect	384	271	385	272
rect	385	271	386	272
rect	386	271	387	272
rect	387	271	388	272
rect	388	271	389	272
rect	0	272	1	273
rect	1	272	2	273
rect	2	272	3	273
rect	3	272	4	273
rect	4	272	5	273
rect	5	272	6	273
rect	7	272	8	273
rect	8	272	9	273
rect	9	272	10	273
rect	10	272	11	273
rect	11	272	12	273
rect	12	272	13	273
rect	14	272	15	273
rect	15	272	16	273
rect	16	272	17	273
rect	17	272	18	273
rect	18	272	19	273
rect	19	272	20	273
rect	20	272	21	273
rect	21	272	22	273
rect	22	272	23	273
rect	23	272	24	273
rect	24	272	25	273
rect	25	272	26	273
rect	26	272	27	273
rect	27	272	28	273
rect	28	272	29	273
rect	29	272	30	273
rect	30	272	31	273
rect	31	272	32	273
rect	32	272	33	273
rect	33	272	34	273
rect	34	272	35	273
rect	35	272	36	273
rect	36	272	37	273
rect	37	272	38	273
rect	38	272	39	273
rect	39	272	40	273
rect	40	272	41	273
rect	41	272	42	273
rect	42	272	43	273
rect	43	272	44	273
rect	44	272	45	273
rect	45	272	46	273
rect	46	272	47	273
rect	47	272	48	273
rect	48	272	49	273
rect	49	272	50	273
rect	50	272	51	273
rect	51	272	52	273
rect	52	272	53	273
rect	53	272	54	273
rect	54	272	55	273
rect	55	272	56	273
rect	56	272	57	273
rect	57	272	58	273
rect	58	272	59	273
rect	59	272	60	273
rect	60	272	61	273
rect	61	272	62	273
rect	62	272	63	273
rect	63	272	64	273
rect	64	272	65	273
rect	65	272	66	273
rect	66	272	67	273
rect	67	272	68	273
rect	68	272	69	273
rect	69	272	70	273
rect	70	272	71	273
rect	71	272	72	273
rect	72	272	73	273
rect	73	272	74	273
rect	74	272	75	273
rect	75	272	76	273
rect	76	272	77	273
rect	77	272	78	273
rect	78	272	79	273
rect	79	272	80	273
rect	80	272	81	273
rect	81	272	82	273
rect	82	272	83	273
rect	84	272	85	273
rect	85	272	86	273
rect	86	272	87	273
rect	87	272	88	273
rect	88	272	89	273
rect	89	272	90	273
rect	90	272	91	273
rect	91	272	92	273
rect	92	272	93	273
rect	93	272	94	273
rect	94	272	95	273
rect	95	272	96	273
rect	96	272	97	273
rect	97	272	98	273
rect	98	272	99	273
rect	99	272	100	273
rect	100	272	101	273
rect	101	272	102	273
rect	102	272	103	273
rect	103	272	104	273
rect	104	272	105	273
rect	105	272	106	273
rect	106	272	107	273
rect	107	272	108	273
rect	108	272	109	273
rect	109	272	110	273
rect	110	272	111	273
rect	111	272	112	273
rect	112	272	113	273
rect	113	272	114	273
rect	114	272	115	273
rect	115	272	116	273
rect	116	272	117	273
rect	117	272	118	273
rect	118	272	119	273
rect	119	272	120	273
rect	120	272	121	273
rect	121	272	122	273
rect	122	272	123	273
rect	123	272	124	273
rect	124	272	125	273
rect	125	272	126	273
rect	126	272	127	273
rect	127	272	128	273
rect	128	272	129	273
rect	129	272	130	273
rect	130	272	131	273
rect	131	272	132	273
rect	132	272	133	273
rect	133	272	134	273
rect	134	272	135	273
rect	135	272	136	273
rect	136	272	137	273
rect	137	272	138	273
rect	138	272	139	273
rect	139	272	140	273
rect	140	272	141	273
rect	141	272	142	273
rect	142	272	143	273
rect	143	272	144	273
rect	144	272	145	273
rect	145	272	146	273
rect	146	272	147	273
rect	147	272	148	273
rect	148	272	149	273
rect	149	272	150	273
rect	150	272	151	273
rect	151	272	152	273
rect	152	272	153	273
rect	153	272	154	273
rect	154	272	155	273
rect	155	272	156	273
rect	156	272	157	273
rect	157	272	158	273
rect	158	272	159	273
rect	159	272	160	273
rect	160	272	161	273
rect	161	272	162	273
rect	162	272	163	273
rect	163	272	164	273
rect	164	272	165	273
rect	165	272	166	273
rect	166	272	167	273
rect	167	272	168	273
rect	168	272	169	273
rect	169	272	170	273
rect	170	272	171	273
rect	171	272	172	273
rect	172	272	173	273
rect	173	272	174	273
rect	174	272	175	273
rect	175	272	176	273
rect	176	272	177	273
rect	177	272	178	273
rect	178	272	179	273
rect	179	272	180	273
rect	180	272	181	273
rect	181	272	182	273
rect	182	272	183	273
rect	184	272	185	273
rect	185	272	186	273
rect	186	272	187	273
rect	187	272	188	273
rect	188	272	189	273
rect	189	272	190	273
rect	190	272	191	273
rect	191	272	192	273
rect	192	272	193	273
rect	193	272	194	273
rect	194	272	195	273
rect	195	272	196	273
rect	196	272	197	273
rect	197	272	198	273
rect	198	272	199	273
rect	199	272	200	273
rect	200	272	201	273
rect	201	272	202	273
rect	203	272	204	273
rect	204	272	205	273
rect	205	272	206	273
rect	206	272	207	273
rect	207	272	208	273
rect	208	272	209	273
rect	210	272	211	273
rect	211	272	212	273
rect	212	272	213	273
rect	213	272	214	273
rect	214	272	215	273
rect	215	272	216	273
rect	217	272	218	273
rect	218	272	219	273
rect	219	272	220	273
rect	220	272	221	273
rect	221	272	222	273
rect	222	272	223	273
rect	223	272	224	273
rect	224	272	225	273
rect	225	272	226	273
rect	226	272	227	273
rect	227	272	228	273
rect	228	272	229	273
rect	229	272	230	273
rect	230	272	231	273
rect	231	272	232	273
rect	232	272	233	273
rect	233	272	234	273
rect	234	272	235	273
rect	235	272	236	273
rect	236	272	237	273
rect	237	272	238	273
rect	238	272	239	273
rect	239	272	240	273
rect	240	272	241	273
rect	241	272	242	273
rect	242	272	243	273
rect	243	272	244	273
rect	245	272	246	273
rect	246	272	247	273
rect	247	272	248	273
rect	248	272	249	273
rect	249	272	250	273
rect	250	272	251	273
rect	252	272	253	273
rect	253	272	254	273
rect	254	272	255	273
rect	255	272	256	273
rect	256	272	257	273
rect	257	272	258	273
rect	258	272	259	273
rect	259	272	260	273
rect	260	272	261	273
rect	261	272	262	273
rect	262	272	263	273
rect	263	272	264	273
rect	264	272	265	273
rect	265	272	266	273
rect	266	272	267	273
rect	267	272	268	273
rect	268	272	269	273
rect	269	272	270	273
rect	270	272	271	273
rect	271	272	272	273
rect	272	272	273	273
rect	273	272	274	273
rect	274	272	275	273
rect	275	272	276	273
rect	276	272	277	273
rect	277	272	278	273
rect	278	272	279	273
rect	279	272	280	273
rect	280	272	281	273
rect	281	272	282	273
rect	282	272	283	273
rect	283	272	284	273
rect	284	272	285	273
rect	285	272	286	273
rect	286	272	287	273
rect	287	272	288	273
rect	288	272	289	273
rect	289	272	290	273
rect	290	272	291	273
rect	291	272	292	273
rect	292	272	293	273
rect	293	272	294	273
rect	294	272	295	273
rect	295	272	296	273
rect	296	272	297	273
rect	297	272	298	273
rect	298	272	299	273
rect	299	272	300	273
rect	301	272	302	273
rect	302	272	303	273
rect	303	272	304	273
rect	304	272	305	273
rect	305	272	306	273
rect	306	272	307	273
rect	307	272	308	273
rect	308	272	309	273
rect	309	272	310	273
rect	310	272	311	273
rect	311	272	312	273
rect	312	272	313	273
rect	313	272	314	273
rect	314	272	315	273
rect	315	272	316	273
rect	316	272	317	273
rect	317	272	318	273
rect	318	272	319	273
rect	319	272	320	273
rect	320	272	321	273
rect	321	272	322	273
rect	322	272	323	273
rect	323	272	324	273
rect	324	272	325	273
rect	325	272	326	273
rect	326	272	327	273
rect	327	272	328	273
rect	328	272	329	273
rect	329	272	330	273
rect	330	272	331	273
rect	331	272	332	273
rect	332	272	333	273
rect	333	272	334	273
rect	334	272	335	273
rect	335	272	336	273
rect	336	272	337	273
rect	337	272	338	273
rect	338	272	339	273
rect	339	272	340	273
rect	340	272	341	273
rect	341	272	342	273
rect	342	272	343	273
rect	343	272	344	273
rect	344	272	345	273
rect	345	272	346	273
rect	346	272	347	273
rect	347	272	348	273
rect	348	272	349	273
rect	349	272	350	273
rect	350	272	351	273
rect	351	272	352	273
rect	353	272	354	273
rect	354	272	355	273
rect	355	272	356	273
rect	356	272	357	273
rect	357	272	358	273
rect	358	272	359	273
rect	359	272	360	273
rect	360	272	361	273
rect	361	272	362	273
rect	362	272	363	273
rect	363	272	364	273
rect	364	272	365	273
rect	365	272	366	273
rect	366	272	367	273
rect	367	272	368	273
rect	368	272	369	273
rect	369	272	370	273
rect	370	272	371	273
rect	371	272	372	273
rect	372	272	373	273
rect	373	272	374	273
rect	374	272	375	273
rect	375	272	376	273
rect	376	272	377	273
rect	377	272	378	273
rect	378	272	379	273
rect	379	272	380	273
rect	380	272	381	273
rect	381	272	382	273
rect	382	272	383	273
rect	383	272	384	273
rect	384	272	385	273
rect	385	272	386	273
rect	386	272	387	273
rect	387	272	388	273
rect	388	272	389	273
rect	0	273	1	274
rect	1	273	2	274
rect	2	273	3	274
rect	3	273	4	274
rect	4	273	5	274
rect	5	273	6	274
rect	7	273	8	274
rect	8	273	9	274
rect	9	273	10	274
rect	10	273	11	274
rect	11	273	12	274
rect	12	273	13	274
rect	14	273	15	274
rect	15	273	16	274
rect	16	273	17	274
rect	17	273	18	274
rect	18	273	19	274
rect	19	273	20	274
rect	20	273	21	274
rect	21	273	22	274
rect	22	273	23	274
rect	23	273	24	274
rect	24	273	25	274
rect	25	273	26	274
rect	26	273	27	274
rect	27	273	28	274
rect	28	273	29	274
rect	29	273	30	274
rect	30	273	31	274
rect	31	273	32	274
rect	32	273	33	274
rect	33	273	34	274
rect	34	273	35	274
rect	35	273	36	274
rect	36	273	37	274
rect	37	273	38	274
rect	38	273	39	274
rect	39	273	40	274
rect	40	273	41	274
rect	41	273	42	274
rect	42	273	43	274
rect	43	273	44	274
rect	44	273	45	274
rect	45	273	46	274
rect	46	273	47	274
rect	47	273	48	274
rect	48	273	49	274
rect	49	273	50	274
rect	50	273	51	274
rect	51	273	52	274
rect	52	273	53	274
rect	53	273	54	274
rect	54	273	55	274
rect	55	273	56	274
rect	56	273	57	274
rect	57	273	58	274
rect	58	273	59	274
rect	59	273	60	274
rect	60	273	61	274
rect	61	273	62	274
rect	62	273	63	274
rect	63	273	64	274
rect	64	273	65	274
rect	65	273	66	274
rect	66	273	67	274
rect	67	273	68	274
rect	68	273	69	274
rect	69	273	70	274
rect	70	273	71	274
rect	71	273	72	274
rect	72	273	73	274
rect	73	273	74	274
rect	74	273	75	274
rect	75	273	76	274
rect	76	273	77	274
rect	77	273	78	274
rect	78	273	79	274
rect	79	273	80	274
rect	80	273	81	274
rect	81	273	82	274
rect	82	273	83	274
rect	84	273	85	274
rect	85	273	86	274
rect	86	273	87	274
rect	87	273	88	274
rect	88	273	89	274
rect	89	273	90	274
rect	90	273	91	274
rect	91	273	92	274
rect	92	273	93	274
rect	93	273	94	274
rect	94	273	95	274
rect	95	273	96	274
rect	96	273	97	274
rect	97	273	98	274
rect	98	273	99	274
rect	99	273	100	274
rect	100	273	101	274
rect	101	273	102	274
rect	102	273	103	274
rect	103	273	104	274
rect	104	273	105	274
rect	105	273	106	274
rect	106	273	107	274
rect	107	273	108	274
rect	108	273	109	274
rect	109	273	110	274
rect	110	273	111	274
rect	111	273	112	274
rect	112	273	113	274
rect	113	273	114	274
rect	114	273	115	274
rect	115	273	116	274
rect	116	273	117	274
rect	117	273	118	274
rect	118	273	119	274
rect	119	273	120	274
rect	120	273	121	274
rect	121	273	122	274
rect	122	273	123	274
rect	123	273	124	274
rect	124	273	125	274
rect	125	273	126	274
rect	126	273	127	274
rect	127	273	128	274
rect	128	273	129	274
rect	129	273	130	274
rect	130	273	131	274
rect	131	273	132	274
rect	132	273	133	274
rect	133	273	134	274
rect	134	273	135	274
rect	135	273	136	274
rect	136	273	137	274
rect	137	273	138	274
rect	138	273	139	274
rect	139	273	140	274
rect	140	273	141	274
rect	141	273	142	274
rect	142	273	143	274
rect	143	273	144	274
rect	144	273	145	274
rect	145	273	146	274
rect	146	273	147	274
rect	147	273	148	274
rect	148	273	149	274
rect	149	273	150	274
rect	150	273	151	274
rect	151	273	152	274
rect	152	273	153	274
rect	153	273	154	274
rect	154	273	155	274
rect	155	273	156	274
rect	156	273	157	274
rect	157	273	158	274
rect	158	273	159	274
rect	159	273	160	274
rect	160	273	161	274
rect	161	273	162	274
rect	162	273	163	274
rect	163	273	164	274
rect	164	273	165	274
rect	165	273	166	274
rect	166	273	167	274
rect	167	273	168	274
rect	168	273	169	274
rect	169	273	170	274
rect	170	273	171	274
rect	171	273	172	274
rect	172	273	173	274
rect	173	273	174	274
rect	174	273	175	274
rect	175	273	176	274
rect	176	273	177	274
rect	177	273	178	274
rect	178	273	179	274
rect	179	273	180	274
rect	180	273	181	274
rect	181	273	182	274
rect	182	273	183	274
rect	184	273	185	274
rect	185	273	186	274
rect	186	273	187	274
rect	187	273	188	274
rect	188	273	189	274
rect	189	273	190	274
rect	190	273	191	274
rect	191	273	192	274
rect	192	273	193	274
rect	193	273	194	274
rect	194	273	195	274
rect	195	273	196	274
rect	196	273	197	274
rect	197	273	198	274
rect	198	273	199	274
rect	199	273	200	274
rect	200	273	201	274
rect	201	273	202	274
rect	203	273	204	274
rect	204	273	205	274
rect	205	273	206	274
rect	206	273	207	274
rect	207	273	208	274
rect	208	273	209	274
rect	210	273	211	274
rect	211	273	212	274
rect	212	273	213	274
rect	213	273	214	274
rect	214	273	215	274
rect	215	273	216	274
rect	217	273	218	274
rect	218	273	219	274
rect	219	273	220	274
rect	220	273	221	274
rect	221	273	222	274
rect	222	273	223	274
rect	223	273	224	274
rect	224	273	225	274
rect	225	273	226	274
rect	226	273	227	274
rect	227	273	228	274
rect	228	273	229	274
rect	229	273	230	274
rect	230	273	231	274
rect	231	273	232	274
rect	232	273	233	274
rect	233	273	234	274
rect	234	273	235	274
rect	235	273	236	274
rect	236	273	237	274
rect	237	273	238	274
rect	238	273	239	274
rect	239	273	240	274
rect	240	273	241	274
rect	241	273	242	274
rect	242	273	243	274
rect	243	273	244	274
rect	245	273	246	274
rect	246	273	247	274
rect	247	273	248	274
rect	248	273	249	274
rect	249	273	250	274
rect	250	273	251	274
rect	252	273	253	274
rect	253	273	254	274
rect	254	273	255	274
rect	255	273	256	274
rect	256	273	257	274
rect	257	273	258	274
rect	258	273	259	274
rect	259	273	260	274
rect	260	273	261	274
rect	261	273	262	274
rect	262	273	263	274
rect	263	273	264	274
rect	264	273	265	274
rect	265	273	266	274
rect	266	273	267	274
rect	267	273	268	274
rect	268	273	269	274
rect	269	273	270	274
rect	270	273	271	274
rect	271	273	272	274
rect	272	273	273	274
rect	273	273	274	274
rect	274	273	275	274
rect	275	273	276	274
rect	276	273	277	274
rect	277	273	278	274
rect	278	273	279	274
rect	279	273	280	274
rect	280	273	281	274
rect	281	273	282	274
rect	282	273	283	274
rect	283	273	284	274
rect	284	273	285	274
rect	285	273	286	274
rect	286	273	287	274
rect	287	273	288	274
rect	288	273	289	274
rect	289	273	290	274
rect	290	273	291	274
rect	291	273	292	274
rect	292	273	293	274
rect	293	273	294	274
rect	294	273	295	274
rect	295	273	296	274
rect	296	273	297	274
rect	297	273	298	274
rect	298	273	299	274
rect	299	273	300	274
rect	301	273	302	274
rect	302	273	303	274
rect	303	273	304	274
rect	304	273	305	274
rect	305	273	306	274
rect	306	273	307	274
rect	307	273	308	274
rect	308	273	309	274
rect	309	273	310	274
rect	310	273	311	274
rect	311	273	312	274
rect	312	273	313	274
rect	313	273	314	274
rect	314	273	315	274
rect	315	273	316	274
rect	316	273	317	274
rect	317	273	318	274
rect	318	273	319	274
rect	319	273	320	274
rect	320	273	321	274
rect	321	273	322	274
rect	322	273	323	274
rect	323	273	324	274
rect	324	273	325	274
rect	325	273	326	274
rect	326	273	327	274
rect	327	273	328	274
rect	328	273	329	274
rect	329	273	330	274
rect	330	273	331	274
rect	331	273	332	274
rect	332	273	333	274
rect	333	273	334	274
rect	334	273	335	274
rect	335	273	336	274
rect	336	273	337	274
rect	337	273	338	274
rect	338	273	339	274
rect	339	273	340	274
rect	340	273	341	274
rect	341	273	342	274
rect	342	273	343	274
rect	343	273	344	274
rect	344	273	345	274
rect	345	273	346	274
rect	346	273	347	274
rect	347	273	348	274
rect	348	273	349	274
rect	349	273	350	274
rect	350	273	351	274
rect	351	273	352	274
rect	353	273	354	274
rect	354	273	355	274
rect	355	273	356	274
rect	356	273	357	274
rect	357	273	358	274
rect	358	273	359	274
rect	359	273	360	274
rect	360	273	361	274
rect	361	273	362	274
rect	362	273	363	274
rect	363	273	364	274
rect	364	273	365	274
rect	365	273	366	274
rect	366	273	367	274
rect	367	273	368	274
rect	368	273	369	274
rect	369	273	370	274
rect	370	273	371	274
rect	371	273	372	274
rect	372	273	373	274
rect	373	273	374	274
rect	374	273	375	274
rect	375	273	376	274
rect	376	273	377	274
rect	377	273	378	274
rect	378	273	379	274
rect	379	273	380	274
rect	380	273	381	274
rect	381	273	382	274
rect	382	273	383	274
rect	383	273	384	274
rect	384	273	385	274
rect	385	273	386	274
rect	386	273	387	274
rect	387	273	388	274
rect	388	273	389	274
rect	0	274	1	275
rect	1	274	2	275
rect	2	274	3	275
rect	3	274	4	275
rect	4	274	5	275
rect	5	274	6	275
rect	7	274	8	275
rect	8	274	9	275
rect	9	274	10	275
rect	10	274	11	275
rect	11	274	12	275
rect	12	274	13	275
rect	14	274	15	275
rect	15	274	16	275
rect	16	274	17	275
rect	17	274	18	275
rect	18	274	19	275
rect	19	274	20	275
rect	20	274	21	275
rect	21	274	22	275
rect	22	274	23	275
rect	23	274	24	275
rect	24	274	25	275
rect	25	274	26	275
rect	26	274	27	275
rect	27	274	28	275
rect	28	274	29	275
rect	29	274	30	275
rect	30	274	31	275
rect	31	274	32	275
rect	32	274	33	275
rect	33	274	34	275
rect	34	274	35	275
rect	35	274	36	275
rect	36	274	37	275
rect	37	274	38	275
rect	38	274	39	275
rect	39	274	40	275
rect	40	274	41	275
rect	41	274	42	275
rect	42	274	43	275
rect	43	274	44	275
rect	44	274	45	275
rect	45	274	46	275
rect	46	274	47	275
rect	47	274	48	275
rect	48	274	49	275
rect	49	274	50	275
rect	50	274	51	275
rect	51	274	52	275
rect	52	274	53	275
rect	53	274	54	275
rect	54	274	55	275
rect	55	274	56	275
rect	56	274	57	275
rect	57	274	58	275
rect	58	274	59	275
rect	59	274	60	275
rect	60	274	61	275
rect	61	274	62	275
rect	62	274	63	275
rect	63	274	64	275
rect	64	274	65	275
rect	65	274	66	275
rect	66	274	67	275
rect	67	274	68	275
rect	68	274	69	275
rect	69	274	70	275
rect	70	274	71	275
rect	71	274	72	275
rect	72	274	73	275
rect	73	274	74	275
rect	74	274	75	275
rect	75	274	76	275
rect	76	274	77	275
rect	77	274	78	275
rect	78	274	79	275
rect	79	274	80	275
rect	80	274	81	275
rect	81	274	82	275
rect	82	274	83	275
rect	84	274	85	275
rect	85	274	86	275
rect	86	274	87	275
rect	87	274	88	275
rect	88	274	89	275
rect	89	274	90	275
rect	90	274	91	275
rect	91	274	92	275
rect	92	274	93	275
rect	93	274	94	275
rect	94	274	95	275
rect	95	274	96	275
rect	96	274	97	275
rect	97	274	98	275
rect	98	274	99	275
rect	99	274	100	275
rect	100	274	101	275
rect	101	274	102	275
rect	102	274	103	275
rect	103	274	104	275
rect	104	274	105	275
rect	105	274	106	275
rect	106	274	107	275
rect	107	274	108	275
rect	108	274	109	275
rect	109	274	110	275
rect	110	274	111	275
rect	111	274	112	275
rect	112	274	113	275
rect	113	274	114	275
rect	114	274	115	275
rect	115	274	116	275
rect	116	274	117	275
rect	117	274	118	275
rect	118	274	119	275
rect	119	274	120	275
rect	120	274	121	275
rect	121	274	122	275
rect	122	274	123	275
rect	123	274	124	275
rect	124	274	125	275
rect	125	274	126	275
rect	126	274	127	275
rect	127	274	128	275
rect	128	274	129	275
rect	129	274	130	275
rect	130	274	131	275
rect	131	274	132	275
rect	132	274	133	275
rect	133	274	134	275
rect	134	274	135	275
rect	135	274	136	275
rect	136	274	137	275
rect	137	274	138	275
rect	138	274	139	275
rect	139	274	140	275
rect	140	274	141	275
rect	141	274	142	275
rect	142	274	143	275
rect	143	274	144	275
rect	144	274	145	275
rect	145	274	146	275
rect	146	274	147	275
rect	147	274	148	275
rect	148	274	149	275
rect	149	274	150	275
rect	150	274	151	275
rect	151	274	152	275
rect	152	274	153	275
rect	153	274	154	275
rect	154	274	155	275
rect	155	274	156	275
rect	156	274	157	275
rect	157	274	158	275
rect	158	274	159	275
rect	159	274	160	275
rect	160	274	161	275
rect	161	274	162	275
rect	162	274	163	275
rect	163	274	164	275
rect	164	274	165	275
rect	165	274	166	275
rect	166	274	167	275
rect	167	274	168	275
rect	168	274	169	275
rect	169	274	170	275
rect	170	274	171	275
rect	171	274	172	275
rect	172	274	173	275
rect	173	274	174	275
rect	174	274	175	275
rect	175	274	176	275
rect	176	274	177	275
rect	177	274	178	275
rect	178	274	179	275
rect	179	274	180	275
rect	180	274	181	275
rect	181	274	182	275
rect	182	274	183	275
rect	184	274	185	275
rect	185	274	186	275
rect	186	274	187	275
rect	187	274	188	275
rect	188	274	189	275
rect	189	274	190	275
rect	190	274	191	275
rect	191	274	192	275
rect	192	274	193	275
rect	193	274	194	275
rect	194	274	195	275
rect	195	274	196	275
rect	196	274	197	275
rect	197	274	198	275
rect	198	274	199	275
rect	199	274	200	275
rect	200	274	201	275
rect	201	274	202	275
rect	203	274	204	275
rect	204	274	205	275
rect	205	274	206	275
rect	206	274	207	275
rect	207	274	208	275
rect	208	274	209	275
rect	210	274	211	275
rect	211	274	212	275
rect	212	274	213	275
rect	213	274	214	275
rect	214	274	215	275
rect	215	274	216	275
rect	217	274	218	275
rect	218	274	219	275
rect	219	274	220	275
rect	220	274	221	275
rect	221	274	222	275
rect	222	274	223	275
rect	223	274	224	275
rect	224	274	225	275
rect	225	274	226	275
rect	226	274	227	275
rect	227	274	228	275
rect	228	274	229	275
rect	229	274	230	275
rect	230	274	231	275
rect	231	274	232	275
rect	232	274	233	275
rect	233	274	234	275
rect	234	274	235	275
rect	235	274	236	275
rect	236	274	237	275
rect	237	274	238	275
rect	238	274	239	275
rect	239	274	240	275
rect	240	274	241	275
rect	241	274	242	275
rect	242	274	243	275
rect	243	274	244	275
rect	245	274	246	275
rect	246	274	247	275
rect	247	274	248	275
rect	248	274	249	275
rect	249	274	250	275
rect	250	274	251	275
rect	252	274	253	275
rect	253	274	254	275
rect	254	274	255	275
rect	255	274	256	275
rect	256	274	257	275
rect	257	274	258	275
rect	258	274	259	275
rect	259	274	260	275
rect	260	274	261	275
rect	261	274	262	275
rect	262	274	263	275
rect	263	274	264	275
rect	264	274	265	275
rect	265	274	266	275
rect	266	274	267	275
rect	267	274	268	275
rect	268	274	269	275
rect	269	274	270	275
rect	270	274	271	275
rect	271	274	272	275
rect	272	274	273	275
rect	273	274	274	275
rect	274	274	275	275
rect	275	274	276	275
rect	276	274	277	275
rect	277	274	278	275
rect	278	274	279	275
rect	279	274	280	275
rect	280	274	281	275
rect	281	274	282	275
rect	282	274	283	275
rect	283	274	284	275
rect	284	274	285	275
rect	285	274	286	275
rect	286	274	287	275
rect	287	274	288	275
rect	288	274	289	275
rect	289	274	290	275
rect	290	274	291	275
rect	291	274	292	275
rect	292	274	293	275
rect	293	274	294	275
rect	294	274	295	275
rect	295	274	296	275
rect	296	274	297	275
rect	297	274	298	275
rect	298	274	299	275
rect	299	274	300	275
rect	301	274	302	275
rect	302	274	303	275
rect	303	274	304	275
rect	304	274	305	275
rect	305	274	306	275
rect	306	274	307	275
rect	307	274	308	275
rect	308	274	309	275
rect	309	274	310	275
rect	310	274	311	275
rect	311	274	312	275
rect	312	274	313	275
rect	313	274	314	275
rect	314	274	315	275
rect	315	274	316	275
rect	316	274	317	275
rect	317	274	318	275
rect	318	274	319	275
rect	319	274	320	275
rect	320	274	321	275
rect	321	274	322	275
rect	322	274	323	275
rect	323	274	324	275
rect	324	274	325	275
rect	325	274	326	275
rect	326	274	327	275
rect	327	274	328	275
rect	328	274	329	275
rect	329	274	330	275
rect	330	274	331	275
rect	331	274	332	275
rect	332	274	333	275
rect	333	274	334	275
rect	334	274	335	275
rect	335	274	336	275
rect	336	274	337	275
rect	337	274	338	275
rect	338	274	339	275
rect	339	274	340	275
rect	340	274	341	275
rect	341	274	342	275
rect	342	274	343	275
rect	343	274	344	275
rect	344	274	345	275
rect	345	274	346	275
rect	346	274	347	275
rect	347	274	348	275
rect	348	274	349	275
rect	349	274	350	275
rect	350	274	351	275
rect	351	274	352	275
rect	353	274	354	275
rect	354	274	355	275
rect	355	274	356	275
rect	356	274	357	275
rect	357	274	358	275
rect	358	274	359	275
rect	359	274	360	275
rect	360	274	361	275
rect	361	274	362	275
rect	362	274	363	275
rect	363	274	364	275
rect	364	274	365	275
rect	365	274	366	275
rect	366	274	367	275
rect	367	274	368	275
rect	368	274	369	275
rect	369	274	370	275
rect	370	274	371	275
rect	371	274	372	275
rect	372	274	373	275
rect	373	274	374	275
rect	374	274	375	275
rect	375	274	376	275
rect	376	274	377	275
rect	377	274	378	275
rect	378	274	379	275
rect	379	274	380	275
rect	380	274	381	275
rect	381	274	382	275
rect	382	274	383	275
rect	383	274	384	275
rect	384	274	385	275
rect	385	274	386	275
rect	386	274	387	275
rect	387	274	388	275
rect	388	274	389	275
rect	0	290	1	291
rect	1	290	2	291
rect	2	290	3	291
rect	3	290	4	291
rect	4	290	5	291
rect	5	290	6	291
rect	7	290	8	291
rect	8	290	9	291
rect	9	290	10	291
rect	10	290	11	291
rect	11	290	12	291
rect	12	290	13	291
rect	13	290	14	291
rect	14	290	15	291
rect	15	290	16	291
rect	16	290	17	291
rect	17	290	18	291
rect	18	290	19	291
rect	19	290	20	291
rect	20	290	21	291
rect	21	290	22	291
rect	22	290	23	291
rect	23	290	24	291
rect	24	290	25	291
rect	25	290	26	291
rect	26	290	27	291
rect	27	290	28	291
rect	28	290	29	291
rect	29	290	30	291
rect	30	290	31	291
rect	32	290	33	291
rect	33	290	34	291
rect	34	290	35	291
rect	35	290	36	291
rect	36	290	37	291
rect	37	290	38	291
rect	38	290	39	291
rect	39	290	40	291
rect	40	290	41	291
rect	41	290	42	291
rect	42	290	43	291
rect	43	290	44	291
rect	44	290	45	291
rect	45	290	46	291
rect	46	290	47	291
rect	47	290	48	291
rect	48	290	49	291
rect	49	290	50	291
rect	50	290	51	291
rect	51	290	52	291
rect	52	290	53	291
rect	53	290	54	291
rect	54	290	55	291
rect	55	290	56	291
rect	56	290	57	291
rect	57	290	58	291
rect	58	290	59	291
rect	59	290	60	291
rect	60	290	61	291
rect	61	290	62	291
rect	62	290	63	291
rect	63	290	64	291
rect	64	290	65	291
rect	65	290	66	291
rect	66	290	67	291
rect	67	290	68	291
rect	68	290	69	291
rect	69	290	70	291
rect	70	290	71	291
rect	71	290	72	291
rect	72	290	73	291
rect	73	290	74	291
rect	74	290	75	291
rect	75	290	76	291
rect	76	290	77	291
rect	77	290	78	291
rect	78	290	79	291
rect	79	290	80	291
rect	80	290	81	291
rect	81	290	82	291
rect	82	290	83	291
rect	83	290	84	291
rect	84	290	85	291
rect	85	290	86	291
rect	86	290	87	291
rect	87	290	88	291
rect	88	290	89	291
rect	90	290	91	291
rect	91	290	92	291
rect	92	290	93	291
rect	93	290	94	291
rect	94	290	95	291
rect	95	290	96	291
rect	96	290	97	291
rect	97	290	98	291
rect	98	290	99	291
rect	99	290	100	291
rect	100	290	101	291
rect	101	290	102	291
rect	102	290	103	291
rect	103	290	104	291
rect	104	290	105	291
rect	105	290	106	291
rect	106	290	107	291
rect	107	290	108	291
rect	108	290	109	291
rect	109	290	110	291
rect	110	290	111	291
rect	111	290	112	291
rect	112	290	113	291
rect	113	290	114	291
rect	114	290	115	291
rect	115	290	116	291
rect	116	290	117	291
rect	117	290	118	291
rect	118	290	119	291
rect	119	290	120	291
rect	120	290	121	291
rect	121	290	122	291
rect	122	290	123	291
rect	123	290	124	291
rect	124	290	125	291
rect	125	290	126	291
rect	126	290	127	291
rect	127	290	128	291
rect	128	290	129	291
rect	129	290	130	291
rect	130	290	131	291
rect	131	290	132	291
rect	132	290	133	291
rect	133	290	134	291
rect	134	290	135	291
rect	135	290	136	291
rect	136	290	137	291
rect	137	290	138	291
rect	138	290	139	291
rect	139	290	140	291
rect	140	290	141	291
rect	141	290	142	291
rect	142	290	143	291
rect	143	290	144	291
rect	144	290	145	291
rect	145	290	146	291
rect	146	290	147	291
rect	147	290	148	291
rect	148	290	149	291
rect	149	290	150	291
rect	150	290	151	291
rect	151	290	152	291
rect	152	290	153	291
rect	153	290	154	291
rect	154	290	155	291
rect	155	290	156	291
rect	157	290	158	291
rect	158	290	159	291
rect	159	290	160	291
rect	160	290	161	291
rect	161	290	162	291
rect	162	290	163	291
rect	163	290	164	291
rect	164	290	165	291
rect	165	290	166	291
rect	166	290	167	291
rect	167	290	168	291
rect	168	290	169	291
rect	169	290	170	291
rect	170	290	171	291
rect	171	290	172	291
rect	172	290	173	291
rect	173	290	174	291
rect	174	290	175	291
rect	175	290	176	291
rect	176	290	177	291
rect	177	290	178	291
rect	178	290	179	291
rect	179	290	180	291
rect	180	290	181	291
rect	181	290	182	291
rect	182	290	183	291
rect	183	290	184	291
rect	184	290	185	291
rect	185	290	186	291
rect	186	290	187	291
rect	187	290	188	291
rect	188	290	189	291
rect	189	290	190	291
rect	190	290	191	291
rect	191	290	192	291
rect	192	290	193	291
rect	193	290	194	291
rect	194	290	195	291
rect	195	290	196	291
rect	196	290	197	291
rect	197	290	198	291
rect	198	290	199	291
rect	199	290	200	291
rect	200	290	201	291
rect	201	290	202	291
rect	202	290	203	291
rect	203	290	204	291
rect	204	290	205	291
rect	205	290	206	291
rect	206	290	207	291
rect	207	290	208	291
rect	208	290	209	291
rect	209	290	210	291
rect	210	290	211	291
rect	211	290	212	291
rect	212	290	213	291
rect	213	290	214	291
rect	214	290	215	291
rect	215	290	216	291
rect	216	290	217	291
rect	217	290	218	291
rect	218	290	219	291
rect	219	290	220	291
rect	220	290	221	291
rect	221	290	222	291
rect	222	290	223	291
rect	223	290	224	291
rect	224	290	225	291
rect	225	290	226	291
rect	226	290	227	291
rect	227	290	228	291
rect	228	290	229	291
rect	229	290	230	291
rect	230	290	231	291
rect	231	290	232	291
rect	232	290	233	291
rect	233	290	234	291
rect	234	290	235	291
rect	235	290	236	291
rect	236	290	237	291
rect	237	290	238	291
rect	239	290	240	291
rect	240	290	241	291
rect	241	290	242	291
rect	242	290	243	291
rect	243	290	244	291
rect	244	290	245	291
rect	245	290	246	291
rect	246	290	247	291
rect	247	290	248	291
rect	248	290	249	291
rect	249	290	250	291
rect	250	290	251	291
rect	251	290	252	291
rect	252	290	253	291
rect	253	290	254	291
rect	254	290	255	291
rect	255	290	256	291
rect	256	290	257	291
rect	257	290	258	291
rect	258	290	259	291
rect	259	290	260	291
rect	260	290	261	291
rect	261	290	262	291
rect	262	290	263	291
rect	264	290	265	291
rect	265	290	266	291
rect	266	290	267	291
rect	267	290	268	291
rect	268	290	269	291
rect	269	290	270	291
rect	270	290	271	291
rect	271	290	272	291
rect	272	290	273	291
rect	273	290	274	291
rect	274	290	275	291
rect	275	290	276	291
rect	276	290	277	291
rect	277	290	278	291
rect	278	290	279	291
rect	279	290	280	291
rect	280	290	281	291
rect	281	290	282	291
rect	282	290	283	291
rect	283	290	284	291
rect	284	290	285	291
rect	285	290	286	291
rect	286	290	287	291
rect	287	290	288	291
rect	288	290	289	291
rect	289	290	290	291
rect	290	290	291	291
rect	291	290	292	291
rect	292	290	293	291
rect	293	290	294	291
rect	294	290	295	291
rect	295	290	296	291
rect	296	290	297	291
rect	297	290	298	291
rect	298	290	299	291
rect	299	290	300	291
rect	301	290	302	291
rect	302	290	303	291
rect	303	290	304	291
rect	304	290	305	291
rect	305	290	306	291
rect	306	290	307	291
rect	307	290	308	291
rect	308	290	309	291
rect	309	290	310	291
rect	310	290	311	291
rect	311	290	312	291
rect	312	290	313	291
rect	313	290	314	291
rect	314	290	315	291
rect	315	290	316	291
rect	317	290	318	291
rect	318	290	319	291
rect	319	290	320	291
rect	320	290	321	291
rect	321	290	322	291
rect	322	290	323	291
rect	323	290	324	291
rect	324	290	325	291
rect	325	290	326	291
rect	326	290	327	291
rect	327	290	328	291
rect	328	290	329	291
rect	329	290	330	291
rect	330	290	331	291
rect	331	290	332	291
rect	332	290	333	291
rect	333	290	334	291
rect	334	290	335	291
rect	335	290	336	291
rect	336	290	337	291
rect	337	290	338	291
rect	338	290	339	291
rect	339	290	340	291
rect	340	290	341	291
rect	341	290	342	291
rect	342	290	343	291
rect	343	290	344	291
rect	344	290	345	291
rect	345	290	346	291
rect	346	290	347	291
rect	347	290	348	291
rect	348	290	349	291
rect	349	290	350	291
rect	350	290	351	291
rect	351	290	352	291
rect	352	290	353	291
rect	353	290	354	291
rect	354	290	355	291
rect	355	290	356	291
rect	356	290	357	291
rect	357	290	358	291
rect	358	290	359	291
rect	359	290	360	291
rect	360	290	361	291
rect	361	290	362	291
rect	362	290	363	291
rect	363	290	364	291
rect	364	290	365	291
rect	365	290	366	291
rect	366	290	367	291
rect	367	290	368	291
rect	368	290	369	291
rect	369	290	370	291
rect	370	290	371	291
rect	371	290	372	291
rect	372	290	373	291
rect	373	290	374	291
rect	374	290	375	291
rect	375	290	376	291
rect	376	290	377	291
rect	377	290	378	291
rect	378	290	379	291
rect	379	290	380	291
rect	380	290	381	291
rect	381	290	382	291
rect	382	290	383	291
rect	383	290	384	291
rect	384	290	385	291
rect	385	290	386	291
rect	386	290	387	291
rect	387	290	388	291
rect	388	290	389	291
rect	389	290	390	291
rect	390	290	391	291
rect	391	290	392	291
rect	392	290	393	291
rect	393	290	394	291
rect	394	290	395	291
rect	396	290	397	291
rect	397	290	398	291
rect	398	290	399	291
rect	399	290	400	291
rect	400	290	401	291
rect	401	290	402	291
rect	0	291	1	292
rect	1	291	2	292
rect	2	291	3	292
rect	3	291	4	292
rect	4	291	5	292
rect	5	291	6	292
rect	7	291	8	292
rect	8	291	9	292
rect	9	291	10	292
rect	10	291	11	292
rect	11	291	12	292
rect	12	291	13	292
rect	13	291	14	292
rect	14	291	15	292
rect	15	291	16	292
rect	16	291	17	292
rect	17	291	18	292
rect	18	291	19	292
rect	19	291	20	292
rect	20	291	21	292
rect	21	291	22	292
rect	22	291	23	292
rect	23	291	24	292
rect	24	291	25	292
rect	25	291	26	292
rect	26	291	27	292
rect	27	291	28	292
rect	28	291	29	292
rect	29	291	30	292
rect	30	291	31	292
rect	32	291	33	292
rect	33	291	34	292
rect	34	291	35	292
rect	35	291	36	292
rect	36	291	37	292
rect	37	291	38	292
rect	38	291	39	292
rect	39	291	40	292
rect	40	291	41	292
rect	41	291	42	292
rect	42	291	43	292
rect	43	291	44	292
rect	44	291	45	292
rect	45	291	46	292
rect	46	291	47	292
rect	47	291	48	292
rect	48	291	49	292
rect	49	291	50	292
rect	50	291	51	292
rect	51	291	52	292
rect	52	291	53	292
rect	53	291	54	292
rect	54	291	55	292
rect	55	291	56	292
rect	56	291	57	292
rect	57	291	58	292
rect	58	291	59	292
rect	59	291	60	292
rect	60	291	61	292
rect	61	291	62	292
rect	62	291	63	292
rect	63	291	64	292
rect	64	291	65	292
rect	65	291	66	292
rect	66	291	67	292
rect	67	291	68	292
rect	68	291	69	292
rect	69	291	70	292
rect	70	291	71	292
rect	71	291	72	292
rect	72	291	73	292
rect	73	291	74	292
rect	74	291	75	292
rect	75	291	76	292
rect	76	291	77	292
rect	77	291	78	292
rect	78	291	79	292
rect	79	291	80	292
rect	80	291	81	292
rect	81	291	82	292
rect	82	291	83	292
rect	83	291	84	292
rect	84	291	85	292
rect	85	291	86	292
rect	86	291	87	292
rect	87	291	88	292
rect	88	291	89	292
rect	90	291	91	292
rect	91	291	92	292
rect	92	291	93	292
rect	93	291	94	292
rect	94	291	95	292
rect	95	291	96	292
rect	96	291	97	292
rect	97	291	98	292
rect	98	291	99	292
rect	99	291	100	292
rect	100	291	101	292
rect	101	291	102	292
rect	102	291	103	292
rect	103	291	104	292
rect	104	291	105	292
rect	105	291	106	292
rect	106	291	107	292
rect	107	291	108	292
rect	108	291	109	292
rect	109	291	110	292
rect	110	291	111	292
rect	111	291	112	292
rect	112	291	113	292
rect	113	291	114	292
rect	114	291	115	292
rect	115	291	116	292
rect	116	291	117	292
rect	117	291	118	292
rect	118	291	119	292
rect	119	291	120	292
rect	120	291	121	292
rect	121	291	122	292
rect	122	291	123	292
rect	123	291	124	292
rect	124	291	125	292
rect	125	291	126	292
rect	126	291	127	292
rect	127	291	128	292
rect	128	291	129	292
rect	129	291	130	292
rect	130	291	131	292
rect	131	291	132	292
rect	132	291	133	292
rect	133	291	134	292
rect	134	291	135	292
rect	135	291	136	292
rect	136	291	137	292
rect	137	291	138	292
rect	138	291	139	292
rect	139	291	140	292
rect	140	291	141	292
rect	141	291	142	292
rect	142	291	143	292
rect	143	291	144	292
rect	144	291	145	292
rect	145	291	146	292
rect	146	291	147	292
rect	147	291	148	292
rect	148	291	149	292
rect	149	291	150	292
rect	150	291	151	292
rect	151	291	152	292
rect	152	291	153	292
rect	153	291	154	292
rect	154	291	155	292
rect	155	291	156	292
rect	157	291	158	292
rect	158	291	159	292
rect	159	291	160	292
rect	160	291	161	292
rect	161	291	162	292
rect	162	291	163	292
rect	163	291	164	292
rect	164	291	165	292
rect	165	291	166	292
rect	166	291	167	292
rect	167	291	168	292
rect	168	291	169	292
rect	169	291	170	292
rect	170	291	171	292
rect	171	291	172	292
rect	172	291	173	292
rect	173	291	174	292
rect	174	291	175	292
rect	175	291	176	292
rect	176	291	177	292
rect	177	291	178	292
rect	178	291	179	292
rect	179	291	180	292
rect	180	291	181	292
rect	181	291	182	292
rect	182	291	183	292
rect	183	291	184	292
rect	184	291	185	292
rect	185	291	186	292
rect	186	291	187	292
rect	187	291	188	292
rect	188	291	189	292
rect	189	291	190	292
rect	190	291	191	292
rect	191	291	192	292
rect	192	291	193	292
rect	193	291	194	292
rect	194	291	195	292
rect	195	291	196	292
rect	196	291	197	292
rect	197	291	198	292
rect	198	291	199	292
rect	199	291	200	292
rect	200	291	201	292
rect	201	291	202	292
rect	202	291	203	292
rect	203	291	204	292
rect	204	291	205	292
rect	205	291	206	292
rect	206	291	207	292
rect	207	291	208	292
rect	208	291	209	292
rect	209	291	210	292
rect	210	291	211	292
rect	211	291	212	292
rect	212	291	213	292
rect	213	291	214	292
rect	214	291	215	292
rect	215	291	216	292
rect	216	291	217	292
rect	217	291	218	292
rect	218	291	219	292
rect	219	291	220	292
rect	220	291	221	292
rect	221	291	222	292
rect	222	291	223	292
rect	223	291	224	292
rect	224	291	225	292
rect	225	291	226	292
rect	226	291	227	292
rect	227	291	228	292
rect	228	291	229	292
rect	229	291	230	292
rect	230	291	231	292
rect	231	291	232	292
rect	232	291	233	292
rect	233	291	234	292
rect	234	291	235	292
rect	235	291	236	292
rect	236	291	237	292
rect	237	291	238	292
rect	239	291	240	292
rect	240	291	241	292
rect	241	291	242	292
rect	242	291	243	292
rect	243	291	244	292
rect	244	291	245	292
rect	245	291	246	292
rect	246	291	247	292
rect	247	291	248	292
rect	248	291	249	292
rect	249	291	250	292
rect	250	291	251	292
rect	251	291	252	292
rect	252	291	253	292
rect	253	291	254	292
rect	254	291	255	292
rect	255	291	256	292
rect	256	291	257	292
rect	257	291	258	292
rect	258	291	259	292
rect	259	291	260	292
rect	260	291	261	292
rect	261	291	262	292
rect	262	291	263	292
rect	264	291	265	292
rect	265	291	266	292
rect	266	291	267	292
rect	267	291	268	292
rect	268	291	269	292
rect	269	291	270	292
rect	270	291	271	292
rect	271	291	272	292
rect	272	291	273	292
rect	273	291	274	292
rect	274	291	275	292
rect	275	291	276	292
rect	276	291	277	292
rect	277	291	278	292
rect	278	291	279	292
rect	279	291	280	292
rect	280	291	281	292
rect	281	291	282	292
rect	282	291	283	292
rect	283	291	284	292
rect	284	291	285	292
rect	285	291	286	292
rect	286	291	287	292
rect	287	291	288	292
rect	288	291	289	292
rect	289	291	290	292
rect	290	291	291	292
rect	291	291	292	292
rect	292	291	293	292
rect	293	291	294	292
rect	294	291	295	292
rect	295	291	296	292
rect	296	291	297	292
rect	297	291	298	292
rect	298	291	299	292
rect	299	291	300	292
rect	301	291	302	292
rect	302	291	303	292
rect	303	291	304	292
rect	304	291	305	292
rect	305	291	306	292
rect	306	291	307	292
rect	307	291	308	292
rect	308	291	309	292
rect	309	291	310	292
rect	310	291	311	292
rect	311	291	312	292
rect	312	291	313	292
rect	313	291	314	292
rect	314	291	315	292
rect	315	291	316	292
rect	317	291	318	292
rect	318	291	319	292
rect	319	291	320	292
rect	320	291	321	292
rect	321	291	322	292
rect	322	291	323	292
rect	323	291	324	292
rect	324	291	325	292
rect	325	291	326	292
rect	326	291	327	292
rect	327	291	328	292
rect	328	291	329	292
rect	329	291	330	292
rect	330	291	331	292
rect	331	291	332	292
rect	332	291	333	292
rect	333	291	334	292
rect	334	291	335	292
rect	335	291	336	292
rect	336	291	337	292
rect	337	291	338	292
rect	338	291	339	292
rect	339	291	340	292
rect	340	291	341	292
rect	341	291	342	292
rect	342	291	343	292
rect	343	291	344	292
rect	344	291	345	292
rect	345	291	346	292
rect	346	291	347	292
rect	347	291	348	292
rect	348	291	349	292
rect	349	291	350	292
rect	350	291	351	292
rect	351	291	352	292
rect	352	291	353	292
rect	353	291	354	292
rect	354	291	355	292
rect	355	291	356	292
rect	356	291	357	292
rect	357	291	358	292
rect	358	291	359	292
rect	359	291	360	292
rect	360	291	361	292
rect	361	291	362	292
rect	362	291	363	292
rect	363	291	364	292
rect	364	291	365	292
rect	365	291	366	292
rect	366	291	367	292
rect	367	291	368	292
rect	368	291	369	292
rect	369	291	370	292
rect	370	291	371	292
rect	371	291	372	292
rect	372	291	373	292
rect	373	291	374	292
rect	374	291	375	292
rect	375	291	376	292
rect	376	291	377	292
rect	377	291	378	292
rect	378	291	379	292
rect	379	291	380	292
rect	380	291	381	292
rect	381	291	382	292
rect	382	291	383	292
rect	383	291	384	292
rect	384	291	385	292
rect	385	291	386	292
rect	386	291	387	292
rect	387	291	388	292
rect	388	291	389	292
rect	389	291	390	292
rect	390	291	391	292
rect	391	291	392	292
rect	392	291	393	292
rect	393	291	394	292
rect	394	291	395	292
rect	396	291	397	292
rect	397	291	398	292
rect	398	291	399	292
rect	399	291	400	292
rect	400	291	401	292
rect	401	291	402	292
rect	0	292	1	293
rect	1	292	2	293
rect	2	292	3	293
rect	3	292	4	293
rect	4	292	5	293
rect	5	292	6	293
rect	7	292	8	293
rect	8	292	9	293
rect	9	292	10	293
rect	10	292	11	293
rect	11	292	12	293
rect	12	292	13	293
rect	13	292	14	293
rect	14	292	15	293
rect	15	292	16	293
rect	16	292	17	293
rect	17	292	18	293
rect	18	292	19	293
rect	19	292	20	293
rect	20	292	21	293
rect	21	292	22	293
rect	22	292	23	293
rect	23	292	24	293
rect	24	292	25	293
rect	25	292	26	293
rect	26	292	27	293
rect	27	292	28	293
rect	28	292	29	293
rect	29	292	30	293
rect	30	292	31	293
rect	32	292	33	293
rect	33	292	34	293
rect	34	292	35	293
rect	35	292	36	293
rect	36	292	37	293
rect	37	292	38	293
rect	38	292	39	293
rect	39	292	40	293
rect	40	292	41	293
rect	41	292	42	293
rect	42	292	43	293
rect	43	292	44	293
rect	44	292	45	293
rect	45	292	46	293
rect	46	292	47	293
rect	47	292	48	293
rect	48	292	49	293
rect	49	292	50	293
rect	50	292	51	293
rect	51	292	52	293
rect	52	292	53	293
rect	53	292	54	293
rect	54	292	55	293
rect	55	292	56	293
rect	56	292	57	293
rect	57	292	58	293
rect	58	292	59	293
rect	59	292	60	293
rect	60	292	61	293
rect	61	292	62	293
rect	62	292	63	293
rect	63	292	64	293
rect	64	292	65	293
rect	65	292	66	293
rect	66	292	67	293
rect	67	292	68	293
rect	68	292	69	293
rect	69	292	70	293
rect	70	292	71	293
rect	71	292	72	293
rect	72	292	73	293
rect	73	292	74	293
rect	74	292	75	293
rect	75	292	76	293
rect	76	292	77	293
rect	77	292	78	293
rect	78	292	79	293
rect	79	292	80	293
rect	80	292	81	293
rect	81	292	82	293
rect	82	292	83	293
rect	83	292	84	293
rect	84	292	85	293
rect	85	292	86	293
rect	86	292	87	293
rect	87	292	88	293
rect	88	292	89	293
rect	90	292	91	293
rect	91	292	92	293
rect	92	292	93	293
rect	93	292	94	293
rect	94	292	95	293
rect	95	292	96	293
rect	96	292	97	293
rect	97	292	98	293
rect	98	292	99	293
rect	99	292	100	293
rect	100	292	101	293
rect	101	292	102	293
rect	102	292	103	293
rect	103	292	104	293
rect	104	292	105	293
rect	105	292	106	293
rect	106	292	107	293
rect	107	292	108	293
rect	108	292	109	293
rect	109	292	110	293
rect	110	292	111	293
rect	111	292	112	293
rect	112	292	113	293
rect	113	292	114	293
rect	114	292	115	293
rect	115	292	116	293
rect	116	292	117	293
rect	117	292	118	293
rect	118	292	119	293
rect	119	292	120	293
rect	120	292	121	293
rect	121	292	122	293
rect	122	292	123	293
rect	123	292	124	293
rect	124	292	125	293
rect	125	292	126	293
rect	126	292	127	293
rect	127	292	128	293
rect	128	292	129	293
rect	129	292	130	293
rect	130	292	131	293
rect	131	292	132	293
rect	132	292	133	293
rect	133	292	134	293
rect	134	292	135	293
rect	135	292	136	293
rect	136	292	137	293
rect	137	292	138	293
rect	138	292	139	293
rect	139	292	140	293
rect	140	292	141	293
rect	141	292	142	293
rect	142	292	143	293
rect	143	292	144	293
rect	144	292	145	293
rect	145	292	146	293
rect	146	292	147	293
rect	147	292	148	293
rect	148	292	149	293
rect	149	292	150	293
rect	150	292	151	293
rect	151	292	152	293
rect	152	292	153	293
rect	153	292	154	293
rect	154	292	155	293
rect	155	292	156	293
rect	157	292	158	293
rect	158	292	159	293
rect	159	292	160	293
rect	160	292	161	293
rect	161	292	162	293
rect	162	292	163	293
rect	163	292	164	293
rect	164	292	165	293
rect	165	292	166	293
rect	166	292	167	293
rect	167	292	168	293
rect	168	292	169	293
rect	169	292	170	293
rect	170	292	171	293
rect	171	292	172	293
rect	172	292	173	293
rect	173	292	174	293
rect	174	292	175	293
rect	175	292	176	293
rect	176	292	177	293
rect	177	292	178	293
rect	178	292	179	293
rect	179	292	180	293
rect	180	292	181	293
rect	181	292	182	293
rect	182	292	183	293
rect	183	292	184	293
rect	184	292	185	293
rect	185	292	186	293
rect	186	292	187	293
rect	187	292	188	293
rect	188	292	189	293
rect	189	292	190	293
rect	190	292	191	293
rect	191	292	192	293
rect	192	292	193	293
rect	193	292	194	293
rect	194	292	195	293
rect	195	292	196	293
rect	196	292	197	293
rect	197	292	198	293
rect	198	292	199	293
rect	199	292	200	293
rect	200	292	201	293
rect	201	292	202	293
rect	202	292	203	293
rect	203	292	204	293
rect	204	292	205	293
rect	205	292	206	293
rect	206	292	207	293
rect	207	292	208	293
rect	208	292	209	293
rect	209	292	210	293
rect	210	292	211	293
rect	211	292	212	293
rect	212	292	213	293
rect	213	292	214	293
rect	214	292	215	293
rect	215	292	216	293
rect	216	292	217	293
rect	217	292	218	293
rect	218	292	219	293
rect	219	292	220	293
rect	220	292	221	293
rect	221	292	222	293
rect	222	292	223	293
rect	223	292	224	293
rect	224	292	225	293
rect	225	292	226	293
rect	226	292	227	293
rect	227	292	228	293
rect	228	292	229	293
rect	229	292	230	293
rect	230	292	231	293
rect	231	292	232	293
rect	232	292	233	293
rect	233	292	234	293
rect	234	292	235	293
rect	235	292	236	293
rect	236	292	237	293
rect	237	292	238	293
rect	239	292	240	293
rect	240	292	241	293
rect	241	292	242	293
rect	242	292	243	293
rect	243	292	244	293
rect	244	292	245	293
rect	245	292	246	293
rect	246	292	247	293
rect	247	292	248	293
rect	248	292	249	293
rect	249	292	250	293
rect	250	292	251	293
rect	251	292	252	293
rect	252	292	253	293
rect	253	292	254	293
rect	254	292	255	293
rect	255	292	256	293
rect	256	292	257	293
rect	257	292	258	293
rect	258	292	259	293
rect	259	292	260	293
rect	260	292	261	293
rect	261	292	262	293
rect	262	292	263	293
rect	264	292	265	293
rect	265	292	266	293
rect	266	292	267	293
rect	267	292	268	293
rect	268	292	269	293
rect	269	292	270	293
rect	270	292	271	293
rect	271	292	272	293
rect	272	292	273	293
rect	273	292	274	293
rect	274	292	275	293
rect	275	292	276	293
rect	276	292	277	293
rect	277	292	278	293
rect	278	292	279	293
rect	279	292	280	293
rect	280	292	281	293
rect	281	292	282	293
rect	282	292	283	293
rect	283	292	284	293
rect	284	292	285	293
rect	285	292	286	293
rect	286	292	287	293
rect	287	292	288	293
rect	288	292	289	293
rect	289	292	290	293
rect	290	292	291	293
rect	291	292	292	293
rect	292	292	293	293
rect	293	292	294	293
rect	294	292	295	293
rect	295	292	296	293
rect	296	292	297	293
rect	297	292	298	293
rect	298	292	299	293
rect	299	292	300	293
rect	301	292	302	293
rect	302	292	303	293
rect	303	292	304	293
rect	304	292	305	293
rect	305	292	306	293
rect	306	292	307	293
rect	307	292	308	293
rect	308	292	309	293
rect	309	292	310	293
rect	310	292	311	293
rect	311	292	312	293
rect	312	292	313	293
rect	313	292	314	293
rect	314	292	315	293
rect	315	292	316	293
rect	317	292	318	293
rect	318	292	319	293
rect	319	292	320	293
rect	320	292	321	293
rect	321	292	322	293
rect	322	292	323	293
rect	323	292	324	293
rect	324	292	325	293
rect	325	292	326	293
rect	326	292	327	293
rect	327	292	328	293
rect	328	292	329	293
rect	329	292	330	293
rect	330	292	331	293
rect	331	292	332	293
rect	332	292	333	293
rect	333	292	334	293
rect	334	292	335	293
rect	335	292	336	293
rect	336	292	337	293
rect	337	292	338	293
rect	338	292	339	293
rect	339	292	340	293
rect	340	292	341	293
rect	341	292	342	293
rect	342	292	343	293
rect	343	292	344	293
rect	344	292	345	293
rect	345	292	346	293
rect	346	292	347	293
rect	347	292	348	293
rect	348	292	349	293
rect	349	292	350	293
rect	350	292	351	293
rect	351	292	352	293
rect	352	292	353	293
rect	353	292	354	293
rect	354	292	355	293
rect	355	292	356	293
rect	356	292	357	293
rect	357	292	358	293
rect	358	292	359	293
rect	359	292	360	293
rect	360	292	361	293
rect	361	292	362	293
rect	362	292	363	293
rect	363	292	364	293
rect	364	292	365	293
rect	365	292	366	293
rect	366	292	367	293
rect	367	292	368	293
rect	368	292	369	293
rect	369	292	370	293
rect	370	292	371	293
rect	371	292	372	293
rect	372	292	373	293
rect	373	292	374	293
rect	374	292	375	293
rect	375	292	376	293
rect	376	292	377	293
rect	377	292	378	293
rect	378	292	379	293
rect	379	292	380	293
rect	380	292	381	293
rect	381	292	382	293
rect	382	292	383	293
rect	383	292	384	293
rect	384	292	385	293
rect	385	292	386	293
rect	386	292	387	293
rect	387	292	388	293
rect	388	292	389	293
rect	389	292	390	293
rect	390	292	391	293
rect	391	292	392	293
rect	392	292	393	293
rect	393	292	394	293
rect	394	292	395	293
rect	396	292	397	293
rect	397	292	398	293
rect	398	292	399	293
rect	399	292	400	293
rect	400	292	401	293
rect	401	292	402	293
rect	0	293	1	294
rect	1	293	2	294
rect	2	293	3	294
rect	3	293	4	294
rect	4	293	5	294
rect	5	293	6	294
rect	7	293	8	294
rect	8	293	9	294
rect	9	293	10	294
rect	10	293	11	294
rect	11	293	12	294
rect	12	293	13	294
rect	13	293	14	294
rect	14	293	15	294
rect	15	293	16	294
rect	16	293	17	294
rect	17	293	18	294
rect	18	293	19	294
rect	19	293	20	294
rect	20	293	21	294
rect	21	293	22	294
rect	22	293	23	294
rect	23	293	24	294
rect	24	293	25	294
rect	25	293	26	294
rect	26	293	27	294
rect	27	293	28	294
rect	28	293	29	294
rect	29	293	30	294
rect	30	293	31	294
rect	32	293	33	294
rect	33	293	34	294
rect	34	293	35	294
rect	35	293	36	294
rect	36	293	37	294
rect	37	293	38	294
rect	38	293	39	294
rect	39	293	40	294
rect	40	293	41	294
rect	41	293	42	294
rect	42	293	43	294
rect	43	293	44	294
rect	44	293	45	294
rect	45	293	46	294
rect	46	293	47	294
rect	47	293	48	294
rect	48	293	49	294
rect	49	293	50	294
rect	50	293	51	294
rect	51	293	52	294
rect	52	293	53	294
rect	53	293	54	294
rect	54	293	55	294
rect	55	293	56	294
rect	56	293	57	294
rect	57	293	58	294
rect	58	293	59	294
rect	59	293	60	294
rect	60	293	61	294
rect	61	293	62	294
rect	62	293	63	294
rect	63	293	64	294
rect	64	293	65	294
rect	65	293	66	294
rect	66	293	67	294
rect	67	293	68	294
rect	68	293	69	294
rect	69	293	70	294
rect	70	293	71	294
rect	71	293	72	294
rect	72	293	73	294
rect	73	293	74	294
rect	74	293	75	294
rect	75	293	76	294
rect	76	293	77	294
rect	77	293	78	294
rect	78	293	79	294
rect	79	293	80	294
rect	80	293	81	294
rect	81	293	82	294
rect	82	293	83	294
rect	83	293	84	294
rect	84	293	85	294
rect	85	293	86	294
rect	86	293	87	294
rect	87	293	88	294
rect	88	293	89	294
rect	90	293	91	294
rect	91	293	92	294
rect	92	293	93	294
rect	93	293	94	294
rect	94	293	95	294
rect	95	293	96	294
rect	96	293	97	294
rect	97	293	98	294
rect	98	293	99	294
rect	99	293	100	294
rect	100	293	101	294
rect	101	293	102	294
rect	102	293	103	294
rect	103	293	104	294
rect	104	293	105	294
rect	105	293	106	294
rect	106	293	107	294
rect	107	293	108	294
rect	108	293	109	294
rect	109	293	110	294
rect	110	293	111	294
rect	111	293	112	294
rect	112	293	113	294
rect	113	293	114	294
rect	114	293	115	294
rect	115	293	116	294
rect	116	293	117	294
rect	117	293	118	294
rect	118	293	119	294
rect	119	293	120	294
rect	120	293	121	294
rect	121	293	122	294
rect	122	293	123	294
rect	123	293	124	294
rect	124	293	125	294
rect	125	293	126	294
rect	126	293	127	294
rect	127	293	128	294
rect	128	293	129	294
rect	129	293	130	294
rect	130	293	131	294
rect	131	293	132	294
rect	132	293	133	294
rect	133	293	134	294
rect	134	293	135	294
rect	135	293	136	294
rect	136	293	137	294
rect	137	293	138	294
rect	138	293	139	294
rect	139	293	140	294
rect	140	293	141	294
rect	141	293	142	294
rect	142	293	143	294
rect	143	293	144	294
rect	144	293	145	294
rect	145	293	146	294
rect	146	293	147	294
rect	147	293	148	294
rect	148	293	149	294
rect	149	293	150	294
rect	150	293	151	294
rect	151	293	152	294
rect	152	293	153	294
rect	153	293	154	294
rect	154	293	155	294
rect	155	293	156	294
rect	157	293	158	294
rect	158	293	159	294
rect	159	293	160	294
rect	160	293	161	294
rect	161	293	162	294
rect	162	293	163	294
rect	163	293	164	294
rect	164	293	165	294
rect	165	293	166	294
rect	166	293	167	294
rect	167	293	168	294
rect	168	293	169	294
rect	169	293	170	294
rect	170	293	171	294
rect	171	293	172	294
rect	172	293	173	294
rect	173	293	174	294
rect	174	293	175	294
rect	175	293	176	294
rect	176	293	177	294
rect	177	293	178	294
rect	178	293	179	294
rect	179	293	180	294
rect	180	293	181	294
rect	181	293	182	294
rect	182	293	183	294
rect	183	293	184	294
rect	184	293	185	294
rect	185	293	186	294
rect	186	293	187	294
rect	187	293	188	294
rect	188	293	189	294
rect	189	293	190	294
rect	190	293	191	294
rect	191	293	192	294
rect	192	293	193	294
rect	193	293	194	294
rect	194	293	195	294
rect	195	293	196	294
rect	196	293	197	294
rect	197	293	198	294
rect	198	293	199	294
rect	199	293	200	294
rect	200	293	201	294
rect	201	293	202	294
rect	202	293	203	294
rect	203	293	204	294
rect	204	293	205	294
rect	205	293	206	294
rect	206	293	207	294
rect	207	293	208	294
rect	208	293	209	294
rect	209	293	210	294
rect	210	293	211	294
rect	211	293	212	294
rect	212	293	213	294
rect	213	293	214	294
rect	214	293	215	294
rect	215	293	216	294
rect	216	293	217	294
rect	217	293	218	294
rect	218	293	219	294
rect	219	293	220	294
rect	220	293	221	294
rect	221	293	222	294
rect	222	293	223	294
rect	223	293	224	294
rect	224	293	225	294
rect	225	293	226	294
rect	226	293	227	294
rect	227	293	228	294
rect	228	293	229	294
rect	229	293	230	294
rect	230	293	231	294
rect	231	293	232	294
rect	232	293	233	294
rect	233	293	234	294
rect	234	293	235	294
rect	235	293	236	294
rect	236	293	237	294
rect	237	293	238	294
rect	239	293	240	294
rect	240	293	241	294
rect	241	293	242	294
rect	242	293	243	294
rect	243	293	244	294
rect	244	293	245	294
rect	245	293	246	294
rect	246	293	247	294
rect	247	293	248	294
rect	248	293	249	294
rect	249	293	250	294
rect	250	293	251	294
rect	251	293	252	294
rect	252	293	253	294
rect	253	293	254	294
rect	254	293	255	294
rect	255	293	256	294
rect	256	293	257	294
rect	257	293	258	294
rect	258	293	259	294
rect	259	293	260	294
rect	260	293	261	294
rect	261	293	262	294
rect	262	293	263	294
rect	264	293	265	294
rect	265	293	266	294
rect	266	293	267	294
rect	267	293	268	294
rect	268	293	269	294
rect	269	293	270	294
rect	270	293	271	294
rect	271	293	272	294
rect	272	293	273	294
rect	273	293	274	294
rect	274	293	275	294
rect	275	293	276	294
rect	276	293	277	294
rect	277	293	278	294
rect	278	293	279	294
rect	279	293	280	294
rect	280	293	281	294
rect	281	293	282	294
rect	282	293	283	294
rect	283	293	284	294
rect	284	293	285	294
rect	285	293	286	294
rect	286	293	287	294
rect	287	293	288	294
rect	288	293	289	294
rect	289	293	290	294
rect	290	293	291	294
rect	291	293	292	294
rect	292	293	293	294
rect	293	293	294	294
rect	294	293	295	294
rect	295	293	296	294
rect	296	293	297	294
rect	297	293	298	294
rect	298	293	299	294
rect	299	293	300	294
rect	301	293	302	294
rect	302	293	303	294
rect	303	293	304	294
rect	304	293	305	294
rect	305	293	306	294
rect	306	293	307	294
rect	307	293	308	294
rect	308	293	309	294
rect	309	293	310	294
rect	310	293	311	294
rect	311	293	312	294
rect	312	293	313	294
rect	313	293	314	294
rect	314	293	315	294
rect	315	293	316	294
rect	317	293	318	294
rect	318	293	319	294
rect	319	293	320	294
rect	320	293	321	294
rect	321	293	322	294
rect	322	293	323	294
rect	323	293	324	294
rect	324	293	325	294
rect	325	293	326	294
rect	326	293	327	294
rect	327	293	328	294
rect	328	293	329	294
rect	329	293	330	294
rect	330	293	331	294
rect	331	293	332	294
rect	332	293	333	294
rect	333	293	334	294
rect	334	293	335	294
rect	335	293	336	294
rect	336	293	337	294
rect	337	293	338	294
rect	338	293	339	294
rect	339	293	340	294
rect	340	293	341	294
rect	341	293	342	294
rect	342	293	343	294
rect	343	293	344	294
rect	344	293	345	294
rect	345	293	346	294
rect	346	293	347	294
rect	347	293	348	294
rect	348	293	349	294
rect	349	293	350	294
rect	350	293	351	294
rect	351	293	352	294
rect	352	293	353	294
rect	353	293	354	294
rect	354	293	355	294
rect	355	293	356	294
rect	356	293	357	294
rect	357	293	358	294
rect	358	293	359	294
rect	359	293	360	294
rect	360	293	361	294
rect	361	293	362	294
rect	362	293	363	294
rect	363	293	364	294
rect	364	293	365	294
rect	365	293	366	294
rect	366	293	367	294
rect	367	293	368	294
rect	368	293	369	294
rect	369	293	370	294
rect	370	293	371	294
rect	371	293	372	294
rect	372	293	373	294
rect	373	293	374	294
rect	374	293	375	294
rect	375	293	376	294
rect	376	293	377	294
rect	377	293	378	294
rect	378	293	379	294
rect	379	293	380	294
rect	380	293	381	294
rect	381	293	382	294
rect	382	293	383	294
rect	383	293	384	294
rect	384	293	385	294
rect	385	293	386	294
rect	386	293	387	294
rect	387	293	388	294
rect	388	293	389	294
rect	389	293	390	294
rect	390	293	391	294
rect	391	293	392	294
rect	392	293	393	294
rect	393	293	394	294
rect	394	293	395	294
rect	396	293	397	294
rect	397	293	398	294
rect	398	293	399	294
rect	399	293	400	294
rect	400	293	401	294
rect	401	293	402	294
rect	0	294	1	295
rect	1	294	2	295
rect	2	294	3	295
rect	3	294	4	295
rect	4	294	5	295
rect	5	294	6	295
rect	7	294	8	295
rect	8	294	9	295
rect	9	294	10	295
rect	10	294	11	295
rect	11	294	12	295
rect	12	294	13	295
rect	13	294	14	295
rect	14	294	15	295
rect	15	294	16	295
rect	16	294	17	295
rect	17	294	18	295
rect	18	294	19	295
rect	19	294	20	295
rect	20	294	21	295
rect	21	294	22	295
rect	22	294	23	295
rect	23	294	24	295
rect	24	294	25	295
rect	25	294	26	295
rect	26	294	27	295
rect	27	294	28	295
rect	28	294	29	295
rect	29	294	30	295
rect	30	294	31	295
rect	32	294	33	295
rect	33	294	34	295
rect	34	294	35	295
rect	35	294	36	295
rect	36	294	37	295
rect	37	294	38	295
rect	38	294	39	295
rect	39	294	40	295
rect	40	294	41	295
rect	41	294	42	295
rect	42	294	43	295
rect	43	294	44	295
rect	44	294	45	295
rect	45	294	46	295
rect	46	294	47	295
rect	47	294	48	295
rect	48	294	49	295
rect	49	294	50	295
rect	50	294	51	295
rect	51	294	52	295
rect	52	294	53	295
rect	53	294	54	295
rect	54	294	55	295
rect	55	294	56	295
rect	56	294	57	295
rect	57	294	58	295
rect	58	294	59	295
rect	59	294	60	295
rect	60	294	61	295
rect	61	294	62	295
rect	62	294	63	295
rect	63	294	64	295
rect	64	294	65	295
rect	65	294	66	295
rect	66	294	67	295
rect	67	294	68	295
rect	68	294	69	295
rect	69	294	70	295
rect	70	294	71	295
rect	71	294	72	295
rect	72	294	73	295
rect	73	294	74	295
rect	74	294	75	295
rect	75	294	76	295
rect	76	294	77	295
rect	77	294	78	295
rect	78	294	79	295
rect	79	294	80	295
rect	80	294	81	295
rect	81	294	82	295
rect	82	294	83	295
rect	83	294	84	295
rect	84	294	85	295
rect	85	294	86	295
rect	86	294	87	295
rect	87	294	88	295
rect	88	294	89	295
rect	90	294	91	295
rect	91	294	92	295
rect	92	294	93	295
rect	93	294	94	295
rect	94	294	95	295
rect	95	294	96	295
rect	96	294	97	295
rect	97	294	98	295
rect	98	294	99	295
rect	99	294	100	295
rect	100	294	101	295
rect	101	294	102	295
rect	102	294	103	295
rect	103	294	104	295
rect	104	294	105	295
rect	105	294	106	295
rect	106	294	107	295
rect	107	294	108	295
rect	108	294	109	295
rect	109	294	110	295
rect	110	294	111	295
rect	111	294	112	295
rect	112	294	113	295
rect	113	294	114	295
rect	114	294	115	295
rect	115	294	116	295
rect	116	294	117	295
rect	117	294	118	295
rect	118	294	119	295
rect	119	294	120	295
rect	120	294	121	295
rect	121	294	122	295
rect	122	294	123	295
rect	123	294	124	295
rect	124	294	125	295
rect	125	294	126	295
rect	126	294	127	295
rect	127	294	128	295
rect	128	294	129	295
rect	129	294	130	295
rect	130	294	131	295
rect	131	294	132	295
rect	132	294	133	295
rect	133	294	134	295
rect	134	294	135	295
rect	135	294	136	295
rect	136	294	137	295
rect	137	294	138	295
rect	138	294	139	295
rect	139	294	140	295
rect	140	294	141	295
rect	141	294	142	295
rect	142	294	143	295
rect	143	294	144	295
rect	144	294	145	295
rect	145	294	146	295
rect	146	294	147	295
rect	147	294	148	295
rect	148	294	149	295
rect	149	294	150	295
rect	150	294	151	295
rect	151	294	152	295
rect	152	294	153	295
rect	153	294	154	295
rect	154	294	155	295
rect	155	294	156	295
rect	157	294	158	295
rect	158	294	159	295
rect	159	294	160	295
rect	160	294	161	295
rect	161	294	162	295
rect	162	294	163	295
rect	163	294	164	295
rect	164	294	165	295
rect	165	294	166	295
rect	166	294	167	295
rect	167	294	168	295
rect	168	294	169	295
rect	169	294	170	295
rect	170	294	171	295
rect	171	294	172	295
rect	172	294	173	295
rect	173	294	174	295
rect	174	294	175	295
rect	175	294	176	295
rect	176	294	177	295
rect	177	294	178	295
rect	178	294	179	295
rect	179	294	180	295
rect	180	294	181	295
rect	181	294	182	295
rect	182	294	183	295
rect	183	294	184	295
rect	184	294	185	295
rect	185	294	186	295
rect	186	294	187	295
rect	187	294	188	295
rect	188	294	189	295
rect	189	294	190	295
rect	190	294	191	295
rect	191	294	192	295
rect	192	294	193	295
rect	193	294	194	295
rect	194	294	195	295
rect	195	294	196	295
rect	196	294	197	295
rect	197	294	198	295
rect	198	294	199	295
rect	199	294	200	295
rect	200	294	201	295
rect	201	294	202	295
rect	202	294	203	295
rect	203	294	204	295
rect	204	294	205	295
rect	205	294	206	295
rect	206	294	207	295
rect	207	294	208	295
rect	208	294	209	295
rect	209	294	210	295
rect	210	294	211	295
rect	211	294	212	295
rect	212	294	213	295
rect	213	294	214	295
rect	214	294	215	295
rect	215	294	216	295
rect	216	294	217	295
rect	217	294	218	295
rect	218	294	219	295
rect	219	294	220	295
rect	220	294	221	295
rect	221	294	222	295
rect	222	294	223	295
rect	223	294	224	295
rect	224	294	225	295
rect	225	294	226	295
rect	226	294	227	295
rect	227	294	228	295
rect	228	294	229	295
rect	229	294	230	295
rect	230	294	231	295
rect	231	294	232	295
rect	232	294	233	295
rect	233	294	234	295
rect	234	294	235	295
rect	235	294	236	295
rect	236	294	237	295
rect	237	294	238	295
rect	239	294	240	295
rect	240	294	241	295
rect	241	294	242	295
rect	242	294	243	295
rect	243	294	244	295
rect	244	294	245	295
rect	245	294	246	295
rect	246	294	247	295
rect	247	294	248	295
rect	248	294	249	295
rect	249	294	250	295
rect	250	294	251	295
rect	251	294	252	295
rect	252	294	253	295
rect	253	294	254	295
rect	254	294	255	295
rect	255	294	256	295
rect	256	294	257	295
rect	257	294	258	295
rect	258	294	259	295
rect	259	294	260	295
rect	260	294	261	295
rect	261	294	262	295
rect	262	294	263	295
rect	264	294	265	295
rect	265	294	266	295
rect	266	294	267	295
rect	267	294	268	295
rect	268	294	269	295
rect	269	294	270	295
rect	270	294	271	295
rect	271	294	272	295
rect	272	294	273	295
rect	273	294	274	295
rect	274	294	275	295
rect	275	294	276	295
rect	276	294	277	295
rect	277	294	278	295
rect	278	294	279	295
rect	279	294	280	295
rect	280	294	281	295
rect	281	294	282	295
rect	282	294	283	295
rect	283	294	284	295
rect	284	294	285	295
rect	285	294	286	295
rect	286	294	287	295
rect	287	294	288	295
rect	288	294	289	295
rect	289	294	290	295
rect	290	294	291	295
rect	291	294	292	295
rect	292	294	293	295
rect	293	294	294	295
rect	294	294	295	295
rect	295	294	296	295
rect	296	294	297	295
rect	297	294	298	295
rect	298	294	299	295
rect	299	294	300	295
rect	301	294	302	295
rect	302	294	303	295
rect	303	294	304	295
rect	304	294	305	295
rect	305	294	306	295
rect	306	294	307	295
rect	307	294	308	295
rect	308	294	309	295
rect	309	294	310	295
rect	310	294	311	295
rect	311	294	312	295
rect	312	294	313	295
rect	313	294	314	295
rect	314	294	315	295
rect	315	294	316	295
rect	317	294	318	295
rect	318	294	319	295
rect	319	294	320	295
rect	320	294	321	295
rect	321	294	322	295
rect	322	294	323	295
rect	323	294	324	295
rect	324	294	325	295
rect	325	294	326	295
rect	326	294	327	295
rect	327	294	328	295
rect	328	294	329	295
rect	329	294	330	295
rect	330	294	331	295
rect	331	294	332	295
rect	332	294	333	295
rect	333	294	334	295
rect	334	294	335	295
rect	335	294	336	295
rect	336	294	337	295
rect	337	294	338	295
rect	338	294	339	295
rect	339	294	340	295
rect	340	294	341	295
rect	341	294	342	295
rect	342	294	343	295
rect	343	294	344	295
rect	344	294	345	295
rect	345	294	346	295
rect	346	294	347	295
rect	347	294	348	295
rect	348	294	349	295
rect	349	294	350	295
rect	350	294	351	295
rect	351	294	352	295
rect	352	294	353	295
rect	353	294	354	295
rect	354	294	355	295
rect	355	294	356	295
rect	356	294	357	295
rect	357	294	358	295
rect	358	294	359	295
rect	359	294	360	295
rect	360	294	361	295
rect	361	294	362	295
rect	362	294	363	295
rect	363	294	364	295
rect	364	294	365	295
rect	365	294	366	295
rect	366	294	367	295
rect	367	294	368	295
rect	368	294	369	295
rect	369	294	370	295
rect	370	294	371	295
rect	371	294	372	295
rect	372	294	373	295
rect	373	294	374	295
rect	374	294	375	295
rect	375	294	376	295
rect	376	294	377	295
rect	377	294	378	295
rect	378	294	379	295
rect	379	294	380	295
rect	380	294	381	295
rect	381	294	382	295
rect	382	294	383	295
rect	383	294	384	295
rect	384	294	385	295
rect	385	294	386	295
rect	386	294	387	295
rect	387	294	388	295
rect	388	294	389	295
rect	389	294	390	295
rect	390	294	391	295
rect	391	294	392	295
rect	392	294	393	295
rect	393	294	394	295
rect	394	294	395	295
rect	396	294	397	295
rect	397	294	398	295
rect	398	294	399	295
rect	399	294	400	295
rect	400	294	401	295
rect	401	294	402	295
rect	0	295	1	296
rect	1	295	2	296
rect	2	295	3	296
rect	3	295	4	296
rect	4	295	5	296
rect	5	295	6	296
rect	7	295	8	296
rect	8	295	9	296
rect	9	295	10	296
rect	10	295	11	296
rect	11	295	12	296
rect	12	295	13	296
rect	13	295	14	296
rect	14	295	15	296
rect	15	295	16	296
rect	16	295	17	296
rect	17	295	18	296
rect	18	295	19	296
rect	19	295	20	296
rect	20	295	21	296
rect	21	295	22	296
rect	22	295	23	296
rect	23	295	24	296
rect	24	295	25	296
rect	25	295	26	296
rect	26	295	27	296
rect	27	295	28	296
rect	28	295	29	296
rect	29	295	30	296
rect	30	295	31	296
rect	32	295	33	296
rect	33	295	34	296
rect	34	295	35	296
rect	35	295	36	296
rect	36	295	37	296
rect	37	295	38	296
rect	38	295	39	296
rect	39	295	40	296
rect	40	295	41	296
rect	41	295	42	296
rect	42	295	43	296
rect	43	295	44	296
rect	44	295	45	296
rect	45	295	46	296
rect	46	295	47	296
rect	47	295	48	296
rect	48	295	49	296
rect	49	295	50	296
rect	50	295	51	296
rect	51	295	52	296
rect	52	295	53	296
rect	53	295	54	296
rect	54	295	55	296
rect	55	295	56	296
rect	56	295	57	296
rect	57	295	58	296
rect	58	295	59	296
rect	59	295	60	296
rect	60	295	61	296
rect	61	295	62	296
rect	62	295	63	296
rect	63	295	64	296
rect	64	295	65	296
rect	65	295	66	296
rect	66	295	67	296
rect	67	295	68	296
rect	68	295	69	296
rect	69	295	70	296
rect	70	295	71	296
rect	71	295	72	296
rect	72	295	73	296
rect	73	295	74	296
rect	74	295	75	296
rect	75	295	76	296
rect	76	295	77	296
rect	77	295	78	296
rect	78	295	79	296
rect	79	295	80	296
rect	80	295	81	296
rect	81	295	82	296
rect	82	295	83	296
rect	83	295	84	296
rect	84	295	85	296
rect	85	295	86	296
rect	86	295	87	296
rect	87	295	88	296
rect	88	295	89	296
rect	90	295	91	296
rect	91	295	92	296
rect	92	295	93	296
rect	93	295	94	296
rect	94	295	95	296
rect	95	295	96	296
rect	96	295	97	296
rect	97	295	98	296
rect	98	295	99	296
rect	99	295	100	296
rect	100	295	101	296
rect	101	295	102	296
rect	102	295	103	296
rect	103	295	104	296
rect	104	295	105	296
rect	105	295	106	296
rect	106	295	107	296
rect	107	295	108	296
rect	108	295	109	296
rect	109	295	110	296
rect	110	295	111	296
rect	111	295	112	296
rect	112	295	113	296
rect	113	295	114	296
rect	114	295	115	296
rect	115	295	116	296
rect	116	295	117	296
rect	117	295	118	296
rect	118	295	119	296
rect	119	295	120	296
rect	120	295	121	296
rect	121	295	122	296
rect	122	295	123	296
rect	123	295	124	296
rect	124	295	125	296
rect	125	295	126	296
rect	126	295	127	296
rect	127	295	128	296
rect	128	295	129	296
rect	129	295	130	296
rect	130	295	131	296
rect	131	295	132	296
rect	132	295	133	296
rect	133	295	134	296
rect	134	295	135	296
rect	135	295	136	296
rect	136	295	137	296
rect	137	295	138	296
rect	138	295	139	296
rect	139	295	140	296
rect	140	295	141	296
rect	141	295	142	296
rect	142	295	143	296
rect	143	295	144	296
rect	144	295	145	296
rect	145	295	146	296
rect	146	295	147	296
rect	147	295	148	296
rect	148	295	149	296
rect	149	295	150	296
rect	150	295	151	296
rect	151	295	152	296
rect	152	295	153	296
rect	153	295	154	296
rect	154	295	155	296
rect	155	295	156	296
rect	157	295	158	296
rect	158	295	159	296
rect	159	295	160	296
rect	160	295	161	296
rect	161	295	162	296
rect	162	295	163	296
rect	163	295	164	296
rect	164	295	165	296
rect	165	295	166	296
rect	166	295	167	296
rect	167	295	168	296
rect	168	295	169	296
rect	169	295	170	296
rect	170	295	171	296
rect	171	295	172	296
rect	172	295	173	296
rect	173	295	174	296
rect	174	295	175	296
rect	175	295	176	296
rect	176	295	177	296
rect	177	295	178	296
rect	178	295	179	296
rect	179	295	180	296
rect	180	295	181	296
rect	181	295	182	296
rect	182	295	183	296
rect	183	295	184	296
rect	184	295	185	296
rect	185	295	186	296
rect	186	295	187	296
rect	187	295	188	296
rect	188	295	189	296
rect	189	295	190	296
rect	190	295	191	296
rect	191	295	192	296
rect	192	295	193	296
rect	193	295	194	296
rect	194	295	195	296
rect	195	295	196	296
rect	196	295	197	296
rect	197	295	198	296
rect	198	295	199	296
rect	199	295	200	296
rect	200	295	201	296
rect	201	295	202	296
rect	202	295	203	296
rect	203	295	204	296
rect	204	295	205	296
rect	205	295	206	296
rect	206	295	207	296
rect	207	295	208	296
rect	208	295	209	296
rect	209	295	210	296
rect	210	295	211	296
rect	211	295	212	296
rect	212	295	213	296
rect	213	295	214	296
rect	214	295	215	296
rect	215	295	216	296
rect	216	295	217	296
rect	217	295	218	296
rect	218	295	219	296
rect	219	295	220	296
rect	220	295	221	296
rect	221	295	222	296
rect	222	295	223	296
rect	223	295	224	296
rect	224	295	225	296
rect	225	295	226	296
rect	226	295	227	296
rect	227	295	228	296
rect	228	295	229	296
rect	229	295	230	296
rect	230	295	231	296
rect	231	295	232	296
rect	232	295	233	296
rect	233	295	234	296
rect	234	295	235	296
rect	235	295	236	296
rect	236	295	237	296
rect	237	295	238	296
rect	239	295	240	296
rect	240	295	241	296
rect	241	295	242	296
rect	242	295	243	296
rect	243	295	244	296
rect	244	295	245	296
rect	245	295	246	296
rect	246	295	247	296
rect	247	295	248	296
rect	248	295	249	296
rect	249	295	250	296
rect	250	295	251	296
rect	251	295	252	296
rect	252	295	253	296
rect	253	295	254	296
rect	254	295	255	296
rect	255	295	256	296
rect	256	295	257	296
rect	257	295	258	296
rect	258	295	259	296
rect	259	295	260	296
rect	260	295	261	296
rect	261	295	262	296
rect	262	295	263	296
rect	264	295	265	296
rect	265	295	266	296
rect	266	295	267	296
rect	267	295	268	296
rect	268	295	269	296
rect	269	295	270	296
rect	270	295	271	296
rect	271	295	272	296
rect	272	295	273	296
rect	273	295	274	296
rect	274	295	275	296
rect	275	295	276	296
rect	276	295	277	296
rect	277	295	278	296
rect	278	295	279	296
rect	279	295	280	296
rect	280	295	281	296
rect	281	295	282	296
rect	282	295	283	296
rect	283	295	284	296
rect	284	295	285	296
rect	285	295	286	296
rect	286	295	287	296
rect	287	295	288	296
rect	288	295	289	296
rect	289	295	290	296
rect	290	295	291	296
rect	291	295	292	296
rect	292	295	293	296
rect	293	295	294	296
rect	294	295	295	296
rect	295	295	296	296
rect	296	295	297	296
rect	297	295	298	296
rect	298	295	299	296
rect	299	295	300	296
rect	301	295	302	296
rect	302	295	303	296
rect	303	295	304	296
rect	304	295	305	296
rect	305	295	306	296
rect	306	295	307	296
rect	307	295	308	296
rect	308	295	309	296
rect	309	295	310	296
rect	310	295	311	296
rect	311	295	312	296
rect	312	295	313	296
rect	313	295	314	296
rect	314	295	315	296
rect	315	295	316	296
rect	317	295	318	296
rect	318	295	319	296
rect	319	295	320	296
rect	320	295	321	296
rect	321	295	322	296
rect	322	295	323	296
rect	323	295	324	296
rect	324	295	325	296
rect	325	295	326	296
rect	326	295	327	296
rect	327	295	328	296
rect	328	295	329	296
rect	329	295	330	296
rect	330	295	331	296
rect	331	295	332	296
rect	332	295	333	296
rect	333	295	334	296
rect	334	295	335	296
rect	335	295	336	296
rect	336	295	337	296
rect	337	295	338	296
rect	338	295	339	296
rect	339	295	340	296
rect	340	295	341	296
rect	341	295	342	296
rect	342	295	343	296
rect	343	295	344	296
rect	344	295	345	296
rect	345	295	346	296
rect	346	295	347	296
rect	347	295	348	296
rect	348	295	349	296
rect	349	295	350	296
rect	350	295	351	296
rect	351	295	352	296
rect	352	295	353	296
rect	353	295	354	296
rect	354	295	355	296
rect	355	295	356	296
rect	356	295	357	296
rect	357	295	358	296
rect	358	295	359	296
rect	359	295	360	296
rect	360	295	361	296
rect	361	295	362	296
rect	362	295	363	296
rect	363	295	364	296
rect	364	295	365	296
rect	365	295	366	296
rect	366	295	367	296
rect	367	295	368	296
rect	368	295	369	296
rect	369	295	370	296
rect	370	295	371	296
rect	371	295	372	296
rect	372	295	373	296
rect	373	295	374	296
rect	374	295	375	296
rect	375	295	376	296
rect	376	295	377	296
rect	377	295	378	296
rect	378	295	379	296
rect	379	295	380	296
rect	380	295	381	296
rect	381	295	382	296
rect	382	295	383	296
rect	383	295	384	296
rect	384	295	385	296
rect	385	295	386	296
rect	386	295	387	296
rect	387	295	388	296
rect	388	295	389	296
rect	389	295	390	296
rect	390	295	391	296
rect	391	295	392	296
rect	392	295	393	296
rect	393	295	394	296
rect	394	295	395	296
rect	396	295	397	296
rect	397	295	398	296
rect	398	295	399	296
rect	399	295	400	296
rect	400	295	401	296
rect	401	295	402	296
rect	0	317	1	318
rect	1	317	2	318
rect	2	317	3	318
rect	3	317	4	318
rect	4	317	5	318
rect	5	317	6	318
rect	7	317	8	318
rect	8	317	9	318
rect	9	317	10	318
rect	10	317	11	318
rect	11	317	12	318
rect	12	317	13	318
rect	13	317	14	318
rect	14	317	15	318
rect	15	317	16	318
rect	16	317	17	318
rect	17	317	18	318
rect	18	317	19	318
rect	19	317	20	318
rect	20	317	21	318
rect	21	317	22	318
rect	23	317	24	318
rect	24	317	25	318
rect	25	317	26	318
rect	26	317	27	318
rect	27	317	28	318
rect	28	317	29	318
rect	30	317	31	318
rect	31	317	32	318
rect	32	317	33	318
rect	33	317	34	318
rect	34	317	35	318
rect	35	317	36	318
rect	37	317	38	318
rect	38	317	39	318
rect	39	317	40	318
rect	40	317	41	318
rect	41	317	42	318
rect	42	317	43	318
rect	43	317	44	318
rect	44	317	45	318
rect	45	317	46	318
rect	46	317	47	318
rect	47	317	48	318
rect	48	317	49	318
rect	49	317	50	318
rect	50	317	51	318
rect	51	317	52	318
rect	52	317	53	318
rect	53	317	54	318
rect	54	317	55	318
rect	55	317	56	318
rect	56	317	57	318
rect	57	317	58	318
rect	58	317	59	318
rect	59	317	60	318
rect	60	317	61	318
rect	61	317	62	318
rect	62	317	63	318
rect	63	317	64	318
rect	64	317	65	318
rect	65	317	66	318
rect	66	317	67	318
rect	67	317	68	318
rect	68	317	69	318
rect	69	317	70	318
rect	70	317	71	318
rect	71	317	72	318
rect	72	317	73	318
rect	73	317	74	318
rect	74	317	75	318
rect	75	317	76	318
rect	76	317	77	318
rect	77	317	78	318
rect	78	317	79	318
rect	79	317	80	318
rect	80	317	81	318
rect	81	317	82	318
rect	82	317	83	318
rect	83	317	84	318
rect	84	317	85	318
rect	85	317	86	318
rect	86	317	87	318
rect	87	317	88	318
rect	88	317	89	318
rect	89	317	90	318
rect	90	317	91	318
rect	91	317	92	318
rect	92	317	93	318
rect	93	317	94	318
rect	94	317	95	318
rect	95	317	96	318
rect	96	317	97	318
rect	97	317	98	318
rect	98	317	99	318
rect	99	317	100	318
rect	100	317	101	318
rect	101	317	102	318
rect	102	317	103	318
rect	103	317	104	318
rect	104	317	105	318
rect	105	317	106	318
rect	106	317	107	318
rect	107	317	108	318
rect	108	317	109	318
rect	109	317	110	318
rect	110	317	111	318
rect	111	317	112	318
rect	112	317	113	318
rect	113	317	114	318
rect	114	317	115	318
rect	115	317	116	318
rect	116	317	117	318
rect	117	317	118	318
rect	118	317	119	318
rect	119	317	120	318
rect	120	317	121	318
rect	121	317	122	318
rect	122	317	123	318
rect	123	317	124	318
rect	124	317	125	318
rect	125	317	126	318
rect	126	317	127	318
rect	127	317	128	318
rect	128	317	129	318
rect	129	317	130	318
rect	130	317	131	318
rect	131	317	132	318
rect	132	317	133	318
rect	133	317	134	318
rect	134	317	135	318
rect	135	317	136	318
rect	136	317	137	318
rect	137	317	138	318
rect	138	317	139	318
rect	139	317	140	318
rect	140	317	141	318
rect	141	317	142	318
rect	142	317	143	318
rect	143	317	144	318
rect	144	317	145	318
rect	145	317	146	318
rect	146	317	147	318
rect	147	317	148	318
rect	148	317	149	318
rect	149	317	150	318
rect	150	317	151	318
rect	151	317	152	318
rect	152	317	153	318
rect	153	317	154	318
rect	154	317	155	318
rect	155	317	156	318
rect	156	317	157	318
rect	157	317	158	318
rect	158	317	159	318
rect	159	317	160	318
rect	160	317	161	318
rect	161	317	162	318
rect	162	317	163	318
rect	163	317	164	318
rect	164	317	165	318
rect	165	317	166	318
rect	166	317	167	318
rect	167	317	168	318
rect	168	317	169	318
rect	169	317	170	318
rect	170	317	171	318
rect	171	317	172	318
rect	172	317	173	318
rect	173	317	174	318
rect	174	317	175	318
rect	175	317	176	318
rect	176	317	177	318
rect	177	317	178	318
rect	178	317	179	318
rect	179	317	180	318
rect	180	317	181	318
rect	181	317	182	318
rect	182	317	183	318
rect	183	317	184	318
rect	184	317	185	318
rect	185	317	186	318
rect	186	317	187	318
rect	187	317	188	318
rect	188	317	189	318
rect	189	317	190	318
rect	190	317	191	318
rect	191	317	192	318
rect	192	317	193	318
rect	193	317	194	318
rect	194	317	195	318
rect	195	317	196	318
rect	196	317	197	318
rect	197	317	198	318
rect	198	317	199	318
rect	199	317	200	318
rect	200	317	201	318
rect	201	317	202	318
rect	202	317	203	318
rect	203	317	204	318
rect	204	317	205	318
rect	205	317	206	318
rect	206	317	207	318
rect	207	317	208	318
rect	208	317	209	318
rect	209	317	210	318
rect	210	317	211	318
rect	211	317	212	318
rect	212	317	213	318
rect	213	317	214	318
rect	214	317	215	318
rect	215	317	216	318
rect	216	317	217	318
rect	217	317	218	318
rect	218	317	219	318
rect	219	317	220	318
rect	220	317	221	318
rect	221	317	222	318
rect	222	317	223	318
rect	223	317	224	318
rect	224	317	225	318
rect	225	317	226	318
rect	226	317	227	318
rect	227	317	228	318
rect	228	317	229	318
rect	229	317	230	318
rect	230	317	231	318
rect	231	317	232	318
rect	232	317	233	318
rect	233	317	234	318
rect	234	317	235	318
rect	235	317	236	318
rect	236	317	237	318
rect	237	317	238	318
rect	238	317	239	318
rect	239	317	240	318
rect	240	317	241	318
rect	241	317	242	318
rect	242	317	243	318
rect	243	317	244	318
rect	244	317	245	318
rect	245	317	246	318
rect	246	317	247	318
rect	247	317	248	318
rect	248	317	249	318
rect	249	317	250	318
rect	250	317	251	318
rect	251	317	252	318
rect	252	317	253	318
rect	253	317	254	318
rect	254	317	255	318
rect	255	317	256	318
rect	256	317	257	318
rect	257	317	258	318
rect	258	317	259	318
rect	259	317	260	318
rect	260	317	261	318
rect	261	317	262	318
rect	262	317	263	318
rect	263	317	264	318
rect	264	317	265	318
rect	265	317	266	318
rect	266	317	267	318
rect	267	317	268	318
rect	268	317	269	318
rect	269	317	270	318
rect	270	317	271	318
rect	271	317	272	318
rect	272	317	273	318
rect	273	317	274	318
rect	274	317	275	318
rect	275	317	276	318
rect	276	317	277	318
rect	277	317	278	318
rect	278	317	279	318
rect	279	317	280	318
rect	280	317	281	318
rect	281	317	282	318
rect	282	317	283	318
rect	283	317	284	318
rect	284	317	285	318
rect	285	317	286	318
rect	286	317	287	318
rect	287	317	288	318
rect	288	317	289	318
rect	289	317	290	318
rect	290	317	291	318
rect	291	317	292	318
rect	292	317	293	318
rect	293	317	294	318
rect	294	317	295	318
rect	295	317	296	318
rect	296	317	297	318
rect	297	317	298	318
rect	298	317	299	318
rect	299	317	300	318
rect	300	317	301	318
rect	302	317	303	318
rect	303	317	304	318
rect	304	317	305	318
rect	305	317	306	318
rect	306	317	307	318
rect	307	317	308	318
rect	309	317	310	318
rect	310	317	311	318
rect	311	317	312	318
rect	312	317	313	318
rect	313	317	314	318
rect	314	317	315	318
rect	316	317	317	318
rect	317	317	318	318
rect	318	317	319	318
rect	319	317	320	318
rect	320	317	321	318
rect	321	317	322	318
rect	322	317	323	318
rect	323	317	324	318
rect	324	317	325	318
rect	325	317	326	318
rect	326	317	327	318
rect	327	317	328	318
rect	328	317	329	318
rect	329	317	330	318
rect	330	317	331	318
rect	331	317	332	318
rect	332	317	333	318
rect	333	317	334	318
rect	334	317	335	318
rect	335	317	336	318
rect	336	317	337	318
rect	337	317	338	318
rect	338	317	339	318
rect	339	317	340	318
rect	340	317	341	318
rect	341	317	342	318
rect	342	317	343	318
rect	344	317	345	318
rect	345	317	346	318
rect	346	317	347	318
rect	347	317	348	318
rect	348	317	349	318
rect	349	317	350	318
rect	351	317	352	318
rect	352	317	353	318
rect	353	317	354	318
rect	354	317	355	318
rect	355	317	356	318
rect	356	317	357	318
rect	357	317	358	318
rect	358	317	359	318
rect	359	317	360	318
rect	360	317	361	318
rect	361	317	362	318
rect	362	317	363	318
rect	363	317	364	318
rect	364	317	365	318
rect	365	317	366	318
rect	366	317	367	318
rect	367	317	368	318
rect	368	317	369	318
rect	369	317	370	318
rect	370	317	371	318
rect	371	317	372	318
rect	372	317	373	318
rect	373	317	374	318
rect	374	317	375	318
rect	375	317	376	318
rect	376	317	377	318
rect	377	317	378	318
rect	378	317	379	318
rect	379	317	380	318
rect	380	317	381	318
rect	381	317	382	318
rect	382	317	383	318
rect	383	317	384	318
rect	384	317	385	318
rect	385	317	386	318
rect	386	317	387	318
rect	387	317	388	318
rect	388	317	389	318
rect	389	317	390	318
rect	390	317	391	318
rect	391	317	392	318
rect	392	317	393	318
rect	393	317	394	318
rect	394	317	395	318
rect	395	317	396	318
rect	396	317	397	318
rect	397	317	398	318
rect	398	317	399	318
rect	399	317	400	318
rect	400	317	401	318
rect	401	317	402	318
rect	403	317	404	318
rect	404	317	405	318
rect	405	317	406	318
rect	406	317	407	318
rect	407	317	408	318
rect	408	317	409	318
rect	409	317	410	318
rect	410	317	411	318
rect	411	317	412	318
rect	412	317	413	318
rect	413	317	414	318
rect	414	317	415	318
rect	415	317	416	318
rect	416	317	417	318
rect	417	317	418	318
rect	418	317	419	318
rect	419	317	420	318
rect	420	317	421	318
rect	0	318	1	319
rect	1	318	2	319
rect	2	318	3	319
rect	3	318	4	319
rect	4	318	5	319
rect	5	318	6	319
rect	7	318	8	319
rect	8	318	9	319
rect	9	318	10	319
rect	10	318	11	319
rect	11	318	12	319
rect	12	318	13	319
rect	13	318	14	319
rect	14	318	15	319
rect	15	318	16	319
rect	16	318	17	319
rect	17	318	18	319
rect	18	318	19	319
rect	19	318	20	319
rect	20	318	21	319
rect	21	318	22	319
rect	23	318	24	319
rect	24	318	25	319
rect	25	318	26	319
rect	26	318	27	319
rect	27	318	28	319
rect	28	318	29	319
rect	30	318	31	319
rect	31	318	32	319
rect	32	318	33	319
rect	33	318	34	319
rect	34	318	35	319
rect	35	318	36	319
rect	37	318	38	319
rect	38	318	39	319
rect	39	318	40	319
rect	40	318	41	319
rect	41	318	42	319
rect	42	318	43	319
rect	43	318	44	319
rect	44	318	45	319
rect	45	318	46	319
rect	46	318	47	319
rect	47	318	48	319
rect	48	318	49	319
rect	49	318	50	319
rect	50	318	51	319
rect	51	318	52	319
rect	52	318	53	319
rect	53	318	54	319
rect	54	318	55	319
rect	55	318	56	319
rect	56	318	57	319
rect	57	318	58	319
rect	58	318	59	319
rect	59	318	60	319
rect	60	318	61	319
rect	61	318	62	319
rect	62	318	63	319
rect	63	318	64	319
rect	64	318	65	319
rect	65	318	66	319
rect	66	318	67	319
rect	67	318	68	319
rect	68	318	69	319
rect	69	318	70	319
rect	70	318	71	319
rect	71	318	72	319
rect	72	318	73	319
rect	73	318	74	319
rect	74	318	75	319
rect	75	318	76	319
rect	76	318	77	319
rect	77	318	78	319
rect	78	318	79	319
rect	79	318	80	319
rect	80	318	81	319
rect	81	318	82	319
rect	82	318	83	319
rect	83	318	84	319
rect	84	318	85	319
rect	85	318	86	319
rect	86	318	87	319
rect	87	318	88	319
rect	88	318	89	319
rect	89	318	90	319
rect	90	318	91	319
rect	91	318	92	319
rect	92	318	93	319
rect	93	318	94	319
rect	94	318	95	319
rect	95	318	96	319
rect	96	318	97	319
rect	97	318	98	319
rect	98	318	99	319
rect	99	318	100	319
rect	100	318	101	319
rect	101	318	102	319
rect	102	318	103	319
rect	103	318	104	319
rect	104	318	105	319
rect	105	318	106	319
rect	106	318	107	319
rect	107	318	108	319
rect	108	318	109	319
rect	109	318	110	319
rect	110	318	111	319
rect	111	318	112	319
rect	112	318	113	319
rect	113	318	114	319
rect	114	318	115	319
rect	115	318	116	319
rect	116	318	117	319
rect	117	318	118	319
rect	118	318	119	319
rect	119	318	120	319
rect	120	318	121	319
rect	121	318	122	319
rect	122	318	123	319
rect	123	318	124	319
rect	124	318	125	319
rect	125	318	126	319
rect	126	318	127	319
rect	127	318	128	319
rect	128	318	129	319
rect	129	318	130	319
rect	130	318	131	319
rect	131	318	132	319
rect	132	318	133	319
rect	133	318	134	319
rect	134	318	135	319
rect	135	318	136	319
rect	136	318	137	319
rect	137	318	138	319
rect	138	318	139	319
rect	139	318	140	319
rect	140	318	141	319
rect	141	318	142	319
rect	142	318	143	319
rect	143	318	144	319
rect	144	318	145	319
rect	145	318	146	319
rect	146	318	147	319
rect	147	318	148	319
rect	148	318	149	319
rect	149	318	150	319
rect	150	318	151	319
rect	151	318	152	319
rect	152	318	153	319
rect	153	318	154	319
rect	154	318	155	319
rect	155	318	156	319
rect	156	318	157	319
rect	157	318	158	319
rect	158	318	159	319
rect	159	318	160	319
rect	160	318	161	319
rect	161	318	162	319
rect	162	318	163	319
rect	163	318	164	319
rect	164	318	165	319
rect	165	318	166	319
rect	166	318	167	319
rect	167	318	168	319
rect	168	318	169	319
rect	169	318	170	319
rect	170	318	171	319
rect	171	318	172	319
rect	172	318	173	319
rect	173	318	174	319
rect	174	318	175	319
rect	175	318	176	319
rect	176	318	177	319
rect	177	318	178	319
rect	178	318	179	319
rect	179	318	180	319
rect	180	318	181	319
rect	181	318	182	319
rect	182	318	183	319
rect	183	318	184	319
rect	184	318	185	319
rect	185	318	186	319
rect	186	318	187	319
rect	187	318	188	319
rect	188	318	189	319
rect	189	318	190	319
rect	190	318	191	319
rect	191	318	192	319
rect	192	318	193	319
rect	193	318	194	319
rect	194	318	195	319
rect	195	318	196	319
rect	196	318	197	319
rect	197	318	198	319
rect	198	318	199	319
rect	199	318	200	319
rect	200	318	201	319
rect	201	318	202	319
rect	202	318	203	319
rect	203	318	204	319
rect	204	318	205	319
rect	205	318	206	319
rect	206	318	207	319
rect	207	318	208	319
rect	208	318	209	319
rect	209	318	210	319
rect	210	318	211	319
rect	211	318	212	319
rect	212	318	213	319
rect	213	318	214	319
rect	214	318	215	319
rect	215	318	216	319
rect	216	318	217	319
rect	217	318	218	319
rect	218	318	219	319
rect	219	318	220	319
rect	220	318	221	319
rect	221	318	222	319
rect	222	318	223	319
rect	223	318	224	319
rect	224	318	225	319
rect	225	318	226	319
rect	226	318	227	319
rect	227	318	228	319
rect	228	318	229	319
rect	229	318	230	319
rect	230	318	231	319
rect	231	318	232	319
rect	232	318	233	319
rect	233	318	234	319
rect	234	318	235	319
rect	235	318	236	319
rect	236	318	237	319
rect	237	318	238	319
rect	238	318	239	319
rect	239	318	240	319
rect	240	318	241	319
rect	241	318	242	319
rect	242	318	243	319
rect	243	318	244	319
rect	244	318	245	319
rect	245	318	246	319
rect	246	318	247	319
rect	247	318	248	319
rect	248	318	249	319
rect	249	318	250	319
rect	250	318	251	319
rect	251	318	252	319
rect	252	318	253	319
rect	253	318	254	319
rect	254	318	255	319
rect	255	318	256	319
rect	256	318	257	319
rect	257	318	258	319
rect	258	318	259	319
rect	259	318	260	319
rect	260	318	261	319
rect	261	318	262	319
rect	262	318	263	319
rect	263	318	264	319
rect	264	318	265	319
rect	265	318	266	319
rect	266	318	267	319
rect	267	318	268	319
rect	268	318	269	319
rect	269	318	270	319
rect	270	318	271	319
rect	271	318	272	319
rect	272	318	273	319
rect	273	318	274	319
rect	274	318	275	319
rect	275	318	276	319
rect	276	318	277	319
rect	277	318	278	319
rect	278	318	279	319
rect	279	318	280	319
rect	280	318	281	319
rect	281	318	282	319
rect	282	318	283	319
rect	283	318	284	319
rect	284	318	285	319
rect	285	318	286	319
rect	286	318	287	319
rect	287	318	288	319
rect	288	318	289	319
rect	289	318	290	319
rect	290	318	291	319
rect	291	318	292	319
rect	292	318	293	319
rect	293	318	294	319
rect	294	318	295	319
rect	295	318	296	319
rect	296	318	297	319
rect	297	318	298	319
rect	298	318	299	319
rect	299	318	300	319
rect	300	318	301	319
rect	302	318	303	319
rect	303	318	304	319
rect	304	318	305	319
rect	305	318	306	319
rect	306	318	307	319
rect	307	318	308	319
rect	309	318	310	319
rect	310	318	311	319
rect	311	318	312	319
rect	312	318	313	319
rect	313	318	314	319
rect	314	318	315	319
rect	316	318	317	319
rect	317	318	318	319
rect	318	318	319	319
rect	319	318	320	319
rect	320	318	321	319
rect	321	318	322	319
rect	322	318	323	319
rect	323	318	324	319
rect	324	318	325	319
rect	325	318	326	319
rect	326	318	327	319
rect	327	318	328	319
rect	328	318	329	319
rect	329	318	330	319
rect	330	318	331	319
rect	331	318	332	319
rect	332	318	333	319
rect	333	318	334	319
rect	334	318	335	319
rect	335	318	336	319
rect	336	318	337	319
rect	337	318	338	319
rect	338	318	339	319
rect	339	318	340	319
rect	340	318	341	319
rect	341	318	342	319
rect	342	318	343	319
rect	344	318	345	319
rect	345	318	346	319
rect	346	318	347	319
rect	347	318	348	319
rect	348	318	349	319
rect	349	318	350	319
rect	351	318	352	319
rect	352	318	353	319
rect	353	318	354	319
rect	354	318	355	319
rect	355	318	356	319
rect	356	318	357	319
rect	357	318	358	319
rect	358	318	359	319
rect	359	318	360	319
rect	360	318	361	319
rect	361	318	362	319
rect	362	318	363	319
rect	363	318	364	319
rect	364	318	365	319
rect	365	318	366	319
rect	366	318	367	319
rect	367	318	368	319
rect	368	318	369	319
rect	369	318	370	319
rect	370	318	371	319
rect	371	318	372	319
rect	372	318	373	319
rect	373	318	374	319
rect	374	318	375	319
rect	375	318	376	319
rect	376	318	377	319
rect	377	318	378	319
rect	378	318	379	319
rect	379	318	380	319
rect	380	318	381	319
rect	381	318	382	319
rect	382	318	383	319
rect	383	318	384	319
rect	384	318	385	319
rect	385	318	386	319
rect	386	318	387	319
rect	387	318	388	319
rect	388	318	389	319
rect	389	318	390	319
rect	390	318	391	319
rect	391	318	392	319
rect	392	318	393	319
rect	393	318	394	319
rect	394	318	395	319
rect	395	318	396	319
rect	396	318	397	319
rect	397	318	398	319
rect	398	318	399	319
rect	399	318	400	319
rect	400	318	401	319
rect	401	318	402	319
rect	403	318	404	319
rect	404	318	405	319
rect	405	318	406	319
rect	406	318	407	319
rect	407	318	408	319
rect	408	318	409	319
rect	409	318	410	319
rect	410	318	411	319
rect	411	318	412	319
rect	412	318	413	319
rect	413	318	414	319
rect	414	318	415	319
rect	415	318	416	319
rect	416	318	417	319
rect	417	318	418	319
rect	418	318	419	319
rect	419	318	420	319
rect	420	318	421	319
rect	0	319	1	320
rect	1	319	2	320
rect	2	319	3	320
rect	3	319	4	320
rect	4	319	5	320
rect	5	319	6	320
rect	7	319	8	320
rect	8	319	9	320
rect	9	319	10	320
rect	10	319	11	320
rect	11	319	12	320
rect	12	319	13	320
rect	13	319	14	320
rect	14	319	15	320
rect	15	319	16	320
rect	16	319	17	320
rect	17	319	18	320
rect	18	319	19	320
rect	19	319	20	320
rect	20	319	21	320
rect	21	319	22	320
rect	23	319	24	320
rect	24	319	25	320
rect	25	319	26	320
rect	26	319	27	320
rect	27	319	28	320
rect	28	319	29	320
rect	30	319	31	320
rect	31	319	32	320
rect	32	319	33	320
rect	33	319	34	320
rect	34	319	35	320
rect	35	319	36	320
rect	37	319	38	320
rect	38	319	39	320
rect	39	319	40	320
rect	40	319	41	320
rect	41	319	42	320
rect	42	319	43	320
rect	43	319	44	320
rect	44	319	45	320
rect	45	319	46	320
rect	46	319	47	320
rect	47	319	48	320
rect	48	319	49	320
rect	49	319	50	320
rect	50	319	51	320
rect	51	319	52	320
rect	52	319	53	320
rect	53	319	54	320
rect	54	319	55	320
rect	55	319	56	320
rect	56	319	57	320
rect	57	319	58	320
rect	58	319	59	320
rect	59	319	60	320
rect	60	319	61	320
rect	61	319	62	320
rect	62	319	63	320
rect	63	319	64	320
rect	64	319	65	320
rect	65	319	66	320
rect	66	319	67	320
rect	67	319	68	320
rect	68	319	69	320
rect	69	319	70	320
rect	70	319	71	320
rect	71	319	72	320
rect	72	319	73	320
rect	73	319	74	320
rect	74	319	75	320
rect	75	319	76	320
rect	76	319	77	320
rect	77	319	78	320
rect	78	319	79	320
rect	79	319	80	320
rect	80	319	81	320
rect	81	319	82	320
rect	82	319	83	320
rect	83	319	84	320
rect	84	319	85	320
rect	85	319	86	320
rect	86	319	87	320
rect	87	319	88	320
rect	88	319	89	320
rect	89	319	90	320
rect	90	319	91	320
rect	91	319	92	320
rect	92	319	93	320
rect	93	319	94	320
rect	94	319	95	320
rect	95	319	96	320
rect	96	319	97	320
rect	97	319	98	320
rect	98	319	99	320
rect	99	319	100	320
rect	100	319	101	320
rect	101	319	102	320
rect	102	319	103	320
rect	103	319	104	320
rect	104	319	105	320
rect	105	319	106	320
rect	106	319	107	320
rect	107	319	108	320
rect	108	319	109	320
rect	109	319	110	320
rect	110	319	111	320
rect	111	319	112	320
rect	112	319	113	320
rect	113	319	114	320
rect	114	319	115	320
rect	115	319	116	320
rect	116	319	117	320
rect	117	319	118	320
rect	118	319	119	320
rect	119	319	120	320
rect	120	319	121	320
rect	121	319	122	320
rect	122	319	123	320
rect	123	319	124	320
rect	124	319	125	320
rect	125	319	126	320
rect	126	319	127	320
rect	127	319	128	320
rect	128	319	129	320
rect	129	319	130	320
rect	130	319	131	320
rect	131	319	132	320
rect	132	319	133	320
rect	133	319	134	320
rect	134	319	135	320
rect	135	319	136	320
rect	136	319	137	320
rect	137	319	138	320
rect	138	319	139	320
rect	139	319	140	320
rect	140	319	141	320
rect	141	319	142	320
rect	142	319	143	320
rect	143	319	144	320
rect	144	319	145	320
rect	145	319	146	320
rect	146	319	147	320
rect	147	319	148	320
rect	148	319	149	320
rect	149	319	150	320
rect	150	319	151	320
rect	151	319	152	320
rect	152	319	153	320
rect	153	319	154	320
rect	154	319	155	320
rect	155	319	156	320
rect	156	319	157	320
rect	157	319	158	320
rect	158	319	159	320
rect	159	319	160	320
rect	160	319	161	320
rect	161	319	162	320
rect	162	319	163	320
rect	163	319	164	320
rect	164	319	165	320
rect	165	319	166	320
rect	166	319	167	320
rect	167	319	168	320
rect	168	319	169	320
rect	169	319	170	320
rect	170	319	171	320
rect	171	319	172	320
rect	172	319	173	320
rect	173	319	174	320
rect	174	319	175	320
rect	175	319	176	320
rect	176	319	177	320
rect	177	319	178	320
rect	178	319	179	320
rect	179	319	180	320
rect	180	319	181	320
rect	181	319	182	320
rect	182	319	183	320
rect	183	319	184	320
rect	184	319	185	320
rect	185	319	186	320
rect	186	319	187	320
rect	187	319	188	320
rect	188	319	189	320
rect	189	319	190	320
rect	190	319	191	320
rect	191	319	192	320
rect	192	319	193	320
rect	193	319	194	320
rect	194	319	195	320
rect	195	319	196	320
rect	196	319	197	320
rect	197	319	198	320
rect	198	319	199	320
rect	199	319	200	320
rect	200	319	201	320
rect	201	319	202	320
rect	202	319	203	320
rect	203	319	204	320
rect	204	319	205	320
rect	205	319	206	320
rect	206	319	207	320
rect	207	319	208	320
rect	208	319	209	320
rect	209	319	210	320
rect	210	319	211	320
rect	211	319	212	320
rect	212	319	213	320
rect	213	319	214	320
rect	214	319	215	320
rect	215	319	216	320
rect	216	319	217	320
rect	217	319	218	320
rect	218	319	219	320
rect	219	319	220	320
rect	220	319	221	320
rect	221	319	222	320
rect	222	319	223	320
rect	223	319	224	320
rect	224	319	225	320
rect	225	319	226	320
rect	226	319	227	320
rect	227	319	228	320
rect	228	319	229	320
rect	229	319	230	320
rect	230	319	231	320
rect	231	319	232	320
rect	232	319	233	320
rect	233	319	234	320
rect	234	319	235	320
rect	235	319	236	320
rect	236	319	237	320
rect	237	319	238	320
rect	238	319	239	320
rect	239	319	240	320
rect	240	319	241	320
rect	241	319	242	320
rect	242	319	243	320
rect	243	319	244	320
rect	244	319	245	320
rect	245	319	246	320
rect	246	319	247	320
rect	247	319	248	320
rect	248	319	249	320
rect	249	319	250	320
rect	250	319	251	320
rect	251	319	252	320
rect	252	319	253	320
rect	253	319	254	320
rect	254	319	255	320
rect	255	319	256	320
rect	256	319	257	320
rect	257	319	258	320
rect	258	319	259	320
rect	259	319	260	320
rect	260	319	261	320
rect	261	319	262	320
rect	262	319	263	320
rect	263	319	264	320
rect	264	319	265	320
rect	265	319	266	320
rect	266	319	267	320
rect	267	319	268	320
rect	268	319	269	320
rect	269	319	270	320
rect	270	319	271	320
rect	271	319	272	320
rect	272	319	273	320
rect	273	319	274	320
rect	274	319	275	320
rect	275	319	276	320
rect	276	319	277	320
rect	277	319	278	320
rect	278	319	279	320
rect	279	319	280	320
rect	280	319	281	320
rect	281	319	282	320
rect	282	319	283	320
rect	283	319	284	320
rect	284	319	285	320
rect	285	319	286	320
rect	286	319	287	320
rect	287	319	288	320
rect	288	319	289	320
rect	289	319	290	320
rect	290	319	291	320
rect	291	319	292	320
rect	292	319	293	320
rect	293	319	294	320
rect	294	319	295	320
rect	295	319	296	320
rect	296	319	297	320
rect	297	319	298	320
rect	298	319	299	320
rect	299	319	300	320
rect	300	319	301	320
rect	302	319	303	320
rect	303	319	304	320
rect	304	319	305	320
rect	305	319	306	320
rect	306	319	307	320
rect	307	319	308	320
rect	309	319	310	320
rect	310	319	311	320
rect	311	319	312	320
rect	312	319	313	320
rect	313	319	314	320
rect	314	319	315	320
rect	316	319	317	320
rect	317	319	318	320
rect	318	319	319	320
rect	319	319	320	320
rect	320	319	321	320
rect	321	319	322	320
rect	322	319	323	320
rect	323	319	324	320
rect	324	319	325	320
rect	325	319	326	320
rect	326	319	327	320
rect	327	319	328	320
rect	328	319	329	320
rect	329	319	330	320
rect	330	319	331	320
rect	331	319	332	320
rect	332	319	333	320
rect	333	319	334	320
rect	334	319	335	320
rect	335	319	336	320
rect	336	319	337	320
rect	337	319	338	320
rect	338	319	339	320
rect	339	319	340	320
rect	340	319	341	320
rect	341	319	342	320
rect	342	319	343	320
rect	344	319	345	320
rect	345	319	346	320
rect	346	319	347	320
rect	347	319	348	320
rect	348	319	349	320
rect	349	319	350	320
rect	351	319	352	320
rect	352	319	353	320
rect	353	319	354	320
rect	354	319	355	320
rect	355	319	356	320
rect	356	319	357	320
rect	357	319	358	320
rect	358	319	359	320
rect	359	319	360	320
rect	360	319	361	320
rect	361	319	362	320
rect	362	319	363	320
rect	363	319	364	320
rect	364	319	365	320
rect	365	319	366	320
rect	366	319	367	320
rect	367	319	368	320
rect	368	319	369	320
rect	369	319	370	320
rect	370	319	371	320
rect	371	319	372	320
rect	372	319	373	320
rect	373	319	374	320
rect	374	319	375	320
rect	375	319	376	320
rect	376	319	377	320
rect	377	319	378	320
rect	378	319	379	320
rect	379	319	380	320
rect	380	319	381	320
rect	381	319	382	320
rect	382	319	383	320
rect	383	319	384	320
rect	384	319	385	320
rect	385	319	386	320
rect	386	319	387	320
rect	387	319	388	320
rect	388	319	389	320
rect	389	319	390	320
rect	390	319	391	320
rect	391	319	392	320
rect	392	319	393	320
rect	393	319	394	320
rect	394	319	395	320
rect	395	319	396	320
rect	396	319	397	320
rect	397	319	398	320
rect	398	319	399	320
rect	399	319	400	320
rect	400	319	401	320
rect	401	319	402	320
rect	403	319	404	320
rect	404	319	405	320
rect	405	319	406	320
rect	406	319	407	320
rect	407	319	408	320
rect	408	319	409	320
rect	409	319	410	320
rect	410	319	411	320
rect	411	319	412	320
rect	412	319	413	320
rect	413	319	414	320
rect	414	319	415	320
rect	415	319	416	320
rect	416	319	417	320
rect	417	319	418	320
rect	418	319	419	320
rect	419	319	420	320
rect	420	319	421	320
rect	0	320	1	321
rect	1	320	2	321
rect	2	320	3	321
rect	3	320	4	321
rect	4	320	5	321
rect	5	320	6	321
rect	7	320	8	321
rect	8	320	9	321
rect	9	320	10	321
rect	10	320	11	321
rect	11	320	12	321
rect	12	320	13	321
rect	13	320	14	321
rect	14	320	15	321
rect	15	320	16	321
rect	16	320	17	321
rect	17	320	18	321
rect	18	320	19	321
rect	19	320	20	321
rect	20	320	21	321
rect	21	320	22	321
rect	23	320	24	321
rect	24	320	25	321
rect	25	320	26	321
rect	26	320	27	321
rect	27	320	28	321
rect	28	320	29	321
rect	30	320	31	321
rect	31	320	32	321
rect	32	320	33	321
rect	33	320	34	321
rect	34	320	35	321
rect	35	320	36	321
rect	37	320	38	321
rect	38	320	39	321
rect	39	320	40	321
rect	40	320	41	321
rect	41	320	42	321
rect	42	320	43	321
rect	43	320	44	321
rect	44	320	45	321
rect	45	320	46	321
rect	46	320	47	321
rect	47	320	48	321
rect	48	320	49	321
rect	49	320	50	321
rect	50	320	51	321
rect	51	320	52	321
rect	52	320	53	321
rect	53	320	54	321
rect	54	320	55	321
rect	55	320	56	321
rect	56	320	57	321
rect	57	320	58	321
rect	58	320	59	321
rect	59	320	60	321
rect	60	320	61	321
rect	61	320	62	321
rect	62	320	63	321
rect	63	320	64	321
rect	64	320	65	321
rect	65	320	66	321
rect	66	320	67	321
rect	67	320	68	321
rect	68	320	69	321
rect	69	320	70	321
rect	70	320	71	321
rect	71	320	72	321
rect	72	320	73	321
rect	73	320	74	321
rect	74	320	75	321
rect	75	320	76	321
rect	76	320	77	321
rect	77	320	78	321
rect	78	320	79	321
rect	79	320	80	321
rect	80	320	81	321
rect	81	320	82	321
rect	82	320	83	321
rect	83	320	84	321
rect	84	320	85	321
rect	85	320	86	321
rect	86	320	87	321
rect	87	320	88	321
rect	88	320	89	321
rect	89	320	90	321
rect	90	320	91	321
rect	91	320	92	321
rect	92	320	93	321
rect	93	320	94	321
rect	94	320	95	321
rect	95	320	96	321
rect	96	320	97	321
rect	97	320	98	321
rect	98	320	99	321
rect	99	320	100	321
rect	100	320	101	321
rect	101	320	102	321
rect	102	320	103	321
rect	103	320	104	321
rect	104	320	105	321
rect	105	320	106	321
rect	106	320	107	321
rect	107	320	108	321
rect	108	320	109	321
rect	109	320	110	321
rect	110	320	111	321
rect	111	320	112	321
rect	112	320	113	321
rect	113	320	114	321
rect	114	320	115	321
rect	115	320	116	321
rect	116	320	117	321
rect	117	320	118	321
rect	118	320	119	321
rect	119	320	120	321
rect	120	320	121	321
rect	121	320	122	321
rect	122	320	123	321
rect	123	320	124	321
rect	124	320	125	321
rect	125	320	126	321
rect	126	320	127	321
rect	127	320	128	321
rect	128	320	129	321
rect	129	320	130	321
rect	130	320	131	321
rect	131	320	132	321
rect	132	320	133	321
rect	133	320	134	321
rect	134	320	135	321
rect	135	320	136	321
rect	136	320	137	321
rect	137	320	138	321
rect	138	320	139	321
rect	139	320	140	321
rect	140	320	141	321
rect	141	320	142	321
rect	142	320	143	321
rect	143	320	144	321
rect	144	320	145	321
rect	145	320	146	321
rect	146	320	147	321
rect	147	320	148	321
rect	148	320	149	321
rect	149	320	150	321
rect	150	320	151	321
rect	151	320	152	321
rect	152	320	153	321
rect	153	320	154	321
rect	154	320	155	321
rect	155	320	156	321
rect	156	320	157	321
rect	157	320	158	321
rect	158	320	159	321
rect	159	320	160	321
rect	160	320	161	321
rect	161	320	162	321
rect	162	320	163	321
rect	163	320	164	321
rect	164	320	165	321
rect	165	320	166	321
rect	166	320	167	321
rect	167	320	168	321
rect	168	320	169	321
rect	169	320	170	321
rect	170	320	171	321
rect	171	320	172	321
rect	172	320	173	321
rect	173	320	174	321
rect	174	320	175	321
rect	175	320	176	321
rect	176	320	177	321
rect	177	320	178	321
rect	178	320	179	321
rect	179	320	180	321
rect	180	320	181	321
rect	181	320	182	321
rect	182	320	183	321
rect	183	320	184	321
rect	184	320	185	321
rect	185	320	186	321
rect	186	320	187	321
rect	187	320	188	321
rect	188	320	189	321
rect	189	320	190	321
rect	190	320	191	321
rect	191	320	192	321
rect	192	320	193	321
rect	193	320	194	321
rect	194	320	195	321
rect	195	320	196	321
rect	196	320	197	321
rect	197	320	198	321
rect	198	320	199	321
rect	199	320	200	321
rect	200	320	201	321
rect	201	320	202	321
rect	202	320	203	321
rect	203	320	204	321
rect	204	320	205	321
rect	205	320	206	321
rect	206	320	207	321
rect	207	320	208	321
rect	208	320	209	321
rect	209	320	210	321
rect	210	320	211	321
rect	211	320	212	321
rect	212	320	213	321
rect	213	320	214	321
rect	214	320	215	321
rect	215	320	216	321
rect	216	320	217	321
rect	217	320	218	321
rect	218	320	219	321
rect	219	320	220	321
rect	220	320	221	321
rect	221	320	222	321
rect	222	320	223	321
rect	223	320	224	321
rect	224	320	225	321
rect	225	320	226	321
rect	226	320	227	321
rect	227	320	228	321
rect	228	320	229	321
rect	229	320	230	321
rect	230	320	231	321
rect	231	320	232	321
rect	232	320	233	321
rect	233	320	234	321
rect	234	320	235	321
rect	235	320	236	321
rect	236	320	237	321
rect	237	320	238	321
rect	238	320	239	321
rect	239	320	240	321
rect	240	320	241	321
rect	241	320	242	321
rect	242	320	243	321
rect	243	320	244	321
rect	244	320	245	321
rect	245	320	246	321
rect	246	320	247	321
rect	247	320	248	321
rect	248	320	249	321
rect	249	320	250	321
rect	250	320	251	321
rect	251	320	252	321
rect	252	320	253	321
rect	253	320	254	321
rect	254	320	255	321
rect	255	320	256	321
rect	256	320	257	321
rect	257	320	258	321
rect	258	320	259	321
rect	259	320	260	321
rect	260	320	261	321
rect	261	320	262	321
rect	262	320	263	321
rect	263	320	264	321
rect	264	320	265	321
rect	265	320	266	321
rect	266	320	267	321
rect	267	320	268	321
rect	268	320	269	321
rect	269	320	270	321
rect	270	320	271	321
rect	271	320	272	321
rect	272	320	273	321
rect	273	320	274	321
rect	274	320	275	321
rect	275	320	276	321
rect	276	320	277	321
rect	277	320	278	321
rect	278	320	279	321
rect	279	320	280	321
rect	280	320	281	321
rect	281	320	282	321
rect	282	320	283	321
rect	283	320	284	321
rect	284	320	285	321
rect	285	320	286	321
rect	286	320	287	321
rect	287	320	288	321
rect	288	320	289	321
rect	289	320	290	321
rect	290	320	291	321
rect	291	320	292	321
rect	292	320	293	321
rect	293	320	294	321
rect	294	320	295	321
rect	295	320	296	321
rect	296	320	297	321
rect	297	320	298	321
rect	298	320	299	321
rect	299	320	300	321
rect	300	320	301	321
rect	302	320	303	321
rect	303	320	304	321
rect	304	320	305	321
rect	305	320	306	321
rect	306	320	307	321
rect	307	320	308	321
rect	309	320	310	321
rect	310	320	311	321
rect	311	320	312	321
rect	312	320	313	321
rect	313	320	314	321
rect	314	320	315	321
rect	316	320	317	321
rect	317	320	318	321
rect	318	320	319	321
rect	319	320	320	321
rect	320	320	321	321
rect	321	320	322	321
rect	322	320	323	321
rect	323	320	324	321
rect	324	320	325	321
rect	325	320	326	321
rect	326	320	327	321
rect	327	320	328	321
rect	328	320	329	321
rect	329	320	330	321
rect	330	320	331	321
rect	331	320	332	321
rect	332	320	333	321
rect	333	320	334	321
rect	334	320	335	321
rect	335	320	336	321
rect	336	320	337	321
rect	337	320	338	321
rect	338	320	339	321
rect	339	320	340	321
rect	340	320	341	321
rect	341	320	342	321
rect	342	320	343	321
rect	344	320	345	321
rect	345	320	346	321
rect	346	320	347	321
rect	347	320	348	321
rect	348	320	349	321
rect	349	320	350	321
rect	351	320	352	321
rect	352	320	353	321
rect	353	320	354	321
rect	354	320	355	321
rect	355	320	356	321
rect	356	320	357	321
rect	357	320	358	321
rect	358	320	359	321
rect	359	320	360	321
rect	360	320	361	321
rect	361	320	362	321
rect	362	320	363	321
rect	363	320	364	321
rect	364	320	365	321
rect	365	320	366	321
rect	366	320	367	321
rect	367	320	368	321
rect	368	320	369	321
rect	369	320	370	321
rect	370	320	371	321
rect	371	320	372	321
rect	372	320	373	321
rect	373	320	374	321
rect	374	320	375	321
rect	375	320	376	321
rect	376	320	377	321
rect	377	320	378	321
rect	378	320	379	321
rect	379	320	380	321
rect	380	320	381	321
rect	381	320	382	321
rect	382	320	383	321
rect	383	320	384	321
rect	384	320	385	321
rect	385	320	386	321
rect	386	320	387	321
rect	387	320	388	321
rect	388	320	389	321
rect	389	320	390	321
rect	390	320	391	321
rect	391	320	392	321
rect	392	320	393	321
rect	393	320	394	321
rect	394	320	395	321
rect	395	320	396	321
rect	396	320	397	321
rect	397	320	398	321
rect	398	320	399	321
rect	399	320	400	321
rect	400	320	401	321
rect	401	320	402	321
rect	403	320	404	321
rect	404	320	405	321
rect	405	320	406	321
rect	406	320	407	321
rect	407	320	408	321
rect	408	320	409	321
rect	409	320	410	321
rect	410	320	411	321
rect	411	320	412	321
rect	412	320	413	321
rect	413	320	414	321
rect	414	320	415	321
rect	415	320	416	321
rect	416	320	417	321
rect	417	320	418	321
rect	418	320	419	321
rect	419	320	420	321
rect	420	320	421	321
rect	0	321	1	322
rect	1	321	2	322
rect	2	321	3	322
rect	3	321	4	322
rect	4	321	5	322
rect	5	321	6	322
rect	7	321	8	322
rect	8	321	9	322
rect	9	321	10	322
rect	10	321	11	322
rect	11	321	12	322
rect	12	321	13	322
rect	13	321	14	322
rect	14	321	15	322
rect	15	321	16	322
rect	16	321	17	322
rect	17	321	18	322
rect	18	321	19	322
rect	19	321	20	322
rect	20	321	21	322
rect	21	321	22	322
rect	23	321	24	322
rect	24	321	25	322
rect	25	321	26	322
rect	26	321	27	322
rect	27	321	28	322
rect	28	321	29	322
rect	30	321	31	322
rect	31	321	32	322
rect	32	321	33	322
rect	33	321	34	322
rect	34	321	35	322
rect	35	321	36	322
rect	37	321	38	322
rect	38	321	39	322
rect	39	321	40	322
rect	40	321	41	322
rect	41	321	42	322
rect	42	321	43	322
rect	43	321	44	322
rect	44	321	45	322
rect	45	321	46	322
rect	46	321	47	322
rect	47	321	48	322
rect	48	321	49	322
rect	49	321	50	322
rect	50	321	51	322
rect	51	321	52	322
rect	52	321	53	322
rect	53	321	54	322
rect	54	321	55	322
rect	55	321	56	322
rect	56	321	57	322
rect	57	321	58	322
rect	58	321	59	322
rect	59	321	60	322
rect	60	321	61	322
rect	61	321	62	322
rect	62	321	63	322
rect	63	321	64	322
rect	64	321	65	322
rect	65	321	66	322
rect	66	321	67	322
rect	67	321	68	322
rect	68	321	69	322
rect	69	321	70	322
rect	70	321	71	322
rect	71	321	72	322
rect	72	321	73	322
rect	73	321	74	322
rect	74	321	75	322
rect	75	321	76	322
rect	76	321	77	322
rect	77	321	78	322
rect	78	321	79	322
rect	79	321	80	322
rect	80	321	81	322
rect	81	321	82	322
rect	82	321	83	322
rect	83	321	84	322
rect	84	321	85	322
rect	85	321	86	322
rect	86	321	87	322
rect	87	321	88	322
rect	88	321	89	322
rect	89	321	90	322
rect	90	321	91	322
rect	91	321	92	322
rect	92	321	93	322
rect	93	321	94	322
rect	94	321	95	322
rect	95	321	96	322
rect	96	321	97	322
rect	97	321	98	322
rect	98	321	99	322
rect	99	321	100	322
rect	100	321	101	322
rect	101	321	102	322
rect	102	321	103	322
rect	103	321	104	322
rect	104	321	105	322
rect	105	321	106	322
rect	106	321	107	322
rect	107	321	108	322
rect	108	321	109	322
rect	109	321	110	322
rect	110	321	111	322
rect	111	321	112	322
rect	112	321	113	322
rect	113	321	114	322
rect	114	321	115	322
rect	115	321	116	322
rect	116	321	117	322
rect	117	321	118	322
rect	118	321	119	322
rect	119	321	120	322
rect	120	321	121	322
rect	121	321	122	322
rect	122	321	123	322
rect	123	321	124	322
rect	124	321	125	322
rect	125	321	126	322
rect	126	321	127	322
rect	127	321	128	322
rect	128	321	129	322
rect	129	321	130	322
rect	130	321	131	322
rect	131	321	132	322
rect	132	321	133	322
rect	133	321	134	322
rect	134	321	135	322
rect	135	321	136	322
rect	136	321	137	322
rect	137	321	138	322
rect	138	321	139	322
rect	139	321	140	322
rect	140	321	141	322
rect	141	321	142	322
rect	142	321	143	322
rect	143	321	144	322
rect	144	321	145	322
rect	145	321	146	322
rect	146	321	147	322
rect	147	321	148	322
rect	148	321	149	322
rect	149	321	150	322
rect	150	321	151	322
rect	151	321	152	322
rect	152	321	153	322
rect	153	321	154	322
rect	154	321	155	322
rect	155	321	156	322
rect	156	321	157	322
rect	157	321	158	322
rect	158	321	159	322
rect	159	321	160	322
rect	160	321	161	322
rect	161	321	162	322
rect	162	321	163	322
rect	163	321	164	322
rect	164	321	165	322
rect	165	321	166	322
rect	166	321	167	322
rect	167	321	168	322
rect	168	321	169	322
rect	169	321	170	322
rect	170	321	171	322
rect	171	321	172	322
rect	172	321	173	322
rect	173	321	174	322
rect	174	321	175	322
rect	175	321	176	322
rect	176	321	177	322
rect	177	321	178	322
rect	178	321	179	322
rect	179	321	180	322
rect	180	321	181	322
rect	181	321	182	322
rect	182	321	183	322
rect	183	321	184	322
rect	184	321	185	322
rect	185	321	186	322
rect	186	321	187	322
rect	187	321	188	322
rect	188	321	189	322
rect	189	321	190	322
rect	190	321	191	322
rect	191	321	192	322
rect	192	321	193	322
rect	193	321	194	322
rect	194	321	195	322
rect	195	321	196	322
rect	196	321	197	322
rect	197	321	198	322
rect	198	321	199	322
rect	199	321	200	322
rect	200	321	201	322
rect	201	321	202	322
rect	202	321	203	322
rect	203	321	204	322
rect	204	321	205	322
rect	205	321	206	322
rect	206	321	207	322
rect	207	321	208	322
rect	208	321	209	322
rect	209	321	210	322
rect	210	321	211	322
rect	211	321	212	322
rect	212	321	213	322
rect	213	321	214	322
rect	214	321	215	322
rect	215	321	216	322
rect	216	321	217	322
rect	217	321	218	322
rect	218	321	219	322
rect	219	321	220	322
rect	220	321	221	322
rect	221	321	222	322
rect	222	321	223	322
rect	223	321	224	322
rect	224	321	225	322
rect	225	321	226	322
rect	226	321	227	322
rect	227	321	228	322
rect	228	321	229	322
rect	229	321	230	322
rect	230	321	231	322
rect	231	321	232	322
rect	232	321	233	322
rect	233	321	234	322
rect	234	321	235	322
rect	235	321	236	322
rect	236	321	237	322
rect	237	321	238	322
rect	238	321	239	322
rect	239	321	240	322
rect	240	321	241	322
rect	241	321	242	322
rect	242	321	243	322
rect	243	321	244	322
rect	244	321	245	322
rect	245	321	246	322
rect	246	321	247	322
rect	247	321	248	322
rect	248	321	249	322
rect	249	321	250	322
rect	250	321	251	322
rect	251	321	252	322
rect	252	321	253	322
rect	253	321	254	322
rect	254	321	255	322
rect	255	321	256	322
rect	256	321	257	322
rect	257	321	258	322
rect	258	321	259	322
rect	259	321	260	322
rect	260	321	261	322
rect	261	321	262	322
rect	262	321	263	322
rect	263	321	264	322
rect	264	321	265	322
rect	265	321	266	322
rect	266	321	267	322
rect	267	321	268	322
rect	268	321	269	322
rect	269	321	270	322
rect	270	321	271	322
rect	271	321	272	322
rect	272	321	273	322
rect	273	321	274	322
rect	274	321	275	322
rect	275	321	276	322
rect	276	321	277	322
rect	277	321	278	322
rect	278	321	279	322
rect	279	321	280	322
rect	280	321	281	322
rect	281	321	282	322
rect	282	321	283	322
rect	283	321	284	322
rect	284	321	285	322
rect	285	321	286	322
rect	286	321	287	322
rect	287	321	288	322
rect	288	321	289	322
rect	289	321	290	322
rect	290	321	291	322
rect	291	321	292	322
rect	292	321	293	322
rect	293	321	294	322
rect	294	321	295	322
rect	295	321	296	322
rect	296	321	297	322
rect	297	321	298	322
rect	298	321	299	322
rect	299	321	300	322
rect	300	321	301	322
rect	302	321	303	322
rect	303	321	304	322
rect	304	321	305	322
rect	305	321	306	322
rect	306	321	307	322
rect	307	321	308	322
rect	309	321	310	322
rect	310	321	311	322
rect	311	321	312	322
rect	312	321	313	322
rect	313	321	314	322
rect	314	321	315	322
rect	316	321	317	322
rect	317	321	318	322
rect	318	321	319	322
rect	319	321	320	322
rect	320	321	321	322
rect	321	321	322	322
rect	322	321	323	322
rect	323	321	324	322
rect	324	321	325	322
rect	325	321	326	322
rect	326	321	327	322
rect	327	321	328	322
rect	328	321	329	322
rect	329	321	330	322
rect	330	321	331	322
rect	331	321	332	322
rect	332	321	333	322
rect	333	321	334	322
rect	334	321	335	322
rect	335	321	336	322
rect	336	321	337	322
rect	337	321	338	322
rect	338	321	339	322
rect	339	321	340	322
rect	340	321	341	322
rect	341	321	342	322
rect	342	321	343	322
rect	344	321	345	322
rect	345	321	346	322
rect	346	321	347	322
rect	347	321	348	322
rect	348	321	349	322
rect	349	321	350	322
rect	351	321	352	322
rect	352	321	353	322
rect	353	321	354	322
rect	354	321	355	322
rect	355	321	356	322
rect	356	321	357	322
rect	357	321	358	322
rect	358	321	359	322
rect	359	321	360	322
rect	360	321	361	322
rect	361	321	362	322
rect	362	321	363	322
rect	363	321	364	322
rect	364	321	365	322
rect	365	321	366	322
rect	366	321	367	322
rect	367	321	368	322
rect	368	321	369	322
rect	369	321	370	322
rect	370	321	371	322
rect	371	321	372	322
rect	372	321	373	322
rect	373	321	374	322
rect	374	321	375	322
rect	375	321	376	322
rect	376	321	377	322
rect	377	321	378	322
rect	378	321	379	322
rect	379	321	380	322
rect	380	321	381	322
rect	381	321	382	322
rect	382	321	383	322
rect	383	321	384	322
rect	384	321	385	322
rect	385	321	386	322
rect	386	321	387	322
rect	387	321	388	322
rect	388	321	389	322
rect	389	321	390	322
rect	390	321	391	322
rect	391	321	392	322
rect	392	321	393	322
rect	393	321	394	322
rect	394	321	395	322
rect	395	321	396	322
rect	396	321	397	322
rect	397	321	398	322
rect	398	321	399	322
rect	399	321	400	322
rect	400	321	401	322
rect	401	321	402	322
rect	403	321	404	322
rect	404	321	405	322
rect	405	321	406	322
rect	406	321	407	322
rect	407	321	408	322
rect	408	321	409	322
rect	409	321	410	322
rect	410	321	411	322
rect	411	321	412	322
rect	412	321	413	322
rect	413	321	414	322
rect	414	321	415	322
rect	415	321	416	322
rect	416	321	417	322
rect	417	321	418	322
rect	418	321	419	322
rect	419	321	420	322
rect	420	321	421	322
rect	0	322	1	323
rect	1	322	2	323
rect	2	322	3	323
rect	3	322	4	323
rect	4	322	5	323
rect	5	322	6	323
rect	7	322	8	323
rect	8	322	9	323
rect	9	322	10	323
rect	10	322	11	323
rect	11	322	12	323
rect	12	322	13	323
rect	13	322	14	323
rect	14	322	15	323
rect	15	322	16	323
rect	16	322	17	323
rect	17	322	18	323
rect	18	322	19	323
rect	19	322	20	323
rect	20	322	21	323
rect	21	322	22	323
rect	23	322	24	323
rect	24	322	25	323
rect	25	322	26	323
rect	26	322	27	323
rect	27	322	28	323
rect	28	322	29	323
rect	30	322	31	323
rect	31	322	32	323
rect	32	322	33	323
rect	33	322	34	323
rect	34	322	35	323
rect	35	322	36	323
rect	37	322	38	323
rect	38	322	39	323
rect	39	322	40	323
rect	40	322	41	323
rect	41	322	42	323
rect	42	322	43	323
rect	43	322	44	323
rect	44	322	45	323
rect	45	322	46	323
rect	46	322	47	323
rect	47	322	48	323
rect	48	322	49	323
rect	49	322	50	323
rect	50	322	51	323
rect	51	322	52	323
rect	52	322	53	323
rect	53	322	54	323
rect	54	322	55	323
rect	55	322	56	323
rect	56	322	57	323
rect	57	322	58	323
rect	58	322	59	323
rect	59	322	60	323
rect	60	322	61	323
rect	61	322	62	323
rect	62	322	63	323
rect	63	322	64	323
rect	64	322	65	323
rect	65	322	66	323
rect	66	322	67	323
rect	67	322	68	323
rect	68	322	69	323
rect	69	322	70	323
rect	70	322	71	323
rect	71	322	72	323
rect	72	322	73	323
rect	73	322	74	323
rect	74	322	75	323
rect	75	322	76	323
rect	76	322	77	323
rect	77	322	78	323
rect	78	322	79	323
rect	79	322	80	323
rect	80	322	81	323
rect	81	322	82	323
rect	82	322	83	323
rect	83	322	84	323
rect	84	322	85	323
rect	85	322	86	323
rect	86	322	87	323
rect	87	322	88	323
rect	88	322	89	323
rect	89	322	90	323
rect	90	322	91	323
rect	91	322	92	323
rect	92	322	93	323
rect	93	322	94	323
rect	94	322	95	323
rect	95	322	96	323
rect	96	322	97	323
rect	97	322	98	323
rect	98	322	99	323
rect	99	322	100	323
rect	100	322	101	323
rect	101	322	102	323
rect	102	322	103	323
rect	103	322	104	323
rect	104	322	105	323
rect	105	322	106	323
rect	106	322	107	323
rect	107	322	108	323
rect	108	322	109	323
rect	109	322	110	323
rect	110	322	111	323
rect	111	322	112	323
rect	112	322	113	323
rect	113	322	114	323
rect	114	322	115	323
rect	115	322	116	323
rect	116	322	117	323
rect	117	322	118	323
rect	118	322	119	323
rect	119	322	120	323
rect	120	322	121	323
rect	121	322	122	323
rect	122	322	123	323
rect	123	322	124	323
rect	124	322	125	323
rect	125	322	126	323
rect	126	322	127	323
rect	127	322	128	323
rect	128	322	129	323
rect	129	322	130	323
rect	130	322	131	323
rect	131	322	132	323
rect	132	322	133	323
rect	133	322	134	323
rect	134	322	135	323
rect	135	322	136	323
rect	136	322	137	323
rect	137	322	138	323
rect	138	322	139	323
rect	139	322	140	323
rect	140	322	141	323
rect	141	322	142	323
rect	142	322	143	323
rect	143	322	144	323
rect	144	322	145	323
rect	145	322	146	323
rect	146	322	147	323
rect	147	322	148	323
rect	148	322	149	323
rect	149	322	150	323
rect	150	322	151	323
rect	151	322	152	323
rect	152	322	153	323
rect	153	322	154	323
rect	154	322	155	323
rect	155	322	156	323
rect	156	322	157	323
rect	157	322	158	323
rect	158	322	159	323
rect	159	322	160	323
rect	160	322	161	323
rect	161	322	162	323
rect	162	322	163	323
rect	163	322	164	323
rect	164	322	165	323
rect	165	322	166	323
rect	166	322	167	323
rect	167	322	168	323
rect	168	322	169	323
rect	169	322	170	323
rect	170	322	171	323
rect	171	322	172	323
rect	172	322	173	323
rect	173	322	174	323
rect	174	322	175	323
rect	175	322	176	323
rect	176	322	177	323
rect	177	322	178	323
rect	178	322	179	323
rect	179	322	180	323
rect	180	322	181	323
rect	181	322	182	323
rect	182	322	183	323
rect	183	322	184	323
rect	184	322	185	323
rect	185	322	186	323
rect	186	322	187	323
rect	187	322	188	323
rect	188	322	189	323
rect	189	322	190	323
rect	190	322	191	323
rect	191	322	192	323
rect	192	322	193	323
rect	193	322	194	323
rect	194	322	195	323
rect	195	322	196	323
rect	196	322	197	323
rect	197	322	198	323
rect	198	322	199	323
rect	199	322	200	323
rect	200	322	201	323
rect	201	322	202	323
rect	202	322	203	323
rect	203	322	204	323
rect	204	322	205	323
rect	205	322	206	323
rect	206	322	207	323
rect	207	322	208	323
rect	208	322	209	323
rect	209	322	210	323
rect	210	322	211	323
rect	211	322	212	323
rect	212	322	213	323
rect	213	322	214	323
rect	214	322	215	323
rect	215	322	216	323
rect	216	322	217	323
rect	217	322	218	323
rect	218	322	219	323
rect	219	322	220	323
rect	220	322	221	323
rect	221	322	222	323
rect	222	322	223	323
rect	223	322	224	323
rect	224	322	225	323
rect	225	322	226	323
rect	226	322	227	323
rect	227	322	228	323
rect	228	322	229	323
rect	229	322	230	323
rect	230	322	231	323
rect	231	322	232	323
rect	232	322	233	323
rect	233	322	234	323
rect	234	322	235	323
rect	235	322	236	323
rect	236	322	237	323
rect	237	322	238	323
rect	238	322	239	323
rect	239	322	240	323
rect	240	322	241	323
rect	241	322	242	323
rect	242	322	243	323
rect	243	322	244	323
rect	244	322	245	323
rect	245	322	246	323
rect	246	322	247	323
rect	247	322	248	323
rect	248	322	249	323
rect	249	322	250	323
rect	250	322	251	323
rect	251	322	252	323
rect	252	322	253	323
rect	253	322	254	323
rect	254	322	255	323
rect	255	322	256	323
rect	256	322	257	323
rect	257	322	258	323
rect	258	322	259	323
rect	259	322	260	323
rect	260	322	261	323
rect	261	322	262	323
rect	262	322	263	323
rect	263	322	264	323
rect	264	322	265	323
rect	265	322	266	323
rect	266	322	267	323
rect	267	322	268	323
rect	268	322	269	323
rect	269	322	270	323
rect	270	322	271	323
rect	271	322	272	323
rect	272	322	273	323
rect	273	322	274	323
rect	274	322	275	323
rect	275	322	276	323
rect	276	322	277	323
rect	277	322	278	323
rect	278	322	279	323
rect	279	322	280	323
rect	280	322	281	323
rect	281	322	282	323
rect	282	322	283	323
rect	283	322	284	323
rect	284	322	285	323
rect	285	322	286	323
rect	286	322	287	323
rect	287	322	288	323
rect	288	322	289	323
rect	289	322	290	323
rect	290	322	291	323
rect	291	322	292	323
rect	292	322	293	323
rect	293	322	294	323
rect	294	322	295	323
rect	295	322	296	323
rect	296	322	297	323
rect	297	322	298	323
rect	298	322	299	323
rect	299	322	300	323
rect	300	322	301	323
rect	302	322	303	323
rect	303	322	304	323
rect	304	322	305	323
rect	305	322	306	323
rect	306	322	307	323
rect	307	322	308	323
rect	309	322	310	323
rect	310	322	311	323
rect	311	322	312	323
rect	312	322	313	323
rect	313	322	314	323
rect	314	322	315	323
rect	316	322	317	323
rect	317	322	318	323
rect	318	322	319	323
rect	319	322	320	323
rect	320	322	321	323
rect	321	322	322	323
rect	322	322	323	323
rect	323	322	324	323
rect	324	322	325	323
rect	325	322	326	323
rect	326	322	327	323
rect	327	322	328	323
rect	328	322	329	323
rect	329	322	330	323
rect	330	322	331	323
rect	331	322	332	323
rect	332	322	333	323
rect	333	322	334	323
rect	334	322	335	323
rect	335	322	336	323
rect	336	322	337	323
rect	337	322	338	323
rect	338	322	339	323
rect	339	322	340	323
rect	340	322	341	323
rect	341	322	342	323
rect	342	322	343	323
rect	344	322	345	323
rect	345	322	346	323
rect	346	322	347	323
rect	347	322	348	323
rect	348	322	349	323
rect	349	322	350	323
rect	351	322	352	323
rect	352	322	353	323
rect	353	322	354	323
rect	354	322	355	323
rect	355	322	356	323
rect	356	322	357	323
rect	357	322	358	323
rect	358	322	359	323
rect	359	322	360	323
rect	360	322	361	323
rect	361	322	362	323
rect	362	322	363	323
rect	363	322	364	323
rect	364	322	365	323
rect	365	322	366	323
rect	366	322	367	323
rect	367	322	368	323
rect	368	322	369	323
rect	369	322	370	323
rect	370	322	371	323
rect	371	322	372	323
rect	372	322	373	323
rect	373	322	374	323
rect	374	322	375	323
rect	375	322	376	323
rect	376	322	377	323
rect	377	322	378	323
rect	378	322	379	323
rect	379	322	380	323
rect	380	322	381	323
rect	381	322	382	323
rect	382	322	383	323
rect	383	322	384	323
rect	384	322	385	323
rect	385	322	386	323
rect	386	322	387	323
rect	387	322	388	323
rect	388	322	389	323
rect	389	322	390	323
rect	390	322	391	323
rect	391	322	392	323
rect	392	322	393	323
rect	393	322	394	323
rect	394	322	395	323
rect	395	322	396	323
rect	396	322	397	323
rect	397	322	398	323
rect	398	322	399	323
rect	399	322	400	323
rect	400	322	401	323
rect	401	322	402	323
rect	403	322	404	323
rect	404	322	405	323
rect	405	322	406	323
rect	406	322	407	323
rect	407	322	408	323
rect	408	322	409	323
rect	409	322	410	323
rect	410	322	411	323
rect	411	322	412	323
rect	412	322	413	323
rect	413	322	414	323
rect	414	322	415	323
rect	415	322	416	323
rect	416	322	417	323
rect	417	322	418	323
rect	418	322	419	323
rect	419	322	420	323
rect	420	322	421	323
rect	0	350	1	351
rect	1	350	2	351
rect	2	350	3	351
rect	3	350	4	351
rect	4	350	5	351
rect	5	350	6	351
rect	6	350	7	351
rect	7	350	8	351
rect	8	350	9	351
rect	9	350	10	351
rect	10	350	11	351
rect	11	350	12	351
rect	12	350	13	351
rect	13	350	14	351
rect	14	350	15	351
rect	16	350	17	351
rect	17	350	18	351
rect	18	350	19	351
rect	19	350	20	351
rect	20	350	21	351
rect	21	350	22	351
rect	23	350	24	351
rect	24	350	25	351
rect	25	350	26	351
rect	26	350	27	351
rect	27	350	28	351
rect	28	350	29	351
rect	30	350	31	351
rect	31	350	32	351
rect	32	350	33	351
rect	33	350	34	351
rect	34	350	35	351
rect	35	350	36	351
rect	37	350	38	351
rect	38	350	39	351
rect	39	350	40	351
rect	40	350	41	351
rect	41	350	42	351
rect	42	350	43	351
rect	44	350	45	351
rect	45	350	46	351
rect	46	350	47	351
rect	47	350	48	351
rect	48	350	49	351
rect	49	350	50	351
rect	50	350	51	351
rect	51	350	52	351
rect	52	350	53	351
rect	53	350	54	351
rect	54	350	55	351
rect	55	350	56	351
rect	56	350	57	351
rect	57	350	58	351
rect	58	350	59	351
rect	59	350	60	351
rect	60	350	61	351
rect	61	350	62	351
rect	62	350	63	351
rect	63	350	64	351
rect	64	350	65	351
rect	65	350	66	351
rect	66	350	67	351
rect	67	350	68	351
rect	68	350	69	351
rect	69	350	70	351
rect	70	350	71	351
rect	71	350	72	351
rect	72	350	73	351
rect	73	350	74	351
rect	74	350	75	351
rect	75	350	76	351
rect	76	350	77	351
rect	77	350	78	351
rect	78	350	79	351
rect	79	350	80	351
rect	80	350	81	351
rect	81	350	82	351
rect	82	350	83	351
rect	83	350	84	351
rect	84	350	85	351
rect	85	350	86	351
rect	86	350	87	351
rect	87	350	88	351
rect	88	350	89	351
rect	89	350	90	351
rect	90	350	91	351
rect	91	350	92	351
rect	92	350	93	351
rect	93	350	94	351
rect	94	350	95	351
rect	95	350	96	351
rect	96	350	97	351
rect	97	350	98	351
rect	98	350	99	351
rect	99	350	100	351
rect	100	350	101	351
rect	101	350	102	351
rect	102	350	103	351
rect	103	350	104	351
rect	104	350	105	351
rect	105	350	106	351
rect	106	350	107	351
rect	107	350	108	351
rect	108	350	109	351
rect	109	350	110	351
rect	110	350	111	351
rect	111	350	112	351
rect	112	350	113	351
rect	113	350	114	351
rect	114	350	115	351
rect	115	350	116	351
rect	116	350	117	351
rect	117	350	118	351
rect	118	350	119	351
rect	119	350	120	351
rect	120	350	121	351
rect	121	350	122	351
rect	122	350	123	351
rect	123	350	124	351
rect	124	350	125	351
rect	125	350	126	351
rect	126	350	127	351
rect	127	350	128	351
rect	128	350	129	351
rect	129	350	130	351
rect	130	350	131	351
rect	131	350	132	351
rect	132	350	133	351
rect	133	350	134	351
rect	134	350	135	351
rect	135	350	136	351
rect	136	350	137	351
rect	137	350	138	351
rect	138	350	139	351
rect	139	350	140	351
rect	140	350	141	351
rect	141	350	142	351
rect	142	350	143	351
rect	143	350	144	351
rect	144	350	145	351
rect	145	350	146	351
rect	146	350	147	351
rect	147	350	148	351
rect	148	350	149	351
rect	149	350	150	351
rect	150	350	151	351
rect	151	350	152	351
rect	152	350	153	351
rect	153	350	154	351
rect	154	350	155	351
rect	155	350	156	351
rect	156	350	157	351
rect	157	350	158	351
rect	158	350	159	351
rect	159	350	160	351
rect	160	350	161	351
rect	161	350	162	351
rect	162	350	163	351
rect	163	350	164	351
rect	164	350	165	351
rect	165	350	166	351
rect	166	350	167	351
rect	167	350	168	351
rect	168	350	169	351
rect	169	350	170	351
rect	170	350	171	351
rect	171	350	172	351
rect	172	350	173	351
rect	173	350	174	351
rect	174	350	175	351
rect	175	350	176	351
rect	176	350	177	351
rect	177	350	178	351
rect	178	350	179	351
rect	179	350	180	351
rect	180	350	181	351
rect	181	350	182	351
rect	182	350	183	351
rect	183	350	184	351
rect	184	350	185	351
rect	185	350	186	351
rect	186	350	187	351
rect	187	350	188	351
rect	188	350	189	351
rect	189	350	190	351
rect	190	350	191	351
rect	191	350	192	351
rect	192	350	193	351
rect	193	350	194	351
rect	194	350	195	351
rect	195	350	196	351
rect	196	350	197	351
rect	197	350	198	351
rect	198	350	199	351
rect	199	350	200	351
rect	200	350	201	351
rect	201	350	202	351
rect	202	350	203	351
rect	203	350	204	351
rect	204	350	205	351
rect	205	350	206	351
rect	206	350	207	351
rect	207	350	208	351
rect	208	350	209	351
rect	209	350	210	351
rect	210	350	211	351
rect	211	350	212	351
rect	212	350	213	351
rect	213	350	214	351
rect	214	350	215	351
rect	215	350	216	351
rect	216	350	217	351
rect	217	350	218	351
rect	219	350	220	351
rect	220	350	221	351
rect	221	350	222	351
rect	222	350	223	351
rect	223	350	224	351
rect	224	350	225	351
rect	225	350	226	351
rect	226	350	227	351
rect	227	350	228	351
rect	228	350	229	351
rect	229	350	230	351
rect	230	350	231	351
rect	231	350	232	351
rect	232	350	233	351
rect	233	350	234	351
rect	234	350	235	351
rect	235	350	236	351
rect	236	350	237	351
rect	237	350	238	351
rect	238	350	239	351
rect	239	350	240	351
rect	240	350	241	351
rect	241	350	242	351
rect	242	350	243	351
rect	243	350	244	351
rect	244	350	245	351
rect	245	350	246	351
rect	246	350	247	351
rect	247	350	248	351
rect	248	350	249	351
rect	249	350	250	351
rect	250	350	251	351
rect	251	350	252	351
rect	252	350	253	351
rect	253	350	254	351
rect	254	350	255	351
rect	255	350	256	351
rect	256	350	257	351
rect	257	350	258	351
rect	258	350	259	351
rect	259	350	260	351
rect	260	350	261	351
rect	261	350	262	351
rect	262	350	263	351
rect	263	350	264	351
rect	264	350	265	351
rect	265	350	266	351
rect	266	350	267	351
rect	267	350	268	351
rect	268	350	269	351
rect	269	350	270	351
rect	270	350	271	351
rect	271	350	272	351
rect	272	350	273	351
rect	273	350	274	351
rect	274	350	275	351
rect	275	350	276	351
rect	276	350	277	351
rect	277	350	278	351
rect	278	350	279	351
rect	279	350	280	351
rect	280	350	281	351
rect	281	350	282	351
rect	282	350	283	351
rect	283	350	284	351
rect	284	350	285	351
rect	285	350	286	351
rect	286	350	287	351
rect	287	350	288	351
rect	288	350	289	351
rect	289	350	290	351
rect	290	350	291	351
rect	291	350	292	351
rect	292	350	293	351
rect	293	350	294	351
rect	294	350	295	351
rect	295	350	296	351
rect	296	350	297	351
rect	298	350	299	351
rect	299	350	300	351
rect	300	350	301	351
rect	301	350	302	351
rect	302	350	303	351
rect	303	350	304	351
rect	304	350	305	351
rect	305	350	306	351
rect	306	350	307	351
rect	307	350	308	351
rect	308	350	309	351
rect	309	350	310	351
rect	310	350	311	351
rect	311	350	312	351
rect	312	350	313	351
rect	313	350	314	351
rect	314	350	315	351
rect	315	350	316	351
rect	316	350	317	351
rect	317	350	318	351
rect	318	350	319	351
rect	319	350	320	351
rect	320	350	321	351
rect	321	350	322	351
rect	322	350	323	351
rect	323	350	324	351
rect	324	350	325	351
rect	325	350	326	351
rect	326	350	327	351
rect	327	350	328	351
rect	328	350	329	351
rect	329	350	330	351
rect	330	350	331	351
rect	332	350	333	351
rect	333	350	334	351
rect	334	350	335	351
rect	335	350	336	351
rect	336	350	337	351
rect	337	350	338	351
rect	339	350	340	351
rect	340	350	341	351
rect	341	350	342	351
rect	342	350	343	351
rect	343	350	344	351
rect	344	350	345	351
rect	345	350	346	351
rect	346	350	347	351
rect	347	350	348	351
rect	348	350	349	351
rect	349	350	350	351
rect	350	350	351	351
rect	351	350	352	351
rect	352	350	353	351
rect	353	350	354	351
rect	354	350	355	351
rect	355	350	356	351
rect	356	350	357	351
rect	357	350	358	351
rect	358	350	359	351
rect	359	350	360	351
rect	360	350	361	351
rect	361	350	362	351
rect	362	350	363	351
rect	363	350	364	351
rect	364	350	365	351
rect	365	350	366	351
rect	367	350	368	351
rect	368	350	369	351
rect	369	350	370	351
rect	370	350	371	351
rect	371	350	372	351
rect	372	350	373	351
rect	374	350	375	351
rect	375	350	376	351
rect	376	350	377	351
rect	377	350	378	351
rect	378	350	379	351
rect	379	350	380	351
rect	381	350	382	351
rect	382	350	383	351
rect	383	350	384	351
rect	384	350	385	351
rect	385	350	386	351
rect	386	350	387	351
rect	388	350	389	351
rect	389	350	390	351
rect	390	350	391	351
rect	391	350	392	351
rect	392	350	393	351
rect	393	350	394	351
rect	394	350	395	351
rect	395	350	396	351
rect	396	350	397	351
rect	0	351	1	352
rect	1	351	2	352
rect	2	351	3	352
rect	3	351	4	352
rect	4	351	5	352
rect	5	351	6	352
rect	6	351	7	352
rect	7	351	8	352
rect	8	351	9	352
rect	9	351	10	352
rect	10	351	11	352
rect	11	351	12	352
rect	12	351	13	352
rect	13	351	14	352
rect	14	351	15	352
rect	16	351	17	352
rect	17	351	18	352
rect	18	351	19	352
rect	19	351	20	352
rect	20	351	21	352
rect	21	351	22	352
rect	23	351	24	352
rect	24	351	25	352
rect	25	351	26	352
rect	26	351	27	352
rect	27	351	28	352
rect	28	351	29	352
rect	30	351	31	352
rect	31	351	32	352
rect	32	351	33	352
rect	33	351	34	352
rect	34	351	35	352
rect	35	351	36	352
rect	37	351	38	352
rect	38	351	39	352
rect	39	351	40	352
rect	40	351	41	352
rect	41	351	42	352
rect	42	351	43	352
rect	44	351	45	352
rect	45	351	46	352
rect	46	351	47	352
rect	47	351	48	352
rect	48	351	49	352
rect	49	351	50	352
rect	50	351	51	352
rect	51	351	52	352
rect	52	351	53	352
rect	53	351	54	352
rect	54	351	55	352
rect	55	351	56	352
rect	56	351	57	352
rect	57	351	58	352
rect	58	351	59	352
rect	59	351	60	352
rect	60	351	61	352
rect	61	351	62	352
rect	62	351	63	352
rect	63	351	64	352
rect	64	351	65	352
rect	65	351	66	352
rect	66	351	67	352
rect	67	351	68	352
rect	68	351	69	352
rect	69	351	70	352
rect	70	351	71	352
rect	71	351	72	352
rect	72	351	73	352
rect	73	351	74	352
rect	74	351	75	352
rect	75	351	76	352
rect	76	351	77	352
rect	77	351	78	352
rect	78	351	79	352
rect	79	351	80	352
rect	80	351	81	352
rect	81	351	82	352
rect	82	351	83	352
rect	83	351	84	352
rect	84	351	85	352
rect	85	351	86	352
rect	86	351	87	352
rect	87	351	88	352
rect	88	351	89	352
rect	89	351	90	352
rect	90	351	91	352
rect	91	351	92	352
rect	92	351	93	352
rect	93	351	94	352
rect	94	351	95	352
rect	95	351	96	352
rect	96	351	97	352
rect	97	351	98	352
rect	98	351	99	352
rect	99	351	100	352
rect	100	351	101	352
rect	101	351	102	352
rect	102	351	103	352
rect	103	351	104	352
rect	104	351	105	352
rect	105	351	106	352
rect	106	351	107	352
rect	107	351	108	352
rect	108	351	109	352
rect	109	351	110	352
rect	110	351	111	352
rect	111	351	112	352
rect	112	351	113	352
rect	113	351	114	352
rect	114	351	115	352
rect	115	351	116	352
rect	116	351	117	352
rect	117	351	118	352
rect	118	351	119	352
rect	119	351	120	352
rect	120	351	121	352
rect	121	351	122	352
rect	122	351	123	352
rect	123	351	124	352
rect	124	351	125	352
rect	125	351	126	352
rect	126	351	127	352
rect	127	351	128	352
rect	128	351	129	352
rect	129	351	130	352
rect	130	351	131	352
rect	131	351	132	352
rect	132	351	133	352
rect	133	351	134	352
rect	134	351	135	352
rect	135	351	136	352
rect	136	351	137	352
rect	137	351	138	352
rect	138	351	139	352
rect	139	351	140	352
rect	140	351	141	352
rect	141	351	142	352
rect	142	351	143	352
rect	143	351	144	352
rect	144	351	145	352
rect	145	351	146	352
rect	146	351	147	352
rect	147	351	148	352
rect	148	351	149	352
rect	149	351	150	352
rect	150	351	151	352
rect	151	351	152	352
rect	152	351	153	352
rect	153	351	154	352
rect	154	351	155	352
rect	155	351	156	352
rect	156	351	157	352
rect	157	351	158	352
rect	158	351	159	352
rect	159	351	160	352
rect	160	351	161	352
rect	161	351	162	352
rect	162	351	163	352
rect	163	351	164	352
rect	164	351	165	352
rect	165	351	166	352
rect	166	351	167	352
rect	167	351	168	352
rect	168	351	169	352
rect	169	351	170	352
rect	170	351	171	352
rect	171	351	172	352
rect	172	351	173	352
rect	173	351	174	352
rect	174	351	175	352
rect	175	351	176	352
rect	176	351	177	352
rect	177	351	178	352
rect	178	351	179	352
rect	179	351	180	352
rect	180	351	181	352
rect	181	351	182	352
rect	182	351	183	352
rect	183	351	184	352
rect	184	351	185	352
rect	185	351	186	352
rect	186	351	187	352
rect	187	351	188	352
rect	188	351	189	352
rect	189	351	190	352
rect	190	351	191	352
rect	191	351	192	352
rect	192	351	193	352
rect	193	351	194	352
rect	194	351	195	352
rect	195	351	196	352
rect	196	351	197	352
rect	197	351	198	352
rect	198	351	199	352
rect	199	351	200	352
rect	200	351	201	352
rect	201	351	202	352
rect	202	351	203	352
rect	203	351	204	352
rect	204	351	205	352
rect	205	351	206	352
rect	206	351	207	352
rect	207	351	208	352
rect	208	351	209	352
rect	209	351	210	352
rect	210	351	211	352
rect	211	351	212	352
rect	212	351	213	352
rect	213	351	214	352
rect	214	351	215	352
rect	215	351	216	352
rect	216	351	217	352
rect	217	351	218	352
rect	219	351	220	352
rect	220	351	221	352
rect	221	351	222	352
rect	222	351	223	352
rect	223	351	224	352
rect	224	351	225	352
rect	225	351	226	352
rect	226	351	227	352
rect	227	351	228	352
rect	228	351	229	352
rect	229	351	230	352
rect	230	351	231	352
rect	231	351	232	352
rect	232	351	233	352
rect	233	351	234	352
rect	234	351	235	352
rect	235	351	236	352
rect	236	351	237	352
rect	237	351	238	352
rect	238	351	239	352
rect	239	351	240	352
rect	240	351	241	352
rect	241	351	242	352
rect	242	351	243	352
rect	243	351	244	352
rect	244	351	245	352
rect	245	351	246	352
rect	246	351	247	352
rect	247	351	248	352
rect	248	351	249	352
rect	249	351	250	352
rect	250	351	251	352
rect	251	351	252	352
rect	252	351	253	352
rect	253	351	254	352
rect	254	351	255	352
rect	255	351	256	352
rect	256	351	257	352
rect	257	351	258	352
rect	258	351	259	352
rect	259	351	260	352
rect	260	351	261	352
rect	261	351	262	352
rect	262	351	263	352
rect	263	351	264	352
rect	264	351	265	352
rect	265	351	266	352
rect	266	351	267	352
rect	267	351	268	352
rect	268	351	269	352
rect	269	351	270	352
rect	270	351	271	352
rect	271	351	272	352
rect	272	351	273	352
rect	273	351	274	352
rect	274	351	275	352
rect	275	351	276	352
rect	276	351	277	352
rect	277	351	278	352
rect	278	351	279	352
rect	279	351	280	352
rect	280	351	281	352
rect	281	351	282	352
rect	282	351	283	352
rect	283	351	284	352
rect	284	351	285	352
rect	285	351	286	352
rect	286	351	287	352
rect	287	351	288	352
rect	288	351	289	352
rect	289	351	290	352
rect	290	351	291	352
rect	291	351	292	352
rect	292	351	293	352
rect	293	351	294	352
rect	294	351	295	352
rect	295	351	296	352
rect	296	351	297	352
rect	298	351	299	352
rect	299	351	300	352
rect	300	351	301	352
rect	301	351	302	352
rect	302	351	303	352
rect	303	351	304	352
rect	304	351	305	352
rect	305	351	306	352
rect	306	351	307	352
rect	307	351	308	352
rect	308	351	309	352
rect	309	351	310	352
rect	310	351	311	352
rect	311	351	312	352
rect	312	351	313	352
rect	313	351	314	352
rect	314	351	315	352
rect	315	351	316	352
rect	316	351	317	352
rect	317	351	318	352
rect	318	351	319	352
rect	319	351	320	352
rect	320	351	321	352
rect	321	351	322	352
rect	322	351	323	352
rect	323	351	324	352
rect	324	351	325	352
rect	325	351	326	352
rect	326	351	327	352
rect	327	351	328	352
rect	328	351	329	352
rect	329	351	330	352
rect	330	351	331	352
rect	332	351	333	352
rect	333	351	334	352
rect	334	351	335	352
rect	335	351	336	352
rect	336	351	337	352
rect	337	351	338	352
rect	339	351	340	352
rect	340	351	341	352
rect	341	351	342	352
rect	342	351	343	352
rect	343	351	344	352
rect	344	351	345	352
rect	345	351	346	352
rect	346	351	347	352
rect	347	351	348	352
rect	348	351	349	352
rect	349	351	350	352
rect	350	351	351	352
rect	351	351	352	352
rect	352	351	353	352
rect	353	351	354	352
rect	354	351	355	352
rect	355	351	356	352
rect	356	351	357	352
rect	357	351	358	352
rect	358	351	359	352
rect	359	351	360	352
rect	360	351	361	352
rect	361	351	362	352
rect	362	351	363	352
rect	363	351	364	352
rect	364	351	365	352
rect	365	351	366	352
rect	367	351	368	352
rect	368	351	369	352
rect	369	351	370	352
rect	370	351	371	352
rect	371	351	372	352
rect	372	351	373	352
rect	374	351	375	352
rect	375	351	376	352
rect	376	351	377	352
rect	377	351	378	352
rect	378	351	379	352
rect	379	351	380	352
rect	381	351	382	352
rect	382	351	383	352
rect	383	351	384	352
rect	384	351	385	352
rect	385	351	386	352
rect	386	351	387	352
rect	388	351	389	352
rect	389	351	390	352
rect	390	351	391	352
rect	391	351	392	352
rect	392	351	393	352
rect	393	351	394	352
rect	394	351	395	352
rect	395	351	396	352
rect	396	351	397	352
rect	0	352	1	353
rect	1	352	2	353
rect	2	352	3	353
rect	3	352	4	353
rect	4	352	5	353
rect	5	352	6	353
rect	6	352	7	353
rect	7	352	8	353
rect	8	352	9	353
rect	9	352	10	353
rect	10	352	11	353
rect	11	352	12	353
rect	12	352	13	353
rect	13	352	14	353
rect	14	352	15	353
rect	16	352	17	353
rect	17	352	18	353
rect	18	352	19	353
rect	19	352	20	353
rect	20	352	21	353
rect	21	352	22	353
rect	23	352	24	353
rect	24	352	25	353
rect	25	352	26	353
rect	26	352	27	353
rect	27	352	28	353
rect	28	352	29	353
rect	30	352	31	353
rect	31	352	32	353
rect	32	352	33	353
rect	33	352	34	353
rect	34	352	35	353
rect	35	352	36	353
rect	37	352	38	353
rect	38	352	39	353
rect	39	352	40	353
rect	40	352	41	353
rect	41	352	42	353
rect	42	352	43	353
rect	44	352	45	353
rect	45	352	46	353
rect	46	352	47	353
rect	47	352	48	353
rect	48	352	49	353
rect	49	352	50	353
rect	50	352	51	353
rect	51	352	52	353
rect	52	352	53	353
rect	53	352	54	353
rect	54	352	55	353
rect	55	352	56	353
rect	56	352	57	353
rect	57	352	58	353
rect	58	352	59	353
rect	59	352	60	353
rect	60	352	61	353
rect	61	352	62	353
rect	62	352	63	353
rect	63	352	64	353
rect	64	352	65	353
rect	65	352	66	353
rect	66	352	67	353
rect	67	352	68	353
rect	68	352	69	353
rect	69	352	70	353
rect	70	352	71	353
rect	71	352	72	353
rect	72	352	73	353
rect	73	352	74	353
rect	74	352	75	353
rect	75	352	76	353
rect	76	352	77	353
rect	77	352	78	353
rect	78	352	79	353
rect	79	352	80	353
rect	80	352	81	353
rect	81	352	82	353
rect	82	352	83	353
rect	83	352	84	353
rect	84	352	85	353
rect	85	352	86	353
rect	86	352	87	353
rect	87	352	88	353
rect	88	352	89	353
rect	89	352	90	353
rect	90	352	91	353
rect	91	352	92	353
rect	92	352	93	353
rect	93	352	94	353
rect	94	352	95	353
rect	95	352	96	353
rect	96	352	97	353
rect	97	352	98	353
rect	98	352	99	353
rect	99	352	100	353
rect	100	352	101	353
rect	101	352	102	353
rect	102	352	103	353
rect	103	352	104	353
rect	104	352	105	353
rect	105	352	106	353
rect	106	352	107	353
rect	107	352	108	353
rect	108	352	109	353
rect	109	352	110	353
rect	110	352	111	353
rect	111	352	112	353
rect	112	352	113	353
rect	113	352	114	353
rect	114	352	115	353
rect	115	352	116	353
rect	116	352	117	353
rect	117	352	118	353
rect	118	352	119	353
rect	119	352	120	353
rect	120	352	121	353
rect	121	352	122	353
rect	122	352	123	353
rect	123	352	124	353
rect	124	352	125	353
rect	125	352	126	353
rect	126	352	127	353
rect	127	352	128	353
rect	128	352	129	353
rect	129	352	130	353
rect	130	352	131	353
rect	131	352	132	353
rect	132	352	133	353
rect	133	352	134	353
rect	134	352	135	353
rect	135	352	136	353
rect	136	352	137	353
rect	137	352	138	353
rect	138	352	139	353
rect	139	352	140	353
rect	140	352	141	353
rect	141	352	142	353
rect	142	352	143	353
rect	143	352	144	353
rect	144	352	145	353
rect	145	352	146	353
rect	146	352	147	353
rect	147	352	148	353
rect	148	352	149	353
rect	149	352	150	353
rect	150	352	151	353
rect	151	352	152	353
rect	152	352	153	353
rect	153	352	154	353
rect	154	352	155	353
rect	155	352	156	353
rect	156	352	157	353
rect	157	352	158	353
rect	158	352	159	353
rect	159	352	160	353
rect	160	352	161	353
rect	161	352	162	353
rect	162	352	163	353
rect	163	352	164	353
rect	164	352	165	353
rect	165	352	166	353
rect	166	352	167	353
rect	167	352	168	353
rect	168	352	169	353
rect	169	352	170	353
rect	170	352	171	353
rect	171	352	172	353
rect	172	352	173	353
rect	173	352	174	353
rect	174	352	175	353
rect	175	352	176	353
rect	176	352	177	353
rect	177	352	178	353
rect	178	352	179	353
rect	179	352	180	353
rect	180	352	181	353
rect	181	352	182	353
rect	182	352	183	353
rect	183	352	184	353
rect	184	352	185	353
rect	185	352	186	353
rect	186	352	187	353
rect	187	352	188	353
rect	188	352	189	353
rect	189	352	190	353
rect	190	352	191	353
rect	191	352	192	353
rect	192	352	193	353
rect	193	352	194	353
rect	194	352	195	353
rect	195	352	196	353
rect	196	352	197	353
rect	197	352	198	353
rect	198	352	199	353
rect	199	352	200	353
rect	200	352	201	353
rect	201	352	202	353
rect	202	352	203	353
rect	203	352	204	353
rect	204	352	205	353
rect	205	352	206	353
rect	206	352	207	353
rect	207	352	208	353
rect	208	352	209	353
rect	209	352	210	353
rect	210	352	211	353
rect	211	352	212	353
rect	212	352	213	353
rect	213	352	214	353
rect	214	352	215	353
rect	215	352	216	353
rect	216	352	217	353
rect	217	352	218	353
rect	219	352	220	353
rect	220	352	221	353
rect	221	352	222	353
rect	222	352	223	353
rect	223	352	224	353
rect	224	352	225	353
rect	225	352	226	353
rect	226	352	227	353
rect	227	352	228	353
rect	228	352	229	353
rect	229	352	230	353
rect	230	352	231	353
rect	231	352	232	353
rect	232	352	233	353
rect	233	352	234	353
rect	234	352	235	353
rect	235	352	236	353
rect	236	352	237	353
rect	237	352	238	353
rect	238	352	239	353
rect	239	352	240	353
rect	240	352	241	353
rect	241	352	242	353
rect	242	352	243	353
rect	243	352	244	353
rect	244	352	245	353
rect	245	352	246	353
rect	246	352	247	353
rect	247	352	248	353
rect	248	352	249	353
rect	249	352	250	353
rect	250	352	251	353
rect	251	352	252	353
rect	252	352	253	353
rect	253	352	254	353
rect	254	352	255	353
rect	255	352	256	353
rect	256	352	257	353
rect	257	352	258	353
rect	258	352	259	353
rect	259	352	260	353
rect	260	352	261	353
rect	261	352	262	353
rect	262	352	263	353
rect	263	352	264	353
rect	264	352	265	353
rect	265	352	266	353
rect	266	352	267	353
rect	267	352	268	353
rect	268	352	269	353
rect	269	352	270	353
rect	270	352	271	353
rect	271	352	272	353
rect	272	352	273	353
rect	273	352	274	353
rect	274	352	275	353
rect	275	352	276	353
rect	276	352	277	353
rect	277	352	278	353
rect	278	352	279	353
rect	279	352	280	353
rect	280	352	281	353
rect	281	352	282	353
rect	282	352	283	353
rect	283	352	284	353
rect	284	352	285	353
rect	285	352	286	353
rect	286	352	287	353
rect	287	352	288	353
rect	288	352	289	353
rect	289	352	290	353
rect	290	352	291	353
rect	291	352	292	353
rect	292	352	293	353
rect	293	352	294	353
rect	294	352	295	353
rect	295	352	296	353
rect	296	352	297	353
rect	298	352	299	353
rect	299	352	300	353
rect	300	352	301	353
rect	301	352	302	353
rect	302	352	303	353
rect	303	352	304	353
rect	304	352	305	353
rect	305	352	306	353
rect	306	352	307	353
rect	307	352	308	353
rect	308	352	309	353
rect	309	352	310	353
rect	310	352	311	353
rect	311	352	312	353
rect	312	352	313	353
rect	313	352	314	353
rect	314	352	315	353
rect	315	352	316	353
rect	316	352	317	353
rect	317	352	318	353
rect	318	352	319	353
rect	319	352	320	353
rect	320	352	321	353
rect	321	352	322	353
rect	322	352	323	353
rect	323	352	324	353
rect	324	352	325	353
rect	325	352	326	353
rect	326	352	327	353
rect	327	352	328	353
rect	328	352	329	353
rect	329	352	330	353
rect	330	352	331	353
rect	332	352	333	353
rect	333	352	334	353
rect	334	352	335	353
rect	335	352	336	353
rect	336	352	337	353
rect	337	352	338	353
rect	339	352	340	353
rect	340	352	341	353
rect	341	352	342	353
rect	342	352	343	353
rect	343	352	344	353
rect	344	352	345	353
rect	345	352	346	353
rect	346	352	347	353
rect	347	352	348	353
rect	348	352	349	353
rect	349	352	350	353
rect	350	352	351	353
rect	351	352	352	353
rect	352	352	353	353
rect	353	352	354	353
rect	354	352	355	353
rect	355	352	356	353
rect	356	352	357	353
rect	357	352	358	353
rect	358	352	359	353
rect	359	352	360	353
rect	360	352	361	353
rect	361	352	362	353
rect	362	352	363	353
rect	363	352	364	353
rect	364	352	365	353
rect	365	352	366	353
rect	367	352	368	353
rect	368	352	369	353
rect	369	352	370	353
rect	370	352	371	353
rect	371	352	372	353
rect	372	352	373	353
rect	374	352	375	353
rect	375	352	376	353
rect	376	352	377	353
rect	377	352	378	353
rect	378	352	379	353
rect	379	352	380	353
rect	381	352	382	353
rect	382	352	383	353
rect	383	352	384	353
rect	384	352	385	353
rect	385	352	386	353
rect	386	352	387	353
rect	388	352	389	353
rect	389	352	390	353
rect	390	352	391	353
rect	391	352	392	353
rect	392	352	393	353
rect	393	352	394	353
rect	394	352	395	353
rect	395	352	396	353
rect	396	352	397	353
rect	0	353	1	354
rect	1	353	2	354
rect	2	353	3	354
rect	3	353	4	354
rect	4	353	5	354
rect	5	353	6	354
rect	6	353	7	354
rect	7	353	8	354
rect	8	353	9	354
rect	9	353	10	354
rect	10	353	11	354
rect	11	353	12	354
rect	12	353	13	354
rect	13	353	14	354
rect	14	353	15	354
rect	16	353	17	354
rect	17	353	18	354
rect	18	353	19	354
rect	19	353	20	354
rect	20	353	21	354
rect	21	353	22	354
rect	23	353	24	354
rect	24	353	25	354
rect	25	353	26	354
rect	26	353	27	354
rect	27	353	28	354
rect	28	353	29	354
rect	30	353	31	354
rect	31	353	32	354
rect	32	353	33	354
rect	33	353	34	354
rect	34	353	35	354
rect	35	353	36	354
rect	37	353	38	354
rect	38	353	39	354
rect	39	353	40	354
rect	40	353	41	354
rect	41	353	42	354
rect	42	353	43	354
rect	44	353	45	354
rect	45	353	46	354
rect	46	353	47	354
rect	47	353	48	354
rect	48	353	49	354
rect	49	353	50	354
rect	50	353	51	354
rect	51	353	52	354
rect	52	353	53	354
rect	53	353	54	354
rect	54	353	55	354
rect	55	353	56	354
rect	56	353	57	354
rect	57	353	58	354
rect	58	353	59	354
rect	59	353	60	354
rect	60	353	61	354
rect	61	353	62	354
rect	62	353	63	354
rect	63	353	64	354
rect	64	353	65	354
rect	65	353	66	354
rect	66	353	67	354
rect	67	353	68	354
rect	68	353	69	354
rect	69	353	70	354
rect	70	353	71	354
rect	71	353	72	354
rect	72	353	73	354
rect	73	353	74	354
rect	74	353	75	354
rect	75	353	76	354
rect	76	353	77	354
rect	77	353	78	354
rect	78	353	79	354
rect	79	353	80	354
rect	80	353	81	354
rect	81	353	82	354
rect	82	353	83	354
rect	83	353	84	354
rect	84	353	85	354
rect	85	353	86	354
rect	86	353	87	354
rect	87	353	88	354
rect	88	353	89	354
rect	89	353	90	354
rect	90	353	91	354
rect	91	353	92	354
rect	92	353	93	354
rect	93	353	94	354
rect	94	353	95	354
rect	95	353	96	354
rect	96	353	97	354
rect	97	353	98	354
rect	98	353	99	354
rect	99	353	100	354
rect	100	353	101	354
rect	101	353	102	354
rect	102	353	103	354
rect	103	353	104	354
rect	104	353	105	354
rect	105	353	106	354
rect	106	353	107	354
rect	107	353	108	354
rect	108	353	109	354
rect	109	353	110	354
rect	110	353	111	354
rect	111	353	112	354
rect	112	353	113	354
rect	113	353	114	354
rect	114	353	115	354
rect	115	353	116	354
rect	116	353	117	354
rect	117	353	118	354
rect	118	353	119	354
rect	119	353	120	354
rect	120	353	121	354
rect	121	353	122	354
rect	122	353	123	354
rect	123	353	124	354
rect	124	353	125	354
rect	125	353	126	354
rect	126	353	127	354
rect	127	353	128	354
rect	128	353	129	354
rect	129	353	130	354
rect	130	353	131	354
rect	131	353	132	354
rect	132	353	133	354
rect	133	353	134	354
rect	134	353	135	354
rect	135	353	136	354
rect	136	353	137	354
rect	137	353	138	354
rect	138	353	139	354
rect	139	353	140	354
rect	140	353	141	354
rect	141	353	142	354
rect	142	353	143	354
rect	143	353	144	354
rect	144	353	145	354
rect	145	353	146	354
rect	146	353	147	354
rect	147	353	148	354
rect	148	353	149	354
rect	149	353	150	354
rect	150	353	151	354
rect	151	353	152	354
rect	152	353	153	354
rect	153	353	154	354
rect	154	353	155	354
rect	155	353	156	354
rect	156	353	157	354
rect	157	353	158	354
rect	158	353	159	354
rect	159	353	160	354
rect	160	353	161	354
rect	161	353	162	354
rect	162	353	163	354
rect	163	353	164	354
rect	164	353	165	354
rect	165	353	166	354
rect	166	353	167	354
rect	167	353	168	354
rect	168	353	169	354
rect	169	353	170	354
rect	170	353	171	354
rect	171	353	172	354
rect	172	353	173	354
rect	173	353	174	354
rect	174	353	175	354
rect	175	353	176	354
rect	176	353	177	354
rect	177	353	178	354
rect	178	353	179	354
rect	179	353	180	354
rect	180	353	181	354
rect	181	353	182	354
rect	182	353	183	354
rect	183	353	184	354
rect	184	353	185	354
rect	185	353	186	354
rect	186	353	187	354
rect	187	353	188	354
rect	188	353	189	354
rect	189	353	190	354
rect	190	353	191	354
rect	191	353	192	354
rect	192	353	193	354
rect	193	353	194	354
rect	194	353	195	354
rect	195	353	196	354
rect	196	353	197	354
rect	197	353	198	354
rect	198	353	199	354
rect	199	353	200	354
rect	200	353	201	354
rect	201	353	202	354
rect	202	353	203	354
rect	203	353	204	354
rect	204	353	205	354
rect	205	353	206	354
rect	206	353	207	354
rect	207	353	208	354
rect	208	353	209	354
rect	209	353	210	354
rect	210	353	211	354
rect	211	353	212	354
rect	212	353	213	354
rect	213	353	214	354
rect	214	353	215	354
rect	215	353	216	354
rect	216	353	217	354
rect	217	353	218	354
rect	219	353	220	354
rect	220	353	221	354
rect	221	353	222	354
rect	222	353	223	354
rect	223	353	224	354
rect	224	353	225	354
rect	225	353	226	354
rect	226	353	227	354
rect	227	353	228	354
rect	228	353	229	354
rect	229	353	230	354
rect	230	353	231	354
rect	231	353	232	354
rect	232	353	233	354
rect	233	353	234	354
rect	234	353	235	354
rect	235	353	236	354
rect	236	353	237	354
rect	237	353	238	354
rect	238	353	239	354
rect	239	353	240	354
rect	240	353	241	354
rect	241	353	242	354
rect	242	353	243	354
rect	243	353	244	354
rect	244	353	245	354
rect	245	353	246	354
rect	246	353	247	354
rect	247	353	248	354
rect	248	353	249	354
rect	249	353	250	354
rect	250	353	251	354
rect	251	353	252	354
rect	252	353	253	354
rect	253	353	254	354
rect	254	353	255	354
rect	255	353	256	354
rect	256	353	257	354
rect	257	353	258	354
rect	258	353	259	354
rect	259	353	260	354
rect	260	353	261	354
rect	261	353	262	354
rect	262	353	263	354
rect	263	353	264	354
rect	264	353	265	354
rect	265	353	266	354
rect	266	353	267	354
rect	267	353	268	354
rect	268	353	269	354
rect	269	353	270	354
rect	270	353	271	354
rect	271	353	272	354
rect	272	353	273	354
rect	273	353	274	354
rect	274	353	275	354
rect	275	353	276	354
rect	276	353	277	354
rect	277	353	278	354
rect	278	353	279	354
rect	279	353	280	354
rect	280	353	281	354
rect	281	353	282	354
rect	282	353	283	354
rect	283	353	284	354
rect	284	353	285	354
rect	285	353	286	354
rect	286	353	287	354
rect	287	353	288	354
rect	288	353	289	354
rect	289	353	290	354
rect	290	353	291	354
rect	291	353	292	354
rect	292	353	293	354
rect	293	353	294	354
rect	294	353	295	354
rect	295	353	296	354
rect	296	353	297	354
rect	298	353	299	354
rect	299	353	300	354
rect	300	353	301	354
rect	301	353	302	354
rect	302	353	303	354
rect	303	353	304	354
rect	304	353	305	354
rect	305	353	306	354
rect	306	353	307	354
rect	307	353	308	354
rect	308	353	309	354
rect	309	353	310	354
rect	310	353	311	354
rect	311	353	312	354
rect	312	353	313	354
rect	313	353	314	354
rect	314	353	315	354
rect	315	353	316	354
rect	316	353	317	354
rect	317	353	318	354
rect	318	353	319	354
rect	319	353	320	354
rect	320	353	321	354
rect	321	353	322	354
rect	322	353	323	354
rect	323	353	324	354
rect	324	353	325	354
rect	325	353	326	354
rect	326	353	327	354
rect	327	353	328	354
rect	328	353	329	354
rect	329	353	330	354
rect	330	353	331	354
rect	332	353	333	354
rect	333	353	334	354
rect	334	353	335	354
rect	335	353	336	354
rect	336	353	337	354
rect	337	353	338	354
rect	339	353	340	354
rect	340	353	341	354
rect	341	353	342	354
rect	342	353	343	354
rect	343	353	344	354
rect	344	353	345	354
rect	345	353	346	354
rect	346	353	347	354
rect	347	353	348	354
rect	348	353	349	354
rect	349	353	350	354
rect	350	353	351	354
rect	351	353	352	354
rect	352	353	353	354
rect	353	353	354	354
rect	354	353	355	354
rect	355	353	356	354
rect	356	353	357	354
rect	357	353	358	354
rect	358	353	359	354
rect	359	353	360	354
rect	360	353	361	354
rect	361	353	362	354
rect	362	353	363	354
rect	363	353	364	354
rect	364	353	365	354
rect	365	353	366	354
rect	367	353	368	354
rect	368	353	369	354
rect	369	353	370	354
rect	370	353	371	354
rect	371	353	372	354
rect	372	353	373	354
rect	374	353	375	354
rect	375	353	376	354
rect	376	353	377	354
rect	377	353	378	354
rect	378	353	379	354
rect	379	353	380	354
rect	381	353	382	354
rect	382	353	383	354
rect	383	353	384	354
rect	384	353	385	354
rect	385	353	386	354
rect	386	353	387	354
rect	388	353	389	354
rect	389	353	390	354
rect	390	353	391	354
rect	391	353	392	354
rect	392	353	393	354
rect	393	353	394	354
rect	394	353	395	354
rect	395	353	396	354
rect	396	353	397	354
rect	0	354	1	355
rect	1	354	2	355
rect	2	354	3	355
rect	3	354	4	355
rect	4	354	5	355
rect	5	354	6	355
rect	6	354	7	355
rect	7	354	8	355
rect	8	354	9	355
rect	9	354	10	355
rect	10	354	11	355
rect	11	354	12	355
rect	12	354	13	355
rect	13	354	14	355
rect	14	354	15	355
rect	16	354	17	355
rect	17	354	18	355
rect	18	354	19	355
rect	19	354	20	355
rect	20	354	21	355
rect	21	354	22	355
rect	23	354	24	355
rect	24	354	25	355
rect	25	354	26	355
rect	26	354	27	355
rect	27	354	28	355
rect	28	354	29	355
rect	30	354	31	355
rect	31	354	32	355
rect	32	354	33	355
rect	33	354	34	355
rect	34	354	35	355
rect	35	354	36	355
rect	37	354	38	355
rect	38	354	39	355
rect	39	354	40	355
rect	40	354	41	355
rect	41	354	42	355
rect	42	354	43	355
rect	44	354	45	355
rect	45	354	46	355
rect	46	354	47	355
rect	47	354	48	355
rect	48	354	49	355
rect	49	354	50	355
rect	50	354	51	355
rect	51	354	52	355
rect	52	354	53	355
rect	53	354	54	355
rect	54	354	55	355
rect	55	354	56	355
rect	56	354	57	355
rect	57	354	58	355
rect	58	354	59	355
rect	59	354	60	355
rect	60	354	61	355
rect	61	354	62	355
rect	62	354	63	355
rect	63	354	64	355
rect	64	354	65	355
rect	65	354	66	355
rect	66	354	67	355
rect	67	354	68	355
rect	68	354	69	355
rect	69	354	70	355
rect	70	354	71	355
rect	71	354	72	355
rect	72	354	73	355
rect	73	354	74	355
rect	74	354	75	355
rect	75	354	76	355
rect	76	354	77	355
rect	77	354	78	355
rect	78	354	79	355
rect	79	354	80	355
rect	80	354	81	355
rect	81	354	82	355
rect	82	354	83	355
rect	83	354	84	355
rect	84	354	85	355
rect	85	354	86	355
rect	86	354	87	355
rect	87	354	88	355
rect	88	354	89	355
rect	89	354	90	355
rect	90	354	91	355
rect	91	354	92	355
rect	92	354	93	355
rect	93	354	94	355
rect	94	354	95	355
rect	95	354	96	355
rect	96	354	97	355
rect	97	354	98	355
rect	98	354	99	355
rect	99	354	100	355
rect	100	354	101	355
rect	101	354	102	355
rect	102	354	103	355
rect	103	354	104	355
rect	104	354	105	355
rect	105	354	106	355
rect	106	354	107	355
rect	107	354	108	355
rect	108	354	109	355
rect	109	354	110	355
rect	110	354	111	355
rect	111	354	112	355
rect	112	354	113	355
rect	113	354	114	355
rect	114	354	115	355
rect	115	354	116	355
rect	116	354	117	355
rect	117	354	118	355
rect	118	354	119	355
rect	119	354	120	355
rect	120	354	121	355
rect	121	354	122	355
rect	122	354	123	355
rect	123	354	124	355
rect	124	354	125	355
rect	125	354	126	355
rect	126	354	127	355
rect	127	354	128	355
rect	128	354	129	355
rect	129	354	130	355
rect	130	354	131	355
rect	131	354	132	355
rect	132	354	133	355
rect	133	354	134	355
rect	134	354	135	355
rect	135	354	136	355
rect	136	354	137	355
rect	137	354	138	355
rect	138	354	139	355
rect	139	354	140	355
rect	140	354	141	355
rect	141	354	142	355
rect	142	354	143	355
rect	143	354	144	355
rect	144	354	145	355
rect	145	354	146	355
rect	146	354	147	355
rect	147	354	148	355
rect	148	354	149	355
rect	149	354	150	355
rect	150	354	151	355
rect	151	354	152	355
rect	152	354	153	355
rect	153	354	154	355
rect	154	354	155	355
rect	155	354	156	355
rect	156	354	157	355
rect	157	354	158	355
rect	158	354	159	355
rect	159	354	160	355
rect	160	354	161	355
rect	161	354	162	355
rect	162	354	163	355
rect	163	354	164	355
rect	164	354	165	355
rect	165	354	166	355
rect	166	354	167	355
rect	167	354	168	355
rect	168	354	169	355
rect	169	354	170	355
rect	170	354	171	355
rect	171	354	172	355
rect	172	354	173	355
rect	173	354	174	355
rect	174	354	175	355
rect	175	354	176	355
rect	176	354	177	355
rect	177	354	178	355
rect	178	354	179	355
rect	179	354	180	355
rect	180	354	181	355
rect	181	354	182	355
rect	182	354	183	355
rect	183	354	184	355
rect	184	354	185	355
rect	185	354	186	355
rect	186	354	187	355
rect	187	354	188	355
rect	188	354	189	355
rect	189	354	190	355
rect	190	354	191	355
rect	191	354	192	355
rect	192	354	193	355
rect	193	354	194	355
rect	194	354	195	355
rect	195	354	196	355
rect	196	354	197	355
rect	197	354	198	355
rect	198	354	199	355
rect	199	354	200	355
rect	200	354	201	355
rect	201	354	202	355
rect	202	354	203	355
rect	203	354	204	355
rect	204	354	205	355
rect	205	354	206	355
rect	206	354	207	355
rect	207	354	208	355
rect	208	354	209	355
rect	209	354	210	355
rect	210	354	211	355
rect	211	354	212	355
rect	212	354	213	355
rect	213	354	214	355
rect	214	354	215	355
rect	215	354	216	355
rect	216	354	217	355
rect	217	354	218	355
rect	219	354	220	355
rect	220	354	221	355
rect	221	354	222	355
rect	222	354	223	355
rect	223	354	224	355
rect	224	354	225	355
rect	225	354	226	355
rect	226	354	227	355
rect	227	354	228	355
rect	228	354	229	355
rect	229	354	230	355
rect	230	354	231	355
rect	231	354	232	355
rect	232	354	233	355
rect	233	354	234	355
rect	234	354	235	355
rect	235	354	236	355
rect	236	354	237	355
rect	237	354	238	355
rect	238	354	239	355
rect	239	354	240	355
rect	240	354	241	355
rect	241	354	242	355
rect	242	354	243	355
rect	243	354	244	355
rect	244	354	245	355
rect	245	354	246	355
rect	246	354	247	355
rect	247	354	248	355
rect	248	354	249	355
rect	249	354	250	355
rect	250	354	251	355
rect	251	354	252	355
rect	252	354	253	355
rect	253	354	254	355
rect	254	354	255	355
rect	255	354	256	355
rect	256	354	257	355
rect	257	354	258	355
rect	258	354	259	355
rect	259	354	260	355
rect	260	354	261	355
rect	261	354	262	355
rect	262	354	263	355
rect	263	354	264	355
rect	264	354	265	355
rect	265	354	266	355
rect	266	354	267	355
rect	267	354	268	355
rect	268	354	269	355
rect	269	354	270	355
rect	270	354	271	355
rect	271	354	272	355
rect	272	354	273	355
rect	273	354	274	355
rect	274	354	275	355
rect	275	354	276	355
rect	276	354	277	355
rect	277	354	278	355
rect	278	354	279	355
rect	279	354	280	355
rect	280	354	281	355
rect	281	354	282	355
rect	282	354	283	355
rect	283	354	284	355
rect	284	354	285	355
rect	285	354	286	355
rect	286	354	287	355
rect	287	354	288	355
rect	288	354	289	355
rect	289	354	290	355
rect	290	354	291	355
rect	291	354	292	355
rect	292	354	293	355
rect	293	354	294	355
rect	294	354	295	355
rect	295	354	296	355
rect	296	354	297	355
rect	298	354	299	355
rect	299	354	300	355
rect	300	354	301	355
rect	301	354	302	355
rect	302	354	303	355
rect	303	354	304	355
rect	304	354	305	355
rect	305	354	306	355
rect	306	354	307	355
rect	307	354	308	355
rect	308	354	309	355
rect	309	354	310	355
rect	310	354	311	355
rect	311	354	312	355
rect	312	354	313	355
rect	313	354	314	355
rect	314	354	315	355
rect	315	354	316	355
rect	316	354	317	355
rect	317	354	318	355
rect	318	354	319	355
rect	319	354	320	355
rect	320	354	321	355
rect	321	354	322	355
rect	322	354	323	355
rect	323	354	324	355
rect	324	354	325	355
rect	325	354	326	355
rect	326	354	327	355
rect	327	354	328	355
rect	328	354	329	355
rect	329	354	330	355
rect	330	354	331	355
rect	332	354	333	355
rect	333	354	334	355
rect	334	354	335	355
rect	335	354	336	355
rect	336	354	337	355
rect	337	354	338	355
rect	339	354	340	355
rect	340	354	341	355
rect	341	354	342	355
rect	342	354	343	355
rect	343	354	344	355
rect	344	354	345	355
rect	345	354	346	355
rect	346	354	347	355
rect	347	354	348	355
rect	348	354	349	355
rect	349	354	350	355
rect	350	354	351	355
rect	351	354	352	355
rect	352	354	353	355
rect	353	354	354	355
rect	354	354	355	355
rect	355	354	356	355
rect	356	354	357	355
rect	357	354	358	355
rect	358	354	359	355
rect	359	354	360	355
rect	360	354	361	355
rect	361	354	362	355
rect	362	354	363	355
rect	363	354	364	355
rect	364	354	365	355
rect	365	354	366	355
rect	367	354	368	355
rect	368	354	369	355
rect	369	354	370	355
rect	370	354	371	355
rect	371	354	372	355
rect	372	354	373	355
rect	374	354	375	355
rect	375	354	376	355
rect	376	354	377	355
rect	377	354	378	355
rect	378	354	379	355
rect	379	354	380	355
rect	381	354	382	355
rect	382	354	383	355
rect	383	354	384	355
rect	384	354	385	355
rect	385	354	386	355
rect	386	354	387	355
rect	388	354	389	355
rect	389	354	390	355
rect	390	354	391	355
rect	391	354	392	355
rect	392	354	393	355
rect	393	354	394	355
rect	394	354	395	355
rect	395	354	396	355
rect	396	354	397	355
rect	0	355	1	356
rect	1	355	2	356
rect	2	355	3	356
rect	3	355	4	356
rect	4	355	5	356
rect	5	355	6	356
rect	6	355	7	356
rect	7	355	8	356
rect	8	355	9	356
rect	9	355	10	356
rect	10	355	11	356
rect	11	355	12	356
rect	12	355	13	356
rect	13	355	14	356
rect	14	355	15	356
rect	16	355	17	356
rect	17	355	18	356
rect	18	355	19	356
rect	19	355	20	356
rect	20	355	21	356
rect	21	355	22	356
rect	23	355	24	356
rect	24	355	25	356
rect	25	355	26	356
rect	26	355	27	356
rect	27	355	28	356
rect	28	355	29	356
rect	30	355	31	356
rect	31	355	32	356
rect	32	355	33	356
rect	33	355	34	356
rect	34	355	35	356
rect	35	355	36	356
rect	37	355	38	356
rect	38	355	39	356
rect	39	355	40	356
rect	40	355	41	356
rect	41	355	42	356
rect	42	355	43	356
rect	44	355	45	356
rect	45	355	46	356
rect	46	355	47	356
rect	47	355	48	356
rect	48	355	49	356
rect	49	355	50	356
rect	50	355	51	356
rect	51	355	52	356
rect	52	355	53	356
rect	53	355	54	356
rect	54	355	55	356
rect	55	355	56	356
rect	56	355	57	356
rect	57	355	58	356
rect	58	355	59	356
rect	59	355	60	356
rect	60	355	61	356
rect	61	355	62	356
rect	62	355	63	356
rect	63	355	64	356
rect	64	355	65	356
rect	65	355	66	356
rect	66	355	67	356
rect	67	355	68	356
rect	68	355	69	356
rect	69	355	70	356
rect	70	355	71	356
rect	71	355	72	356
rect	72	355	73	356
rect	73	355	74	356
rect	74	355	75	356
rect	75	355	76	356
rect	76	355	77	356
rect	77	355	78	356
rect	78	355	79	356
rect	79	355	80	356
rect	80	355	81	356
rect	81	355	82	356
rect	82	355	83	356
rect	83	355	84	356
rect	84	355	85	356
rect	85	355	86	356
rect	86	355	87	356
rect	87	355	88	356
rect	88	355	89	356
rect	89	355	90	356
rect	90	355	91	356
rect	91	355	92	356
rect	92	355	93	356
rect	93	355	94	356
rect	94	355	95	356
rect	95	355	96	356
rect	96	355	97	356
rect	97	355	98	356
rect	98	355	99	356
rect	99	355	100	356
rect	100	355	101	356
rect	101	355	102	356
rect	102	355	103	356
rect	103	355	104	356
rect	104	355	105	356
rect	105	355	106	356
rect	106	355	107	356
rect	107	355	108	356
rect	108	355	109	356
rect	109	355	110	356
rect	110	355	111	356
rect	111	355	112	356
rect	112	355	113	356
rect	113	355	114	356
rect	114	355	115	356
rect	115	355	116	356
rect	116	355	117	356
rect	117	355	118	356
rect	118	355	119	356
rect	119	355	120	356
rect	120	355	121	356
rect	121	355	122	356
rect	122	355	123	356
rect	123	355	124	356
rect	124	355	125	356
rect	125	355	126	356
rect	126	355	127	356
rect	127	355	128	356
rect	128	355	129	356
rect	129	355	130	356
rect	130	355	131	356
rect	131	355	132	356
rect	132	355	133	356
rect	133	355	134	356
rect	134	355	135	356
rect	135	355	136	356
rect	136	355	137	356
rect	137	355	138	356
rect	138	355	139	356
rect	139	355	140	356
rect	140	355	141	356
rect	141	355	142	356
rect	142	355	143	356
rect	143	355	144	356
rect	144	355	145	356
rect	145	355	146	356
rect	146	355	147	356
rect	147	355	148	356
rect	148	355	149	356
rect	149	355	150	356
rect	150	355	151	356
rect	151	355	152	356
rect	152	355	153	356
rect	153	355	154	356
rect	154	355	155	356
rect	155	355	156	356
rect	156	355	157	356
rect	157	355	158	356
rect	158	355	159	356
rect	159	355	160	356
rect	160	355	161	356
rect	161	355	162	356
rect	162	355	163	356
rect	163	355	164	356
rect	164	355	165	356
rect	165	355	166	356
rect	166	355	167	356
rect	167	355	168	356
rect	168	355	169	356
rect	169	355	170	356
rect	170	355	171	356
rect	171	355	172	356
rect	172	355	173	356
rect	173	355	174	356
rect	174	355	175	356
rect	175	355	176	356
rect	176	355	177	356
rect	177	355	178	356
rect	178	355	179	356
rect	179	355	180	356
rect	180	355	181	356
rect	181	355	182	356
rect	182	355	183	356
rect	183	355	184	356
rect	184	355	185	356
rect	185	355	186	356
rect	186	355	187	356
rect	187	355	188	356
rect	188	355	189	356
rect	189	355	190	356
rect	190	355	191	356
rect	191	355	192	356
rect	192	355	193	356
rect	193	355	194	356
rect	194	355	195	356
rect	195	355	196	356
rect	196	355	197	356
rect	197	355	198	356
rect	198	355	199	356
rect	199	355	200	356
rect	200	355	201	356
rect	201	355	202	356
rect	202	355	203	356
rect	203	355	204	356
rect	204	355	205	356
rect	205	355	206	356
rect	206	355	207	356
rect	207	355	208	356
rect	208	355	209	356
rect	209	355	210	356
rect	210	355	211	356
rect	211	355	212	356
rect	212	355	213	356
rect	213	355	214	356
rect	214	355	215	356
rect	215	355	216	356
rect	216	355	217	356
rect	217	355	218	356
rect	219	355	220	356
rect	220	355	221	356
rect	221	355	222	356
rect	222	355	223	356
rect	223	355	224	356
rect	224	355	225	356
rect	225	355	226	356
rect	226	355	227	356
rect	227	355	228	356
rect	228	355	229	356
rect	229	355	230	356
rect	230	355	231	356
rect	231	355	232	356
rect	232	355	233	356
rect	233	355	234	356
rect	234	355	235	356
rect	235	355	236	356
rect	236	355	237	356
rect	237	355	238	356
rect	238	355	239	356
rect	239	355	240	356
rect	240	355	241	356
rect	241	355	242	356
rect	242	355	243	356
rect	243	355	244	356
rect	244	355	245	356
rect	245	355	246	356
rect	246	355	247	356
rect	247	355	248	356
rect	248	355	249	356
rect	249	355	250	356
rect	250	355	251	356
rect	251	355	252	356
rect	252	355	253	356
rect	253	355	254	356
rect	254	355	255	356
rect	255	355	256	356
rect	256	355	257	356
rect	257	355	258	356
rect	258	355	259	356
rect	259	355	260	356
rect	260	355	261	356
rect	261	355	262	356
rect	262	355	263	356
rect	263	355	264	356
rect	264	355	265	356
rect	265	355	266	356
rect	266	355	267	356
rect	267	355	268	356
rect	268	355	269	356
rect	269	355	270	356
rect	270	355	271	356
rect	271	355	272	356
rect	272	355	273	356
rect	273	355	274	356
rect	274	355	275	356
rect	275	355	276	356
rect	276	355	277	356
rect	277	355	278	356
rect	278	355	279	356
rect	279	355	280	356
rect	280	355	281	356
rect	281	355	282	356
rect	282	355	283	356
rect	283	355	284	356
rect	284	355	285	356
rect	285	355	286	356
rect	286	355	287	356
rect	287	355	288	356
rect	288	355	289	356
rect	289	355	290	356
rect	290	355	291	356
rect	291	355	292	356
rect	292	355	293	356
rect	293	355	294	356
rect	294	355	295	356
rect	295	355	296	356
rect	296	355	297	356
rect	298	355	299	356
rect	299	355	300	356
rect	300	355	301	356
rect	301	355	302	356
rect	302	355	303	356
rect	303	355	304	356
rect	304	355	305	356
rect	305	355	306	356
rect	306	355	307	356
rect	307	355	308	356
rect	308	355	309	356
rect	309	355	310	356
rect	310	355	311	356
rect	311	355	312	356
rect	312	355	313	356
rect	313	355	314	356
rect	314	355	315	356
rect	315	355	316	356
rect	316	355	317	356
rect	317	355	318	356
rect	318	355	319	356
rect	319	355	320	356
rect	320	355	321	356
rect	321	355	322	356
rect	322	355	323	356
rect	323	355	324	356
rect	324	355	325	356
rect	325	355	326	356
rect	326	355	327	356
rect	327	355	328	356
rect	328	355	329	356
rect	329	355	330	356
rect	330	355	331	356
rect	332	355	333	356
rect	333	355	334	356
rect	334	355	335	356
rect	335	355	336	356
rect	336	355	337	356
rect	337	355	338	356
rect	339	355	340	356
rect	340	355	341	356
rect	341	355	342	356
rect	342	355	343	356
rect	343	355	344	356
rect	344	355	345	356
rect	345	355	346	356
rect	346	355	347	356
rect	347	355	348	356
rect	348	355	349	356
rect	349	355	350	356
rect	350	355	351	356
rect	351	355	352	356
rect	352	355	353	356
rect	353	355	354	356
rect	354	355	355	356
rect	355	355	356	356
rect	356	355	357	356
rect	357	355	358	356
rect	358	355	359	356
rect	359	355	360	356
rect	360	355	361	356
rect	361	355	362	356
rect	362	355	363	356
rect	363	355	364	356
rect	364	355	365	356
rect	365	355	366	356
rect	367	355	368	356
rect	368	355	369	356
rect	369	355	370	356
rect	370	355	371	356
rect	371	355	372	356
rect	372	355	373	356
rect	374	355	375	356
rect	375	355	376	356
rect	376	355	377	356
rect	377	355	378	356
rect	378	355	379	356
rect	379	355	380	356
rect	381	355	382	356
rect	382	355	383	356
rect	383	355	384	356
rect	384	355	385	356
rect	385	355	386	356
rect	386	355	387	356
rect	388	355	389	356
rect	389	355	390	356
rect	390	355	391	356
rect	391	355	392	356
rect	392	355	393	356
rect	393	355	394	356
rect	394	355	395	356
rect	395	355	396	356
rect	396	355	397	356
rect	0	381	1	382
rect	1	381	2	382
rect	2	381	3	382
rect	3	381	4	382
rect	4	381	5	382
rect	5	381	6	382
rect	7	381	8	382
rect	8	381	9	382
rect	9	381	10	382
rect	10	381	11	382
rect	11	381	12	382
rect	12	381	13	382
rect	13	381	14	382
rect	14	381	15	382
rect	15	381	16	382
rect	16	381	17	382
rect	17	381	18	382
rect	18	381	19	382
rect	19	381	20	382
rect	20	381	21	382
rect	21	381	22	382
rect	23	381	24	382
rect	24	381	25	382
rect	25	381	26	382
rect	26	381	27	382
rect	27	381	28	382
rect	28	381	29	382
rect	30	381	31	382
rect	31	381	32	382
rect	32	381	33	382
rect	33	381	34	382
rect	34	381	35	382
rect	35	381	36	382
rect	37	381	38	382
rect	38	381	39	382
rect	39	381	40	382
rect	40	381	41	382
rect	41	381	42	382
rect	42	381	43	382
rect	44	381	45	382
rect	45	381	46	382
rect	46	381	47	382
rect	47	381	48	382
rect	48	381	49	382
rect	49	381	50	382
rect	51	381	52	382
rect	52	381	53	382
rect	53	381	54	382
rect	54	381	55	382
rect	55	381	56	382
rect	56	381	57	382
rect	57	381	58	382
rect	58	381	59	382
rect	59	381	60	382
rect	60	381	61	382
rect	61	381	62	382
rect	62	381	63	382
rect	63	381	64	382
rect	64	381	65	382
rect	65	381	66	382
rect	66	381	67	382
rect	67	381	68	382
rect	68	381	69	382
rect	69	381	70	382
rect	70	381	71	382
rect	71	381	72	382
rect	72	381	73	382
rect	73	381	74	382
rect	74	381	75	382
rect	75	381	76	382
rect	76	381	77	382
rect	77	381	78	382
rect	78	381	79	382
rect	79	381	80	382
rect	80	381	81	382
rect	81	381	82	382
rect	82	381	83	382
rect	83	381	84	382
rect	84	381	85	382
rect	85	381	86	382
rect	86	381	87	382
rect	87	381	88	382
rect	88	381	89	382
rect	89	381	90	382
rect	90	381	91	382
rect	91	381	92	382
rect	92	381	93	382
rect	93	381	94	382
rect	94	381	95	382
rect	95	381	96	382
rect	96	381	97	382
rect	97	381	98	382
rect	98	381	99	382
rect	99	381	100	382
rect	100	381	101	382
rect	101	381	102	382
rect	102	381	103	382
rect	103	381	104	382
rect	104	381	105	382
rect	105	381	106	382
rect	106	381	107	382
rect	107	381	108	382
rect	108	381	109	382
rect	109	381	110	382
rect	110	381	111	382
rect	111	381	112	382
rect	112	381	113	382
rect	113	381	114	382
rect	114	381	115	382
rect	115	381	116	382
rect	116	381	117	382
rect	117	381	118	382
rect	118	381	119	382
rect	119	381	120	382
rect	120	381	121	382
rect	121	381	122	382
rect	122	381	123	382
rect	123	381	124	382
rect	124	381	125	382
rect	125	381	126	382
rect	126	381	127	382
rect	127	381	128	382
rect	128	381	129	382
rect	129	381	130	382
rect	130	381	131	382
rect	131	381	132	382
rect	132	381	133	382
rect	133	381	134	382
rect	134	381	135	382
rect	135	381	136	382
rect	136	381	137	382
rect	137	381	138	382
rect	138	381	139	382
rect	139	381	140	382
rect	140	381	141	382
rect	141	381	142	382
rect	142	381	143	382
rect	143	381	144	382
rect	144	381	145	382
rect	145	381	146	382
rect	146	381	147	382
rect	147	381	148	382
rect	148	381	149	382
rect	149	381	150	382
rect	150	381	151	382
rect	151	381	152	382
rect	152	381	153	382
rect	153	381	154	382
rect	154	381	155	382
rect	155	381	156	382
rect	156	381	157	382
rect	157	381	158	382
rect	158	381	159	382
rect	160	381	161	382
rect	161	381	162	382
rect	162	381	163	382
rect	163	381	164	382
rect	164	381	165	382
rect	165	381	166	382
rect	166	381	167	382
rect	167	381	168	382
rect	168	381	169	382
rect	169	381	170	382
rect	170	381	171	382
rect	171	381	172	382
rect	172	381	173	382
rect	173	381	174	382
rect	174	381	175	382
rect	176	381	177	382
rect	177	381	178	382
rect	178	381	179	382
rect	179	381	180	382
rect	180	381	181	382
rect	181	381	182	382
rect	182	381	183	382
rect	183	381	184	382
rect	184	381	185	382
rect	185	381	186	382
rect	186	381	187	382
rect	187	381	188	382
rect	188	381	189	382
rect	189	381	190	382
rect	190	381	191	382
rect	191	381	192	382
rect	192	381	193	382
rect	193	381	194	382
rect	194	381	195	382
rect	195	381	196	382
rect	196	381	197	382
rect	197	381	198	382
rect	198	381	199	382
rect	199	381	200	382
rect	200	381	201	382
rect	201	381	202	382
rect	202	381	203	382
rect	203	381	204	382
rect	204	381	205	382
rect	205	381	206	382
rect	206	381	207	382
rect	207	381	208	382
rect	208	381	209	382
rect	210	381	211	382
rect	211	381	212	382
rect	212	381	213	382
rect	213	381	214	382
rect	214	381	215	382
rect	215	381	216	382
rect	216	381	217	382
rect	217	381	218	382
rect	218	381	219	382
rect	219	381	220	382
rect	220	381	221	382
rect	221	381	222	382
rect	222	381	223	382
rect	223	381	224	382
rect	224	381	225	382
rect	225	381	226	382
rect	226	381	227	382
rect	227	381	228	382
rect	228	381	229	382
rect	229	381	230	382
rect	230	381	231	382
rect	231	381	232	382
rect	232	381	233	382
rect	233	381	234	382
rect	234	381	235	382
rect	235	381	236	382
rect	236	381	237	382
rect	237	381	238	382
rect	238	381	239	382
rect	239	381	240	382
rect	240	381	241	382
rect	241	381	242	382
rect	242	381	243	382
rect	243	381	244	382
rect	244	381	245	382
rect	245	381	246	382
rect	246	381	247	382
rect	247	381	248	382
rect	248	381	249	382
rect	249	381	250	382
rect	250	381	251	382
rect	251	381	252	382
rect	252	381	253	382
rect	253	381	254	382
rect	254	381	255	382
rect	255	381	256	382
rect	256	381	257	382
rect	257	381	258	382
rect	258	381	259	382
rect	259	381	260	382
rect	260	381	261	382
rect	261	381	262	382
rect	262	381	263	382
rect	263	381	264	382
rect	264	381	265	382
rect	265	381	266	382
rect	266	381	267	382
rect	267	381	268	382
rect	268	381	269	382
rect	269	381	270	382
rect	270	381	271	382
rect	271	381	272	382
rect	272	381	273	382
rect	273	381	274	382
rect	274	381	275	382
rect	275	381	276	382
rect	276	381	277	382
rect	277	381	278	382
rect	278	381	279	382
rect	279	381	280	382
rect	280	381	281	382
rect	281	381	282	382
rect	282	381	283	382
rect	283	381	284	382
rect	284	381	285	382
rect	285	381	286	382
rect	286	381	287	382
rect	287	381	288	382
rect	288	381	289	382
rect	289	381	290	382
rect	290	381	291	382
rect	291	381	292	382
rect	292	381	293	382
rect	293	381	294	382
rect	294	381	295	382
rect	295	381	296	382
rect	296	381	297	382
rect	297	381	298	382
rect	298	381	299	382
rect	299	381	300	382
rect	300	381	301	382
rect	301	381	302	382
rect	302	381	303	382
rect	304	381	305	382
rect	305	381	306	382
rect	306	381	307	382
rect	307	381	308	382
rect	308	381	309	382
rect	309	381	310	382
rect	310	381	311	382
rect	311	381	312	382
rect	312	381	313	382
rect	313	381	314	382
rect	314	381	315	382
rect	315	381	316	382
rect	316	381	317	382
rect	317	381	318	382
rect	318	381	319	382
rect	319	381	320	382
rect	320	381	321	382
rect	321	381	322	382
rect	322	381	323	382
rect	323	381	324	382
rect	324	381	325	382
rect	325	381	326	382
rect	326	381	327	382
rect	327	381	328	382
rect	328	381	329	382
rect	329	381	330	382
rect	330	381	331	382
rect	331	381	332	382
rect	332	381	333	382
rect	333	381	334	382
rect	334	381	335	382
rect	335	381	336	382
rect	336	381	337	382
rect	337	381	338	382
rect	338	381	339	382
rect	339	381	340	382
rect	341	381	342	382
rect	342	381	343	382
rect	343	381	344	382
rect	344	381	345	382
rect	345	381	346	382
rect	346	381	347	382
rect	347	381	348	382
rect	348	381	349	382
rect	349	381	350	382
rect	350	381	351	382
rect	351	381	352	382
rect	352	381	353	382
rect	353	381	354	382
rect	354	381	355	382
rect	355	381	356	382
rect	357	381	358	382
rect	358	381	359	382
rect	359	381	360	382
rect	360	381	361	382
rect	361	381	362	382
rect	362	381	363	382
rect	363	381	364	382
rect	364	381	365	382
rect	365	381	366	382
rect	0	382	1	383
rect	1	382	2	383
rect	2	382	3	383
rect	3	382	4	383
rect	4	382	5	383
rect	5	382	6	383
rect	7	382	8	383
rect	8	382	9	383
rect	9	382	10	383
rect	10	382	11	383
rect	11	382	12	383
rect	12	382	13	383
rect	13	382	14	383
rect	14	382	15	383
rect	15	382	16	383
rect	16	382	17	383
rect	17	382	18	383
rect	18	382	19	383
rect	19	382	20	383
rect	20	382	21	383
rect	21	382	22	383
rect	23	382	24	383
rect	24	382	25	383
rect	25	382	26	383
rect	26	382	27	383
rect	27	382	28	383
rect	28	382	29	383
rect	30	382	31	383
rect	31	382	32	383
rect	32	382	33	383
rect	33	382	34	383
rect	34	382	35	383
rect	35	382	36	383
rect	37	382	38	383
rect	38	382	39	383
rect	39	382	40	383
rect	40	382	41	383
rect	41	382	42	383
rect	42	382	43	383
rect	44	382	45	383
rect	45	382	46	383
rect	46	382	47	383
rect	47	382	48	383
rect	48	382	49	383
rect	49	382	50	383
rect	51	382	52	383
rect	52	382	53	383
rect	53	382	54	383
rect	54	382	55	383
rect	55	382	56	383
rect	56	382	57	383
rect	57	382	58	383
rect	58	382	59	383
rect	59	382	60	383
rect	60	382	61	383
rect	61	382	62	383
rect	62	382	63	383
rect	63	382	64	383
rect	64	382	65	383
rect	65	382	66	383
rect	66	382	67	383
rect	67	382	68	383
rect	68	382	69	383
rect	69	382	70	383
rect	70	382	71	383
rect	71	382	72	383
rect	72	382	73	383
rect	73	382	74	383
rect	74	382	75	383
rect	75	382	76	383
rect	76	382	77	383
rect	77	382	78	383
rect	78	382	79	383
rect	79	382	80	383
rect	80	382	81	383
rect	81	382	82	383
rect	82	382	83	383
rect	83	382	84	383
rect	84	382	85	383
rect	85	382	86	383
rect	86	382	87	383
rect	87	382	88	383
rect	88	382	89	383
rect	89	382	90	383
rect	90	382	91	383
rect	91	382	92	383
rect	92	382	93	383
rect	93	382	94	383
rect	94	382	95	383
rect	95	382	96	383
rect	96	382	97	383
rect	97	382	98	383
rect	98	382	99	383
rect	99	382	100	383
rect	100	382	101	383
rect	101	382	102	383
rect	102	382	103	383
rect	103	382	104	383
rect	104	382	105	383
rect	105	382	106	383
rect	106	382	107	383
rect	107	382	108	383
rect	108	382	109	383
rect	109	382	110	383
rect	110	382	111	383
rect	111	382	112	383
rect	112	382	113	383
rect	113	382	114	383
rect	114	382	115	383
rect	115	382	116	383
rect	116	382	117	383
rect	117	382	118	383
rect	118	382	119	383
rect	119	382	120	383
rect	120	382	121	383
rect	121	382	122	383
rect	122	382	123	383
rect	123	382	124	383
rect	124	382	125	383
rect	125	382	126	383
rect	126	382	127	383
rect	127	382	128	383
rect	128	382	129	383
rect	129	382	130	383
rect	130	382	131	383
rect	131	382	132	383
rect	132	382	133	383
rect	133	382	134	383
rect	134	382	135	383
rect	135	382	136	383
rect	136	382	137	383
rect	137	382	138	383
rect	138	382	139	383
rect	139	382	140	383
rect	140	382	141	383
rect	141	382	142	383
rect	142	382	143	383
rect	143	382	144	383
rect	144	382	145	383
rect	145	382	146	383
rect	146	382	147	383
rect	147	382	148	383
rect	148	382	149	383
rect	149	382	150	383
rect	150	382	151	383
rect	151	382	152	383
rect	152	382	153	383
rect	153	382	154	383
rect	154	382	155	383
rect	155	382	156	383
rect	156	382	157	383
rect	157	382	158	383
rect	158	382	159	383
rect	160	382	161	383
rect	161	382	162	383
rect	162	382	163	383
rect	163	382	164	383
rect	164	382	165	383
rect	165	382	166	383
rect	166	382	167	383
rect	167	382	168	383
rect	168	382	169	383
rect	169	382	170	383
rect	170	382	171	383
rect	171	382	172	383
rect	172	382	173	383
rect	173	382	174	383
rect	174	382	175	383
rect	176	382	177	383
rect	177	382	178	383
rect	178	382	179	383
rect	179	382	180	383
rect	180	382	181	383
rect	181	382	182	383
rect	182	382	183	383
rect	183	382	184	383
rect	184	382	185	383
rect	185	382	186	383
rect	186	382	187	383
rect	187	382	188	383
rect	188	382	189	383
rect	189	382	190	383
rect	190	382	191	383
rect	191	382	192	383
rect	192	382	193	383
rect	193	382	194	383
rect	194	382	195	383
rect	195	382	196	383
rect	196	382	197	383
rect	197	382	198	383
rect	198	382	199	383
rect	199	382	200	383
rect	200	382	201	383
rect	201	382	202	383
rect	202	382	203	383
rect	203	382	204	383
rect	204	382	205	383
rect	205	382	206	383
rect	206	382	207	383
rect	207	382	208	383
rect	208	382	209	383
rect	210	382	211	383
rect	211	382	212	383
rect	212	382	213	383
rect	213	382	214	383
rect	214	382	215	383
rect	215	382	216	383
rect	216	382	217	383
rect	217	382	218	383
rect	218	382	219	383
rect	219	382	220	383
rect	220	382	221	383
rect	221	382	222	383
rect	222	382	223	383
rect	223	382	224	383
rect	224	382	225	383
rect	225	382	226	383
rect	226	382	227	383
rect	227	382	228	383
rect	228	382	229	383
rect	229	382	230	383
rect	230	382	231	383
rect	231	382	232	383
rect	232	382	233	383
rect	233	382	234	383
rect	234	382	235	383
rect	235	382	236	383
rect	236	382	237	383
rect	237	382	238	383
rect	238	382	239	383
rect	239	382	240	383
rect	240	382	241	383
rect	241	382	242	383
rect	242	382	243	383
rect	243	382	244	383
rect	244	382	245	383
rect	245	382	246	383
rect	246	382	247	383
rect	247	382	248	383
rect	248	382	249	383
rect	249	382	250	383
rect	250	382	251	383
rect	251	382	252	383
rect	252	382	253	383
rect	253	382	254	383
rect	254	382	255	383
rect	255	382	256	383
rect	256	382	257	383
rect	257	382	258	383
rect	258	382	259	383
rect	259	382	260	383
rect	260	382	261	383
rect	261	382	262	383
rect	262	382	263	383
rect	263	382	264	383
rect	264	382	265	383
rect	265	382	266	383
rect	266	382	267	383
rect	267	382	268	383
rect	268	382	269	383
rect	269	382	270	383
rect	270	382	271	383
rect	271	382	272	383
rect	272	382	273	383
rect	273	382	274	383
rect	274	382	275	383
rect	275	382	276	383
rect	276	382	277	383
rect	277	382	278	383
rect	278	382	279	383
rect	279	382	280	383
rect	280	382	281	383
rect	281	382	282	383
rect	282	382	283	383
rect	283	382	284	383
rect	284	382	285	383
rect	285	382	286	383
rect	286	382	287	383
rect	287	382	288	383
rect	288	382	289	383
rect	289	382	290	383
rect	290	382	291	383
rect	291	382	292	383
rect	292	382	293	383
rect	293	382	294	383
rect	294	382	295	383
rect	295	382	296	383
rect	296	382	297	383
rect	297	382	298	383
rect	298	382	299	383
rect	299	382	300	383
rect	300	382	301	383
rect	301	382	302	383
rect	302	382	303	383
rect	304	382	305	383
rect	305	382	306	383
rect	306	382	307	383
rect	307	382	308	383
rect	308	382	309	383
rect	309	382	310	383
rect	310	382	311	383
rect	311	382	312	383
rect	312	382	313	383
rect	313	382	314	383
rect	314	382	315	383
rect	315	382	316	383
rect	316	382	317	383
rect	317	382	318	383
rect	318	382	319	383
rect	319	382	320	383
rect	320	382	321	383
rect	321	382	322	383
rect	322	382	323	383
rect	323	382	324	383
rect	324	382	325	383
rect	325	382	326	383
rect	326	382	327	383
rect	327	382	328	383
rect	328	382	329	383
rect	329	382	330	383
rect	330	382	331	383
rect	331	382	332	383
rect	332	382	333	383
rect	333	382	334	383
rect	334	382	335	383
rect	335	382	336	383
rect	336	382	337	383
rect	337	382	338	383
rect	338	382	339	383
rect	339	382	340	383
rect	341	382	342	383
rect	342	382	343	383
rect	343	382	344	383
rect	344	382	345	383
rect	345	382	346	383
rect	346	382	347	383
rect	347	382	348	383
rect	348	382	349	383
rect	349	382	350	383
rect	350	382	351	383
rect	351	382	352	383
rect	352	382	353	383
rect	353	382	354	383
rect	354	382	355	383
rect	355	382	356	383
rect	357	382	358	383
rect	358	382	359	383
rect	359	382	360	383
rect	360	382	361	383
rect	361	382	362	383
rect	362	382	363	383
rect	363	382	364	383
rect	364	382	365	383
rect	365	382	366	383
rect	0	383	1	384
rect	1	383	2	384
rect	2	383	3	384
rect	3	383	4	384
rect	4	383	5	384
rect	5	383	6	384
rect	7	383	8	384
rect	8	383	9	384
rect	9	383	10	384
rect	10	383	11	384
rect	11	383	12	384
rect	12	383	13	384
rect	13	383	14	384
rect	14	383	15	384
rect	15	383	16	384
rect	16	383	17	384
rect	17	383	18	384
rect	18	383	19	384
rect	19	383	20	384
rect	20	383	21	384
rect	21	383	22	384
rect	23	383	24	384
rect	24	383	25	384
rect	25	383	26	384
rect	26	383	27	384
rect	27	383	28	384
rect	28	383	29	384
rect	30	383	31	384
rect	31	383	32	384
rect	32	383	33	384
rect	33	383	34	384
rect	34	383	35	384
rect	35	383	36	384
rect	37	383	38	384
rect	38	383	39	384
rect	39	383	40	384
rect	40	383	41	384
rect	41	383	42	384
rect	42	383	43	384
rect	44	383	45	384
rect	45	383	46	384
rect	46	383	47	384
rect	47	383	48	384
rect	48	383	49	384
rect	49	383	50	384
rect	51	383	52	384
rect	52	383	53	384
rect	53	383	54	384
rect	54	383	55	384
rect	55	383	56	384
rect	56	383	57	384
rect	57	383	58	384
rect	58	383	59	384
rect	59	383	60	384
rect	60	383	61	384
rect	61	383	62	384
rect	62	383	63	384
rect	63	383	64	384
rect	64	383	65	384
rect	65	383	66	384
rect	66	383	67	384
rect	67	383	68	384
rect	68	383	69	384
rect	69	383	70	384
rect	70	383	71	384
rect	71	383	72	384
rect	72	383	73	384
rect	73	383	74	384
rect	74	383	75	384
rect	75	383	76	384
rect	76	383	77	384
rect	77	383	78	384
rect	78	383	79	384
rect	79	383	80	384
rect	80	383	81	384
rect	81	383	82	384
rect	82	383	83	384
rect	83	383	84	384
rect	84	383	85	384
rect	85	383	86	384
rect	86	383	87	384
rect	87	383	88	384
rect	88	383	89	384
rect	89	383	90	384
rect	90	383	91	384
rect	91	383	92	384
rect	92	383	93	384
rect	93	383	94	384
rect	94	383	95	384
rect	95	383	96	384
rect	96	383	97	384
rect	97	383	98	384
rect	98	383	99	384
rect	99	383	100	384
rect	100	383	101	384
rect	101	383	102	384
rect	102	383	103	384
rect	103	383	104	384
rect	104	383	105	384
rect	105	383	106	384
rect	106	383	107	384
rect	107	383	108	384
rect	108	383	109	384
rect	109	383	110	384
rect	110	383	111	384
rect	111	383	112	384
rect	112	383	113	384
rect	113	383	114	384
rect	114	383	115	384
rect	115	383	116	384
rect	116	383	117	384
rect	117	383	118	384
rect	118	383	119	384
rect	119	383	120	384
rect	120	383	121	384
rect	121	383	122	384
rect	122	383	123	384
rect	123	383	124	384
rect	124	383	125	384
rect	125	383	126	384
rect	126	383	127	384
rect	127	383	128	384
rect	128	383	129	384
rect	129	383	130	384
rect	130	383	131	384
rect	131	383	132	384
rect	132	383	133	384
rect	133	383	134	384
rect	134	383	135	384
rect	135	383	136	384
rect	136	383	137	384
rect	137	383	138	384
rect	138	383	139	384
rect	139	383	140	384
rect	140	383	141	384
rect	141	383	142	384
rect	142	383	143	384
rect	143	383	144	384
rect	144	383	145	384
rect	145	383	146	384
rect	146	383	147	384
rect	147	383	148	384
rect	148	383	149	384
rect	149	383	150	384
rect	150	383	151	384
rect	151	383	152	384
rect	152	383	153	384
rect	153	383	154	384
rect	154	383	155	384
rect	155	383	156	384
rect	156	383	157	384
rect	157	383	158	384
rect	158	383	159	384
rect	160	383	161	384
rect	161	383	162	384
rect	162	383	163	384
rect	163	383	164	384
rect	164	383	165	384
rect	165	383	166	384
rect	166	383	167	384
rect	167	383	168	384
rect	168	383	169	384
rect	169	383	170	384
rect	170	383	171	384
rect	171	383	172	384
rect	172	383	173	384
rect	173	383	174	384
rect	174	383	175	384
rect	176	383	177	384
rect	177	383	178	384
rect	178	383	179	384
rect	179	383	180	384
rect	180	383	181	384
rect	181	383	182	384
rect	182	383	183	384
rect	183	383	184	384
rect	184	383	185	384
rect	185	383	186	384
rect	186	383	187	384
rect	187	383	188	384
rect	188	383	189	384
rect	189	383	190	384
rect	190	383	191	384
rect	191	383	192	384
rect	192	383	193	384
rect	193	383	194	384
rect	194	383	195	384
rect	195	383	196	384
rect	196	383	197	384
rect	197	383	198	384
rect	198	383	199	384
rect	199	383	200	384
rect	200	383	201	384
rect	201	383	202	384
rect	202	383	203	384
rect	203	383	204	384
rect	204	383	205	384
rect	205	383	206	384
rect	206	383	207	384
rect	207	383	208	384
rect	208	383	209	384
rect	210	383	211	384
rect	211	383	212	384
rect	212	383	213	384
rect	213	383	214	384
rect	214	383	215	384
rect	215	383	216	384
rect	216	383	217	384
rect	217	383	218	384
rect	218	383	219	384
rect	219	383	220	384
rect	220	383	221	384
rect	221	383	222	384
rect	222	383	223	384
rect	223	383	224	384
rect	224	383	225	384
rect	225	383	226	384
rect	226	383	227	384
rect	227	383	228	384
rect	228	383	229	384
rect	229	383	230	384
rect	230	383	231	384
rect	231	383	232	384
rect	232	383	233	384
rect	233	383	234	384
rect	234	383	235	384
rect	235	383	236	384
rect	236	383	237	384
rect	237	383	238	384
rect	238	383	239	384
rect	239	383	240	384
rect	240	383	241	384
rect	241	383	242	384
rect	242	383	243	384
rect	243	383	244	384
rect	244	383	245	384
rect	245	383	246	384
rect	246	383	247	384
rect	247	383	248	384
rect	248	383	249	384
rect	249	383	250	384
rect	250	383	251	384
rect	251	383	252	384
rect	252	383	253	384
rect	253	383	254	384
rect	254	383	255	384
rect	255	383	256	384
rect	256	383	257	384
rect	257	383	258	384
rect	258	383	259	384
rect	259	383	260	384
rect	260	383	261	384
rect	261	383	262	384
rect	262	383	263	384
rect	263	383	264	384
rect	264	383	265	384
rect	265	383	266	384
rect	266	383	267	384
rect	267	383	268	384
rect	268	383	269	384
rect	269	383	270	384
rect	270	383	271	384
rect	271	383	272	384
rect	272	383	273	384
rect	273	383	274	384
rect	274	383	275	384
rect	275	383	276	384
rect	276	383	277	384
rect	277	383	278	384
rect	278	383	279	384
rect	279	383	280	384
rect	280	383	281	384
rect	281	383	282	384
rect	282	383	283	384
rect	283	383	284	384
rect	284	383	285	384
rect	285	383	286	384
rect	286	383	287	384
rect	287	383	288	384
rect	288	383	289	384
rect	289	383	290	384
rect	290	383	291	384
rect	291	383	292	384
rect	292	383	293	384
rect	293	383	294	384
rect	294	383	295	384
rect	295	383	296	384
rect	296	383	297	384
rect	297	383	298	384
rect	298	383	299	384
rect	299	383	300	384
rect	300	383	301	384
rect	301	383	302	384
rect	302	383	303	384
rect	304	383	305	384
rect	305	383	306	384
rect	306	383	307	384
rect	307	383	308	384
rect	308	383	309	384
rect	309	383	310	384
rect	310	383	311	384
rect	311	383	312	384
rect	312	383	313	384
rect	313	383	314	384
rect	314	383	315	384
rect	315	383	316	384
rect	316	383	317	384
rect	317	383	318	384
rect	318	383	319	384
rect	319	383	320	384
rect	320	383	321	384
rect	321	383	322	384
rect	322	383	323	384
rect	323	383	324	384
rect	324	383	325	384
rect	325	383	326	384
rect	326	383	327	384
rect	327	383	328	384
rect	328	383	329	384
rect	329	383	330	384
rect	330	383	331	384
rect	331	383	332	384
rect	332	383	333	384
rect	333	383	334	384
rect	334	383	335	384
rect	335	383	336	384
rect	336	383	337	384
rect	337	383	338	384
rect	338	383	339	384
rect	339	383	340	384
rect	341	383	342	384
rect	342	383	343	384
rect	343	383	344	384
rect	344	383	345	384
rect	345	383	346	384
rect	346	383	347	384
rect	347	383	348	384
rect	348	383	349	384
rect	349	383	350	384
rect	350	383	351	384
rect	351	383	352	384
rect	352	383	353	384
rect	353	383	354	384
rect	354	383	355	384
rect	355	383	356	384
rect	357	383	358	384
rect	358	383	359	384
rect	359	383	360	384
rect	360	383	361	384
rect	361	383	362	384
rect	362	383	363	384
rect	363	383	364	384
rect	364	383	365	384
rect	365	383	366	384
rect	0	384	1	385
rect	1	384	2	385
rect	2	384	3	385
rect	3	384	4	385
rect	4	384	5	385
rect	5	384	6	385
rect	7	384	8	385
rect	8	384	9	385
rect	9	384	10	385
rect	10	384	11	385
rect	11	384	12	385
rect	12	384	13	385
rect	13	384	14	385
rect	14	384	15	385
rect	15	384	16	385
rect	16	384	17	385
rect	17	384	18	385
rect	18	384	19	385
rect	19	384	20	385
rect	20	384	21	385
rect	21	384	22	385
rect	23	384	24	385
rect	24	384	25	385
rect	25	384	26	385
rect	26	384	27	385
rect	27	384	28	385
rect	28	384	29	385
rect	30	384	31	385
rect	31	384	32	385
rect	32	384	33	385
rect	33	384	34	385
rect	34	384	35	385
rect	35	384	36	385
rect	37	384	38	385
rect	38	384	39	385
rect	39	384	40	385
rect	40	384	41	385
rect	41	384	42	385
rect	42	384	43	385
rect	44	384	45	385
rect	45	384	46	385
rect	46	384	47	385
rect	47	384	48	385
rect	48	384	49	385
rect	49	384	50	385
rect	51	384	52	385
rect	52	384	53	385
rect	53	384	54	385
rect	54	384	55	385
rect	55	384	56	385
rect	56	384	57	385
rect	57	384	58	385
rect	58	384	59	385
rect	59	384	60	385
rect	60	384	61	385
rect	61	384	62	385
rect	62	384	63	385
rect	63	384	64	385
rect	64	384	65	385
rect	65	384	66	385
rect	66	384	67	385
rect	67	384	68	385
rect	68	384	69	385
rect	69	384	70	385
rect	70	384	71	385
rect	71	384	72	385
rect	72	384	73	385
rect	73	384	74	385
rect	74	384	75	385
rect	75	384	76	385
rect	76	384	77	385
rect	77	384	78	385
rect	78	384	79	385
rect	79	384	80	385
rect	80	384	81	385
rect	81	384	82	385
rect	82	384	83	385
rect	83	384	84	385
rect	84	384	85	385
rect	85	384	86	385
rect	86	384	87	385
rect	87	384	88	385
rect	88	384	89	385
rect	89	384	90	385
rect	90	384	91	385
rect	91	384	92	385
rect	92	384	93	385
rect	93	384	94	385
rect	94	384	95	385
rect	95	384	96	385
rect	96	384	97	385
rect	97	384	98	385
rect	98	384	99	385
rect	99	384	100	385
rect	100	384	101	385
rect	101	384	102	385
rect	102	384	103	385
rect	103	384	104	385
rect	104	384	105	385
rect	105	384	106	385
rect	106	384	107	385
rect	107	384	108	385
rect	108	384	109	385
rect	109	384	110	385
rect	110	384	111	385
rect	111	384	112	385
rect	112	384	113	385
rect	113	384	114	385
rect	114	384	115	385
rect	115	384	116	385
rect	116	384	117	385
rect	117	384	118	385
rect	118	384	119	385
rect	119	384	120	385
rect	120	384	121	385
rect	121	384	122	385
rect	122	384	123	385
rect	123	384	124	385
rect	124	384	125	385
rect	125	384	126	385
rect	126	384	127	385
rect	127	384	128	385
rect	128	384	129	385
rect	129	384	130	385
rect	130	384	131	385
rect	131	384	132	385
rect	132	384	133	385
rect	133	384	134	385
rect	134	384	135	385
rect	135	384	136	385
rect	136	384	137	385
rect	137	384	138	385
rect	138	384	139	385
rect	139	384	140	385
rect	140	384	141	385
rect	141	384	142	385
rect	142	384	143	385
rect	143	384	144	385
rect	144	384	145	385
rect	145	384	146	385
rect	146	384	147	385
rect	147	384	148	385
rect	148	384	149	385
rect	149	384	150	385
rect	150	384	151	385
rect	151	384	152	385
rect	152	384	153	385
rect	153	384	154	385
rect	154	384	155	385
rect	155	384	156	385
rect	156	384	157	385
rect	157	384	158	385
rect	158	384	159	385
rect	160	384	161	385
rect	161	384	162	385
rect	162	384	163	385
rect	163	384	164	385
rect	164	384	165	385
rect	165	384	166	385
rect	166	384	167	385
rect	167	384	168	385
rect	168	384	169	385
rect	169	384	170	385
rect	170	384	171	385
rect	171	384	172	385
rect	172	384	173	385
rect	173	384	174	385
rect	174	384	175	385
rect	176	384	177	385
rect	177	384	178	385
rect	178	384	179	385
rect	179	384	180	385
rect	180	384	181	385
rect	181	384	182	385
rect	182	384	183	385
rect	183	384	184	385
rect	184	384	185	385
rect	185	384	186	385
rect	186	384	187	385
rect	187	384	188	385
rect	188	384	189	385
rect	189	384	190	385
rect	190	384	191	385
rect	191	384	192	385
rect	192	384	193	385
rect	193	384	194	385
rect	194	384	195	385
rect	195	384	196	385
rect	196	384	197	385
rect	197	384	198	385
rect	198	384	199	385
rect	199	384	200	385
rect	200	384	201	385
rect	201	384	202	385
rect	202	384	203	385
rect	203	384	204	385
rect	204	384	205	385
rect	205	384	206	385
rect	206	384	207	385
rect	207	384	208	385
rect	208	384	209	385
rect	210	384	211	385
rect	211	384	212	385
rect	212	384	213	385
rect	213	384	214	385
rect	214	384	215	385
rect	215	384	216	385
rect	216	384	217	385
rect	217	384	218	385
rect	218	384	219	385
rect	219	384	220	385
rect	220	384	221	385
rect	221	384	222	385
rect	222	384	223	385
rect	223	384	224	385
rect	224	384	225	385
rect	225	384	226	385
rect	226	384	227	385
rect	227	384	228	385
rect	228	384	229	385
rect	229	384	230	385
rect	230	384	231	385
rect	231	384	232	385
rect	232	384	233	385
rect	233	384	234	385
rect	234	384	235	385
rect	235	384	236	385
rect	236	384	237	385
rect	237	384	238	385
rect	238	384	239	385
rect	239	384	240	385
rect	240	384	241	385
rect	241	384	242	385
rect	242	384	243	385
rect	243	384	244	385
rect	244	384	245	385
rect	245	384	246	385
rect	246	384	247	385
rect	247	384	248	385
rect	248	384	249	385
rect	249	384	250	385
rect	250	384	251	385
rect	251	384	252	385
rect	252	384	253	385
rect	253	384	254	385
rect	254	384	255	385
rect	255	384	256	385
rect	256	384	257	385
rect	257	384	258	385
rect	258	384	259	385
rect	259	384	260	385
rect	260	384	261	385
rect	261	384	262	385
rect	262	384	263	385
rect	263	384	264	385
rect	264	384	265	385
rect	265	384	266	385
rect	266	384	267	385
rect	267	384	268	385
rect	268	384	269	385
rect	269	384	270	385
rect	270	384	271	385
rect	271	384	272	385
rect	272	384	273	385
rect	273	384	274	385
rect	274	384	275	385
rect	275	384	276	385
rect	276	384	277	385
rect	277	384	278	385
rect	278	384	279	385
rect	279	384	280	385
rect	280	384	281	385
rect	281	384	282	385
rect	282	384	283	385
rect	283	384	284	385
rect	284	384	285	385
rect	285	384	286	385
rect	286	384	287	385
rect	287	384	288	385
rect	288	384	289	385
rect	289	384	290	385
rect	290	384	291	385
rect	291	384	292	385
rect	292	384	293	385
rect	293	384	294	385
rect	294	384	295	385
rect	295	384	296	385
rect	296	384	297	385
rect	297	384	298	385
rect	298	384	299	385
rect	299	384	300	385
rect	300	384	301	385
rect	301	384	302	385
rect	302	384	303	385
rect	304	384	305	385
rect	305	384	306	385
rect	306	384	307	385
rect	307	384	308	385
rect	308	384	309	385
rect	309	384	310	385
rect	310	384	311	385
rect	311	384	312	385
rect	312	384	313	385
rect	313	384	314	385
rect	314	384	315	385
rect	315	384	316	385
rect	316	384	317	385
rect	317	384	318	385
rect	318	384	319	385
rect	319	384	320	385
rect	320	384	321	385
rect	321	384	322	385
rect	322	384	323	385
rect	323	384	324	385
rect	324	384	325	385
rect	325	384	326	385
rect	326	384	327	385
rect	327	384	328	385
rect	328	384	329	385
rect	329	384	330	385
rect	330	384	331	385
rect	331	384	332	385
rect	332	384	333	385
rect	333	384	334	385
rect	334	384	335	385
rect	335	384	336	385
rect	336	384	337	385
rect	337	384	338	385
rect	338	384	339	385
rect	339	384	340	385
rect	341	384	342	385
rect	342	384	343	385
rect	343	384	344	385
rect	344	384	345	385
rect	345	384	346	385
rect	346	384	347	385
rect	347	384	348	385
rect	348	384	349	385
rect	349	384	350	385
rect	350	384	351	385
rect	351	384	352	385
rect	352	384	353	385
rect	353	384	354	385
rect	354	384	355	385
rect	355	384	356	385
rect	357	384	358	385
rect	358	384	359	385
rect	359	384	360	385
rect	360	384	361	385
rect	361	384	362	385
rect	362	384	363	385
rect	363	384	364	385
rect	364	384	365	385
rect	365	384	366	385
rect	0	385	1	386
rect	1	385	2	386
rect	2	385	3	386
rect	3	385	4	386
rect	4	385	5	386
rect	5	385	6	386
rect	7	385	8	386
rect	8	385	9	386
rect	9	385	10	386
rect	10	385	11	386
rect	11	385	12	386
rect	12	385	13	386
rect	13	385	14	386
rect	14	385	15	386
rect	15	385	16	386
rect	16	385	17	386
rect	17	385	18	386
rect	18	385	19	386
rect	19	385	20	386
rect	20	385	21	386
rect	21	385	22	386
rect	23	385	24	386
rect	24	385	25	386
rect	25	385	26	386
rect	26	385	27	386
rect	27	385	28	386
rect	28	385	29	386
rect	30	385	31	386
rect	31	385	32	386
rect	32	385	33	386
rect	33	385	34	386
rect	34	385	35	386
rect	35	385	36	386
rect	37	385	38	386
rect	38	385	39	386
rect	39	385	40	386
rect	40	385	41	386
rect	41	385	42	386
rect	42	385	43	386
rect	44	385	45	386
rect	45	385	46	386
rect	46	385	47	386
rect	47	385	48	386
rect	48	385	49	386
rect	49	385	50	386
rect	51	385	52	386
rect	52	385	53	386
rect	53	385	54	386
rect	54	385	55	386
rect	55	385	56	386
rect	56	385	57	386
rect	57	385	58	386
rect	58	385	59	386
rect	59	385	60	386
rect	60	385	61	386
rect	61	385	62	386
rect	62	385	63	386
rect	63	385	64	386
rect	64	385	65	386
rect	65	385	66	386
rect	66	385	67	386
rect	67	385	68	386
rect	68	385	69	386
rect	69	385	70	386
rect	70	385	71	386
rect	71	385	72	386
rect	72	385	73	386
rect	73	385	74	386
rect	74	385	75	386
rect	75	385	76	386
rect	76	385	77	386
rect	77	385	78	386
rect	78	385	79	386
rect	79	385	80	386
rect	80	385	81	386
rect	81	385	82	386
rect	82	385	83	386
rect	83	385	84	386
rect	84	385	85	386
rect	85	385	86	386
rect	86	385	87	386
rect	87	385	88	386
rect	88	385	89	386
rect	89	385	90	386
rect	90	385	91	386
rect	91	385	92	386
rect	92	385	93	386
rect	93	385	94	386
rect	94	385	95	386
rect	95	385	96	386
rect	96	385	97	386
rect	97	385	98	386
rect	98	385	99	386
rect	99	385	100	386
rect	100	385	101	386
rect	101	385	102	386
rect	102	385	103	386
rect	103	385	104	386
rect	104	385	105	386
rect	105	385	106	386
rect	106	385	107	386
rect	107	385	108	386
rect	108	385	109	386
rect	109	385	110	386
rect	110	385	111	386
rect	111	385	112	386
rect	112	385	113	386
rect	113	385	114	386
rect	114	385	115	386
rect	115	385	116	386
rect	116	385	117	386
rect	117	385	118	386
rect	118	385	119	386
rect	119	385	120	386
rect	120	385	121	386
rect	121	385	122	386
rect	122	385	123	386
rect	123	385	124	386
rect	124	385	125	386
rect	125	385	126	386
rect	126	385	127	386
rect	127	385	128	386
rect	128	385	129	386
rect	129	385	130	386
rect	130	385	131	386
rect	131	385	132	386
rect	132	385	133	386
rect	133	385	134	386
rect	134	385	135	386
rect	135	385	136	386
rect	136	385	137	386
rect	137	385	138	386
rect	138	385	139	386
rect	139	385	140	386
rect	140	385	141	386
rect	141	385	142	386
rect	142	385	143	386
rect	143	385	144	386
rect	144	385	145	386
rect	145	385	146	386
rect	146	385	147	386
rect	147	385	148	386
rect	148	385	149	386
rect	149	385	150	386
rect	150	385	151	386
rect	151	385	152	386
rect	152	385	153	386
rect	153	385	154	386
rect	154	385	155	386
rect	155	385	156	386
rect	156	385	157	386
rect	157	385	158	386
rect	158	385	159	386
rect	160	385	161	386
rect	161	385	162	386
rect	162	385	163	386
rect	163	385	164	386
rect	164	385	165	386
rect	165	385	166	386
rect	166	385	167	386
rect	167	385	168	386
rect	168	385	169	386
rect	169	385	170	386
rect	170	385	171	386
rect	171	385	172	386
rect	172	385	173	386
rect	173	385	174	386
rect	174	385	175	386
rect	176	385	177	386
rect	177	385	178	386
rect	178	385	179	386
rect	179	385	180	386
rect	180	385	181	386
rect	181	385	182	386
rect	182	385	183	386
rect	183	385	184	386
rect	184	385	185	386
rect	185	385	186	386
rect	186	385	187	386
rect	187	385	188	386
rect	188	385	189	386
rect	189	385	190	386
rect	190	385	191	386
rect	191	385	192	386
rect	192	385	193	386
rect	193	385	194	386
rect	194	385	195	386
rect	195	385	196	386
rect	196	385	197	386
rect	197	385	198	386
rect	198	385	199	386
rect	199	385	200	386
rect	200	385	201	386
rect	201	385	202	386
rect	202	385	203	386
rect	203	385	204	386
rect	204	385	205	386
rect	205	385	206	386
rect	206	385	207	386
rect	207	385	208	386
rect	208	385	209	386
rect	210	385	211	386
rect	211	385	212	386
rect	212	385	213	386
rect	213	385	214	386
rect	214	385	215	386
rect	215	385	216	386
rect	216	385	217	386
rect	217	385	218	386
rect	218	385	219	386
rect	219	385	220	386
rect	220	385	221	386
rect	221	385	222	386
rect	222	385	223	386
rect	223	385	224	386
rect	224	385	225	386
rect	225	385	226	386
rect	226	385	227	386
rect	227	385	228	386
rect	228	385	229	386
rect	229	385	230	386
rect	230	385	231	386
rect	231	385	232	386
rect	232	385	233	386
rect	233	385	234	386
rect	234	385	235	386
rect	235	385	236	386
rect	236	385	237	386
rect	237	385	238	386
rect	238	385	239	386
rect	239	385	240	386
rect	240	385	241	386
rect	241	385	242	386
rect	242	385	243	386
rect	243	385	244	386
rect	244	385	245	386
rect	245	385	246	386
rect	246	385	247	386
rect	247	385	248	386
rect	248	385	249	386
rect	249	385	250	386
rect	250	385	251	386
rect	251	385	252	386
rect	252	385	253	386
rect	253	385	254	386
rect	254	385	255	386
rect	255	385	256	386
rect	256	385	257	386
rect	257	385	258	386
rect	258	385	259	386
rect	259	385	260	386
rect	260	385	261	386
rect	261	385	262	386
rect	262	385	263	386
rect	263	385	264	386
rect	264	385	265	386
rect	265	385	266	386
rect	266	385	267	386
rect	267	385	268	386
rect	268	385	269	386
rect	269	385	270	386
rect	270	385	271	386
rect	271	385	272	386
rect	272	385	273	386
rect	273	385	274	386
rect	274	385	275	386
rect	275	385	276	386
rect	276	385	277	386
rect	277	385	278	386
rect	278	385	279	386
rect	279	385	280	386
rect	280	385	281	386
rect	281	385	282	386
rect	282	385	283	386
rect	283	385	284	386
rect	284	385	285	386
rect	285	385	286	386
rect	286	385	287	386
rect	287	385	288	386
rect	288	385	289	386
rect	289	385	290	386
rect	290	385	291	386
rect	291	385	292	386
rect	292	385	293	386
rect	293	385	294	386
rect	294	385	295	386
rect	295	385	296	386
rect	296	385	297	386
rect	297	385	298	386
rect	298	385	299	386
rect	299	385	300	386
rect	300	385	301	386
rect	301	385	302	386
rect	302	385	303	386
rect	304	385	305	386
rect	305	385	306	386
rect	306	385	307	386
rect	307	385	308	386
rect	308	385	309	386
rect	309	385	310	386
rect	310	385	311	386
rect	311	385	312	386
rect	312	385	313	386
rect	313	385	314	386
rect	314	385	315	386
rect	315	385	316	386
rect	316	385	317	386
rect	317	385	318	386
rect	318	385	319	386
rect	319	385	320	386
rect	320	385	321	386
rect	321	385	322	386
rect	322	385	323	386
rect	323	385	324	386
rect	324	385	325	386
rect	325	385	326	386
rect	326	385	327	386
rect	327	385	328	386
rect	328	385	329	386
rect	329	385	330	386
rect	330	385	331	386
rect	331	385	332	386
rect	332	385	333	386
rect	333	385	334	386
rect	334	385	335	386
rect	335	385	336	386
rect	336	385	337	386
rect	337	385	338	386
rect	338	385	339	386
rect	339	385	340	386
rect	341	385	342	386
rect	342	385	343	386
rect	343	385	344	386
rect	344	385	345	386
rect	345	385	346	386
rect	346	385	347	386
rect	347	385	348	386
rect	348	385	349	386
rect	349	385	350	386
rect	350	385	351	386
rect	351	385	352	386
rect	352	385	353	386
rect	353	385	354	386
rect	354	385	355	386
rect	355	385	356	386
rect	357	385	358	386
rect	358	385	359	386
rect	359	385	360	386
rect	360	385	361	386
rect	361	385	362	386
rect	362	385	363	386
rect	363	385	364	386
rect	364	385	365	386
rect	365	385	366	386
rect	0	386	1	387
rect	1	386	2	387
rect	2	386	3	387
rect	3	386	4	387
rect	4	386	5	387
rect	5	386	6	387
rect	7	386	8	387
rect	8	386	9	387
rect	9	386	10	387
rect	10	386	11	387
rect	11	386	12	387
rect	12	386	13	387
rect	13	386	14	387
rect	14	386	15	387
rect	15	386	16	387
rect	16	386	17	387
rect	17	386	18	387
rect	18	386	19	387
rect	19	386	20	387
rect	20	386	21	387
rect	21	386	22	387
rect	23	386	24	387
rect	24	386	25	387
rect	25	386	26	387
rect	26	386	27	387
rect	27	386	28	387
rect	28	386	29	387
rect	30	386	31	387
rect	31	386	32	387
rect	32	386	33	387
rect	33	386	34	387
rect	34	386	35	387
rect	35	386	36	387
rect	37	386	38	387
rect	38	386	39	387
rect	39	386	40	387
rect	40	386	41	387
rect	41	386	42	387
rect	42	386	43	387
rect	44	386	45	387
rect	45	386	46	387
rect	46	386	47	387
rect	47	386	48	387
rect	48	386	49	387
rect	49	386	50	387
rect	51	386	52	387
rect	52	386	53	387
rect	53	386	54	387
rect	54	386	55	387
rect	55	386	56	387
rect	56	386	57	387
rect	57	386	58	387
rect	58	386	59	387
rect	59	386	60	387
rect	60	386	61	387
rect	61	386	62	387
rect	62	386	63	387
rect	63	386	64	387
rect	64	386	65	387
rect	65	386	66	387
rect	66	386	67	387
rect	67	386	68	387
rect	68	386	69	387
rect	69	386	70	387
rect	70	386	71	387
rect	71	386	72	387
rect	72	386	73	387
rect	73	386	74	387
rect	74	386	75	387
rect	75	386	76	387
rect	76	386	77	387
rect	77	386	78	387
rect	78	386	79	387
rect	79	386	80	387
rect	80	386	81	387
rect	81	386	82	387
rect	82	386	83	387
rect	83	386	84	387
rect	84	386	85	387
rect	85	386	86	387
rect	86	386	87	387
rect	87	386	88	387
rect	88	386	89	387
rect	89	386	90	387
rect	90	386	91	387
rect	91	386	92	387
rect	92	386	93	387
rect	93	386	94	387
rect	94	386	95	387
rect	95	386	96	387
rect	96	386	97	387
rect	97	386	98	387
rect	98	386	99	387
rect	99	386	100	387
rect	100	386	101	387
rect	101	386	102	387
rect	102	386	103	387
rect	103	386	104	387
rect	104	386	105	387
rect	105	386	106	387
rect	106	386	107	387
rect	107	386	108	387
rect	108	386	109	387
rect	109	386	110	387
rect	110	386	111	387
rect	111	386	112	387
rect	112	386	113	387
rect	113	386	114	387
rect	114	386	115	387
rect	115	386	116	387
rect	116	386	117	387
rect	117	386	118	387
rect	118	386	119	387
rect	119	386	120	387
rect	120	386	121	387
rect	121	386	122	387
rect	122	386	123	387
rect	123	386	124	387
rect	124	386	125	387
rect	125	386	126	387
rect	126	386	127	387
rect	127	386	128	387
rect	128	386	129	387
rect	129	386	130	387
rect	130	386	131	387
rect	131	386	132	387
rect	132	386	133	387
rect	133	386	134	387
rect	134	386	135	387
rect	135	386	136	387
rect	136	386	137	387
rect	137	386	138	387
rect	138	386	139	387
rect	139	386	140	387
rect	140	386	141	387
rect	141	386	142	387
rect	142	386	143	387
rect	143	386	144	387
rect	144	386	145	387
rect	145	386	146	387
rect	146	386	147	387
rect	147	386	148	387
rect	148	386	149	387
rect	149	386	150	387
rect	150	386	151	387
rect	151	386	152	387
rect	152	386	153	387
rect	153	386	154	387
rect	154	386	155	387
rect	155	386	156	387
rect	156	386	157	387
rect	157	386	158	387
rect	158	386	159	387
rect	160	386	161	387
rect	161	386	162	387
rect	162	386	163	387
rect	163	386	164	387
rect	164	386	165	387
rect	165	386	166	387
rect	166	386	167	387
rect	167	386	168	387
rect	168	386	169	387
rect	169	386	170	387
rect	170	386	171	387
rect	171	386	172	387
rect	172	386	173	387
rect	173	386	174	387
rect	174	386	175	387
rect	176	386	177	387
rect	177	386	178	387
rect	178	386	179	387
rect	179	386	180	387
rect	180	386	181	387
rect	181	386	182	387
rect	182	386	183	387
rect	183	386	184	387
rect	184	386	185	387
rect	185	386	186	387
rect	186	386	187	387
rect	187	386	188	387
rect	188	386	189	387
rect	189	386	190	387
rect	190	386	191	387
rect	191	386	192	387
rect	192	386	193	387
rect	193	386	194	387
rect	194	386	195	387
rect	195	386	196	387
rect	196	386	197	387
rect	197	386	198	387
rect	198	386	199	387
rect	199	386	200	387
rect	200	386	201	387
rect	201	386	202	387
rect	202	386	203	387
rect	203	386	204	387
rect	204	386	205	387
rect	205	386	206	387
rect	206	386	207	387
rect	207	386	208	387
rect	208	386	209	387
rect	210	386	211	387
rect	211	386	212	387
rect	212	386	213	387
rect	213	386	214	387
rect	214	386	215	387
rect	215	386	216	387
rect	216	386	217	387
rect	217	386	218	387
rect	218	386	219	387
rect	219	386	220	387
rect	220	386	221	387
rect	221	386	222	387
rect	222	386	223	387
rect	223	386	224	387
rect	224	386	225	387
rect	225	386	226	387
rect	226	386	227	387
rect	227	386	228	387
rect	228	386	229	387
rect	229	386	230	387
rect	230	386	231	387
rect	231	386	232	387
rect	232	386	233	387
rect	233	386	234	387
rect	234	386	235	387
rect	235	386	236	387
rect	236	386	237	387
rect	237	386	238	387
rect	238	386	239	387
rect	239	386	240	387
rect	240	386	241	387
rect	241	386	242	387
rect	242	386	243	387
rect	243	386	244	387
rect	244	386	245	387
rect	245	386	246	387
rect	246	386	247	387
rect	247	386	248	387
rect	248	386	249	387
rect	249	386	250	387
rect	250	386	251	387
rect	251	386	252	387
rect	252	386	253	387
rect	253	386	254	387
rect	254	386	255	387
rect	255	386	256	387
rect	256	386	257	387
rect	257	386	258	387
rect	258	386	259	387
rect	259	386	260	387
rect	260	386	261	387
rect	261	386	262	387
rect	262	386	263	387
rect	263	386	264	387
rect	264	386	265	387
rect	265	386	266	387
rect	266	386	267	387
rect	267	386	268	387
rect	268	386	269	387
rect	269	386	270	387
rect	270	386	271	387
rect	271	386	272	387
rect	272	386	273	387
rect	273	386	274	387
rect	274	386	275	387
rect	275	386	276	387
rect	276	386	277	387
rect	277	386	278	387
rect	278	386	279	387
rect	279	386	280	387
rect	280	386	281	387
rect	281	386	282	387
rect	282	386	283	387
rect	283	386	284	387
rect	284	386	285	387
rect	285	386	286	387
rect	286	386	287	387
rect	287	386	288	387
rect	288	386	289	387
rect	289	386	290	387
rect	290	386	291	387
rect	291	386	292	387
rect	292	386	293	387
rect	293	386	294	387
rect	294	386	295	387
rect	295	386	296	387
rect	296	386	297	387
rect	297	386	298	387
rect	298	386	299	387
rect	299	386	300	387
rect	300	386	301	387
rect	301	386	302	387
rect	302	386	303	387
rect	304	386	305	387
rect	305	386	306	387
rect	306	386	307	387
rect	307	386	308	387
rect	308	386	309	387
rect	309	386	310	387
rect	310	386	311	387
rect	311	386	312	387
rect	312	386	313	387
rect	313	386	314	387
rect	314	386	315	387
rect	315	386	316	387
rect	316	386	317	387
rect	317	386	318	387
rect	318	386	319	387
rect	319	386	320	387
rect	320	386	321	387
rect	321	386	322	387
rect	322	386	323	387
rect	323	386	324	387
rect	324	386	325	387
rect	325	386	326	387
rect	326	386	327	387
rect	327	386	328	387
rect	328	386	329	387
rect	329	386	330	387
rect	330	386	331	387
rect	331	386	332	387
rect	332	386	333	387
rect	333	386	334	387
rect	334	386	335	387
rect	335	386	336	387
rect	336	386	337	387
rect	337	386	338	387
rect	338	386	339	387
rect	339	386	340	387
rect	341	386	342	387
rect	342	386	343	387
rect	343	386	344	387
rect	344	386	345	387
rect	345	386	346	387
rect	346	386	347	387
rect	347	386	348	387
rect	348	386	349	387
rect	349	386	350	387
rect	350	386	351	387
rect	351	386	352	387
rect	352	386	353	387
rect	353	386	354	387
rect	354	386	355	387
rect	355	386	356	387
rect	357	386	358	387
rect	358	386	359	387
rect	359	386	360	387
rect	360	386	361	387
rect	361	386	362	387
rect	362	386	363	387
rect	363	386	364	387
rect	364	386	365	387
rect	365	386	366	387
rect	0	406	1	407
rect	1	406	2	407
rect	2	406	3	407
rect	3	406	4	407
rect	4	406	5	407
rect	5	406	6	407
rect	7	406	8	407
rect	8	406	9	407
rect	9	406	10	407
rect	10	406	11	407
rect	11	406	12	407
rect	12	406	13	407
rect	14	406	15	407
rect	15	406	16	407
rect	16	406	17	407
rect	17	406	18	407
rect	18	406	19	407
rect	19	406	20	407
rect	21	406	22	407
rect	22	406	23	407
rect	23	406	24	407
rect	24	406	25	407
rect	25	406	26	407
rect	26	406	27	407
rect	28	406	29	407
rect	29	406	30	407
rect	30	406	31	407
rect	31	406	32	407
rect	32	406	33	407
rect	33	406	34	407
rect	35	406	36	407
rect	36	406	37	407
rect	37	406	38	407
rect	38	406	39	407
rect	39	406	40	407
rect	40	406	41	407
rect	42	406	43	407
rect	43	406	44	407
rect	44	406	45	407
rect	45	406	46	407
rect	46	406	47	407
rect	47	406	48	407
rect	49	406	50	407
rect	50	406	51	407
rect	51	406	52	407
rect	52	406	53	407
rect	53	406	54	407
rect	54	406	55	407
rect	56	406	57	407
rect	57	406	58	407
rect	58	406	59	407
rect	59	406	60	407
rect	60	406	61	407
rect	61	406	62	407
rect	62	406	63	407
rect	63	406	64	407
rect	64	406	65	407
rect	65	406	66	407
rect	66	406	67	407
rect	67	406	68	407
rect	68	406	69	407
rect	69	406	70	407
rect	70	406	71	407
rect	71	406	72	407
rect	72	406	73	407
rect	73	406	74	407
rect	74	406	75	407
rect	75	406	76	407
rect	76	406	77	407
rect	77	406	78	407
rect	78	406	79	407
rect	79	406	80	407
rect	80	406	81	407
rect	81	406	82	407
rect	82	406	83	407
rect	83	406	84	407
rect	84	406	85	407
rect	85	406	86	407
rect	86	406	87	407
rect	87	406	88	407
rect	88	406	89	407
rect	90	406	91	407
rect	91	406	92	407
rect	92	406	93	407
rect	93	406	94	407
rect	94	406	95	407
rect	95	406	96	407
rect	96	406	97	407
rect	97	406	98	407
rect	98	406	99	407
rect	99	406	100	407
rect	100	406	101	407
rect	101	406	102	407
rect	102	406	103	407
rect	103	406	104	407
rect	104	406	105	407
rect	105	406	106	407
rect	106	406	107	407
rect	107	406	108	407
rect	108	406	109	407
rect	109	406	110	407
rect	110	406	111	407
rect	111	406	112	407
rect	112	406	113	407
rect	113	406	114	407
rect	114	406	115	407
rect	115	406	116	407
rect	116	406	117	407
rect	117	406	118	407
rect	118	406	119	407
rect	119	406	120	407
rect	120	406	121	407
rect	121	406	122	407
rect	122	406	123	407
rect	123	406	124	407
rect	124	406	125	407
rect	125	406	126	407
rect	126	406	127	407
rect	127	406	128	407
rect	128	406	129	407
rect	129	406	130	407
rect	130	406	131	407
rect	131	406	132	407
rect	132	406	133	407
rect	133	406	134	407
rect	134	406	135	407
rect	135	406	136	407
rect	136	406	137	407
rect	137	406	138	407
rect	139	406	140	407
rect	140	406	141	407
rect	141	406	142	407
rect	142	406	143	407
rect	143	406	144	407
rect	144	406	145	407
rect	145	406	146	407
rect	146	406	147	407
rect	147	406	148	407
rect	148	406	149	407
rect	149	406	150	407
rect	150	406	151	407
rect	151	406	152	407
rect	152	406	153	407
rect	153	406	154	407
rect	155	406	156	407
rect	156	406	157	407
rect	157	406	158	407
rect	158	406	159	407
rect	159	406	160	407
rect	160	406	161	407
rect	162	406	163	407
rect	163	406	164	407
rect	164	406	165	407
rect	165	406	166	407
rect	166	406	167	407
rect	167	406	168	407
rect	169	406	170	407
rect	170	406	171	407
rect	171	406	172	407
rect	172	406	173	407
rect	173	406	174	407
rect	174	406	175	407
rect	176	406	177	407
rect	177	406	178	407
rect	178	406	179	407
rect	179	406	180	407
rect	180	406	181	407
rect	181	406	182	407
rect	183	406	184	407
rect	184	406	185	407
rect	185	406	186	407
rect	186	406	187	407
rect	187	406	188	407
rect	188	406	189	407
rect	190	406	191	407
rect	191	406	192	407
rect	192	406	193	407
rect	193	406	194	407
rect	194	406	195	407
rect	195	406	196	407
rect	196	406	197	407
rect	197	406	198	407
rect	198	406	199	407
rect	199	406	200	407
rect	200	406	201	407
rect	201	406	202	407
rect	202	406	203	407
rect	203	406	204	407
rect	204	406	205	407
rect	205	406	206	407
rect	206	406	207	407
rect	207	406	208	407
rect	208	406	209	407
rect	209	406	210	407
rect	210	406	211	407
rect	211	406	212	407
rect	212	406	213	407
rect	213	406	214	407
rect	214	406	215	407
rect	215	406	216	407
rect	216	406	217	407
rect	217	406	218	407
rect	218	406	219	407
rect	219	406	220	407
rect	220	406	221	407
rect	221	406	222	407
rect	222	406	223	407
rect	223	406	224	407
rect	224	406	225	407
rect	225	406	226	407
rect	226	406	227	407
rect	227	406	228	407
rect	228	406	229	407
rect	229	406	230	407
rect	230	406	231	407
rect	231	406	232	407
rect	232	406	233	407
rect	233	406	234	407
rect	234	406	235	407
rect	235	406	236	407
rect	236	406	237	407
rect	237	406	238	407
rect	238	406	239	407
rect	239	406	240	407
rect	240	406	241	407
rect	241	406	242	407
rect	242	406	243	407
rect	243	406	244	407
rect	244	406	245	407
rect	245	406	246	407
rect	246	406	247	407
rect	247	406	248	407
rect	248	406	249	407
rect	249	406	250	407
rect	250	406	251	407
rect	251	406	252	407
rect	252	406	253	407
rect	253	406	254	407
rect	254	406	255	407
rect	255	406	256	407
rect	256	406	257	407
rect	257	406	258	407
rect	258	406	259	407
rect	259	406	260	407
rect	260	406	261	407
rect	261	406	262	407
rect	262	406	263	407
rect	263	406	264	407
rect	264	406	265	407
rect	265	406	266	407
rect	266	406	267	407
rect	267	406	268	407
rect	268	406	269	407
rect	269	406	270	407
rect	270	406	271	407
rect	271	406	272	407
rect	272	406	273	407
rect	273	406	274	407
rect	274	406	275	407
rect	275	406	276	407
rect	276	406	277	407
rect	277	406	278	407
rect	278	406	279	407
rect	279	406	280	407
rect	280	406	281	407
rect	281	406	282	407
rect	282	406	283	407
rect	283	406	284	407
rect	284	406	285	407
rect	285	406	286	407
rect	286	406	287	407
rect	287	406	288	407
rect	288	406	289	407
rect	289	406	290	407
rect	290	406	291	407
rect	291	406	292	407
rect	292	406	293	407
rect	293	406	294	407
rect	294	406	295	407
rect	296	406	297	407
rect	297	406	298	407
rect	298	406	299	407
rect	299	406	300	407
rect	300	406	301	407
rect	301	406	302	407
rect	302	406	303	407
rect	303	406	304	407
rect	304	406	305	407
rect	305	406	306	407
rect	306	406	307	407
rect	307	406	308	407
rect	308	406	309	407
rect	309	406	310	407
rect	310	406	311	407
rect	311	406	312	407
rect	312	406	313	407
rect	313	406	314	407
rect	314	406	315	407
rect	315	406	316	407
rect	316	406	317	407
rect	317	406	318	407
rect	318	406	319	407
rect	319	406	320	407
rect	321	406	322	407
rect	322	406	323	407
rect	323	406	324	407
rect	324	406	325	407
rect	325	406	326	407
rect	326	406	327	407
rect	327	406	328	407
rect	328	406	329	407
rect	329	406	330	407
rect	330	406	331	407
rect	331	406	332	407
rect	332	406	333	407
rect	0	407	1	408
rect	1	407	2	408
rect	2	407	3	408
rect	3	407	4	408
rect	4	407	5	408
rect	5	407	6	408
rect	7	407	8	408
rect	8	407	9	408
rect	9	407	10	408
rect	10	407	11	408
rect	11	407	12	408
rect	12	407	13	408
rect	14	407	15	408
rect	15	407	16	408
rect	16	407	17	408
rect	17	407	18	408
rect	18	407	19	408
rect	19	407	20	408
rect	21	407	22	408
rect	22	407	23	408
rect	23	407	24	408
rect	24	407	25	408
rect	25	407	26	408
rect	26	407	27	408
rect	28	407	29	408
rect	29	407	30	408
rect	30	407	31	408
rect	31	407	32	408
rect	32	407	33	408
rect	33	407	34	408
rect	35	407	36	408
rect	36	407	37	408
rect	37	407	38	408
rect	38	407	39	408
rect	39	407	40	408
rect	40	407	41	408
rect	42	407	43	408
rect	43	407	44	408
rect	44	407	45	408
rect	45	407	46	408
rect	46	407	47	408
rect	47	407	48	408
rect	49	407	50	408
rect	50	407	51	408
rect	51	407	52	408
rect	52	407	53	408
rect	53	407	54	408
rect	54	407	55	408
rect	56	407	57	408
rect	57	407	58	408
rect	58	407	59	408
rect	59	407	60	408
rect	60	407	61	408
rect	61	407	62	408
rect	62	407	63	408
rect	63	407	64	408
rect	64	407	65	408
rect	65	407	66	408
rect	66	407	67	408
rect	67	407	68	408
rect	68	407	69	408
rect	69	407	70	408
rect	70	407	71	408
rect	71	407	72	408
rect	72	407	73	408
rect	73	407	74	408
rect	74	407	75	408
rect	75	407	76	408
rect	76	407	77	408
rect	77	407	78	408
rect	78	407	79	408
rect	79	407	80	408
rect	80	407	81	408
rect	81	407	82	408
rect	82	407	83	408
rect	83	407	84	408
rect	84	407	85	408
rect	85	407	86	408
rect	86	407	87	408
rect	87	407	88	408
rect	88	407	89	408
rect	90	407	91	408
rect	91	407	92	408
rect	92	407	93	408
rect	93	407	94	408
rect	94	407	95	408
rect	95	407	96	408
rect	96	407	97	408
rect	97	407	98	408
rect	98	407	99	408
rect	99	407	100	408
rect	100	407	101	408
rect	101	407	102	408
rect	102	407	103	408
rect	103	407	104	408
rect	104	407	105	408
rect	105	407	106	408
rect	106	407	107	408
rect	107	407	108	408
rect	108	407	109	408
rect	109	407	110	408
rect	110	407	111	408
rect	111	407	112	408
rect	112	407	113	408
rect	113	407	114	408
rect	114	407	115	408
rect	115	407	116	408
rect	116	407	117	408
rect	117	407	118	408
rect	118	407	119	408
rect	119	407	120	408
rect	120	407	121	408
rect	121	407	122	408
rect	122	407	123	408
rect	123	407	124	408
rect	124	407	125	408
rect	125	407	126	408
rect	126	407	127	408
rect	127	407	128	408
rect	128	407	129	408
rect	129	407	130	408
rect	130	407	131	408
rect	131	407	132	408
rect	132	407	133	408
rect	133	407	134	408
rect	134	407	135	408
rect	135	407	136	408
rect	136	407	137	408
rect	137	407	138	408
rect	139	407	140	408
rect	140	407	141	408
rect	141	407	142	408
rect	142	407	143	408
rect	143	407	144	408
rect	144	407	145	408
rect	145	407	146	408
rect	146	407	147	408
rect	147	407	148	408
rect	148	407	149	408
rect	149	407	150	408
rect	150	407	151	408
rect	151	407	152	408
rect	152	407	153	408
rect	153	407	154	408
rect	155	407	156	408
rect	156	407	157	408
rect	157	407	158	408
rect	158	407	159	408
rect	159	407	160	408
rect	160	407	161	408
rect	162	407	163	408
rect	163	407	164	408
rect	164	407	165	408
rect	165	407	166	408
rect	166	407	167	408
rect	167	407	168	408
rect	169	407	170	408
rect	170	407	171	408
rect	171	407	172	408
rect	172	407	173	408
rect	173	407	174	408
rect	174	407	175	408
rect	176	407	177	408
rect	177	407	178	408
rect	178	407	179	408
rect	179	407	180	408
rect	180	407	181	408
rect	181	407	182	408
rect	183	407	184	408
rect	184	407	185	408
rect	185	407	186	408
rect	186	407	187	408
rect	187	407	188	408
rect	188	407	189	408
rect	190	407	191	408
rect	191	407	192	408
rect	192	407	193	408
rect	193	407	194	408
rect	194	407	195	408
rect	195	407	196	408
rect	196	407	197	408
rect	197	407	198	408
rect	198	407	199	408
rect	199	407	200	408
rect	200	407	201	408
rect	201	407	202	408
rect	202	407	203	408
rect	203	407	204	408
rect	204	407	205	408
rect	205	407	206	408
rect	206	407	207	408
rect	207	407	208	408
rect	208	407	209	408
rect	209	407	210	408
rect	210	407	211	408
rect	211	407	212	408
rect	212	407	213	408
rect	213	407	214	408
rect	214	407	215	408
rect	215	407	216	408
rect	216	407	217	408
rect	217	407	218	408
rect	218	407	219	408
rect	219	407	220	408
rect	220	407	221	408
rect	221	407	222	408
rect	222	407	223	408
rect	223	407	224	408
rect	224	407	225	408
rect	225	407	226	408
rect	226	407	227	408
rect	227	407	228	408
rect	228	407	229	408
rect	229	407	230	408
rect	230	407	231	408
rect	231	407	232	408
rect	232	407	233	408
rect	233	407	234	408
rect	234	407	235	408
rect	235	407	236	408
rect	236	407	237	408
rect	237	407	238	408
rect	238	407	239	408
rect	239	407	240	408
rect	240	407	241	408
rect	241	407	242	408
rect	242	407	243	408
rect	243	407	244	408
rect	244	407	245	408
rect	245	407	246	408
rect	246	407	247	408
rect	247	407	248	408
rect	248	407	249	408
rect	249	407	250	408
rect	250	407	251	408
rect	251	407	252	408
rect	252	407	253	408
rect	253	407	254	408
rect	254	407	255	408
rect	255	407	256	408
rect	256	407	257	408
rect	257	407	258	408
rect	258	407	259	408
rect	259	407	260	408
rect	260	407	261	408
rect	261	407	262	408
rect	262	407	263	408
rect	263	407	264	408
rect	264	407	265	408
rect	265	407	266	408
rect	266	407	267	408
rect	267	407	268	408
rect	268	407	269	408
rect	269	407	270	408
rect	270	407	271	408
rect	271	407	272	408
rect	272	407	273	408
rect	273	407	274	408
rect	274	407	275	408
rect	275	407	276	408
rect	276	407	277	408
rect	277	407	278	408
rect	278	407	279	408
rect	279	407	280	408
rect	280	407	281	408
rect	281	407	282	408
rect	282	407	283	408
rect	283	407	284	408
rect	284	407	285	408
rect	285	407	286	408
rect	286	407	287	408
rect	287	407	288	408
rect	288	407	289	408
rect	289	407	290	408
rect	290	407	291	408
rect	291	407	292	408
rect	292	407	293	408
rect	293	407	294	408
rect	294	407	295	408
rect	296	407	297	408
rect	297	407	298	408
rect	298	407	299	408
rect	299	407	300	408
rect	300	407	301	408
rect	301	407	302	408
rect	302	407	303	408
rect	303	407	304	408
rect	304	407	305	408
rect	305	407	306	408
rect	306	407	307	408
rect	307	407	308	408
rect	308	407	309	408
rect	309	407	310	408
rect	310	407	311	408
rect	311	407	312	408
rect	312	407	313	408
rect	313	407	314	408
rect	314	407	315	408
rect	315	407	316	408
rect	316	407	317	408
rect	317	407	318	408
rect	318	407	319	408
rect	319	407	320	408
rect	321	407	322	408
rect	322	407	323	408
rect	323	407	324	408
rect	324	407	325	408
rect	325	407	326	408
rect	326	407	327	408
rect	327	407	328	408
rect	328	407	329	408
rect	329	407	330	408
rect	330	407	331	408
rect	331	407	332	408
rect	332	407	333	408
rect	0	408	1	409
rect	1	408	2	409
rect	2	408	3	409
rect	3	408	4	409
rect	4	408	5	409
rect	5	408	6	409
rect	7	408	8	409
rect	8	408	9	409
rect	9	408	10	409
rect	10	408	11	409
rect	11	408	12	409
rect	12	408	13	409
rect	14	408	15	409
rect	15	408	16	409
rect	16	408	17	409
rect	17	408	18	409
rect	18	408	19	409
rect	19	408	20	409
rect	21	408	22	409
rect	22	408	23	409
rect	23	408	24	409
rect	24	408	25	409
rect	25	408	26	409
rect	26	408	27	409
rect	28	408	29	409
rect	29	408	30	409
rect	30	408	31	409
rect	31	408	32	409
rect	32	408	33	409
rect	33	408	34	409
rect	35	408	36	409
rect	36	408	37	409
rect	37	408	38	409
rect	38	408	39	409
rect	39	408	40	409
rect	40	408	41	409
rect	42	408	43	409
rect	43	408	44	409
rect	44	408	45	409
rect	45	408	46	409
rect	46	408	47	409
rect	47	408	48	409
rect	49	408	50	409
rect	50	408	51	409
rect	51	408	52	409
rect	52	408	53	409
rect	53	408	54	409
rect	54	408	55	409
rect	56	408	57	409
rect	57	408	58	409
rect	58	408	59	409
rect	59	408	60	409
rect	60	408	61	409
rect	61	408	62	409
rect	62	408	63	409
rect	63	408	64	409
rect	64	408	65	409
rect	65	408	66	409
rect	66	408	67	409
rect	67	408	68	409
rect	68	408	69	409
rect	69	408	70	409
rect	70	408	71	409
rect	71	408	72	409
rect	72	408	73	409
rect	73	408	74	409
rect	74	408	75	409
rect	75	408	76	409
rect	76	408	77	409
rect	77	408	78	409
rect	78	408	79	409
rect	79	408	80	409
rect	80	408	81	409
rect	81	408	82	409
rect	82	408	83	409
rect	83	408	84	409
rect	84	408	85	409
rect	85	408	86	409
rect	86	408	87	409
rect	87	408	88	409
rect	88	408	89	409
rect	90	408	91	409
rect	91	408	92	409
rect	92	408	93	409
rect	93	408	94	409
rect	94	408	95	409
rect	95	408	96	409
rect	96	408	97	409
rect	97	408	98	409
rect	98	408	99	409
rect	99	408	100	409
rect	100	408	101	409
rect	101	408	102	409
rect	102	408	103	409
rect	103	408	104	409
rect	104	408	105	409
rect	105	408	106	409
rect	106	408	107	409
rect	107	408	108	409
rect	108	408	109	409
rect	109	408	110	409
rect	110	408	111	409
rect	111	408	112	409
rect	112	408	113	409
rect	113	408	114	409
rect	114	408	115	409
rect	115	408	116	409
rect	116	408	117	409
rect	117	408	118	409
rect	118	408	119	409
rect	119	408	120	409
rect	120	408	121	409
rect	121	408	122	409
rect	122	408	123	409
rect	123	408	124	409
rect	124	408	125	409
rect	125	408	126	409
rect	126	408	127	409
rect	127	408	128	409
rect	128	408	129	409
rect	129	408	130	409
rect	130	408	131	409
rect	131	408	132	409
rect	132	408	133	409
rect	133	408	134	409
rect	134	408	135	409
rect	135	408	136	409
rect	136	408	137	409
rect	137	408	138	409
rect	139	408	140	409
rect	140	408	141	409
rect	141	408	142	409
rect	142	408	143	409
rect	143	408	144	409
rect	144	408	145	409
rect	145	408	146	409
rect	146	408	147	409
rect	147	408	148	409
rect	148	408	149	409
rect	149	408	150	409
rect	150	408	151	409
rect	151	408	152	409
rect	152	408	153	409
rect	153	408	154	409
rect	155	408	156	409
rect	156	408	157	409
rect	157	408	158	409
rect	158	408	159	409
rect	159	408	160	409
rect	160	408	161	409
rect	162	408	163	409
rect	163	408	164	409
rect	164	408	165	409
rect	165	408	166	409
rect	166	408	167	409
rect	167	408	168	409
rect	169	408	170	409
rect	170	408	171	409
rect	171	408	172	409
rect	172	408	173	409
rect	173	408	174	409
rect	174	408	175	409
rect	176	408	177	409
rect	177	408	178	409
rect	178	408	179	409
rect	179	408	180	409
rect	180	408	181	409
rect	181	408	182	409
rect	183	408	184	409
rect	184	408	185	409
rect	185	408	186	409
rect	186	408	187	409
rect	187	408	188	409
rect	188	408	189	409
rect	190	408	191	409
rect	191	408	192	409
rect	192	408	193	409
rect	193	408	194	409
rect	194	408	195	409
rect	195	408	196	409
rect	196	408	197	409
rect	197	408	198	409
rect	198	408	199	409
rect	199	408	200	409
rect	200	408	201	409
rect	201	408	202	409
rect	202	408	203	409
rect	203	408	204	409
rect	204	408	205	409
rect	205	408	206	409
rect	206	408	207	409
rect	207	408	208	409
rect	208	408	209	409
rect	209	408	210	409
rect	210	408	211	409
rect	211	408	212	409
rect	212	408	213	409
rect	213	408	214	409
rect	214	408	215	409
rect	215	408	216	409
rect	216	408	217	409
rect	217	408	218	409
rect	218	408	219	409
rect	219	408	220	409
rect	220	408	221	409
rect	221	408	222	409
rect	222	408	223	409
rect	223	408	224	409
rect	224	408	225	409
rect	225	408	226	409
rect	226	408	227	409
rect	227	408	228	409
rect	228	408	229	409
rect	229	408	230	409
rect	230	408	231	409
rect	231	408	232	409
rect	232	408	233	409
rect	233	408	234	409
rect	234	408	235	409
rect	235	408	236	409
rect	236	408	237	409
rect	237	408	238	409
rect	238	408	239	409
rect	239	408	240	409
rect	240	408	241	409
rect	241	408	242	409
rect	242	408	243	409
rect	243	408	244	409
rect	244	408	245	409
rect	245	408	246	409
rect	246	408	247	409
rect	247	408	248	409
rect	248	408	249	409
rect	249	408	250	409
rect	250	408	251	409
rect	251	408	252	409
rect	252	408	253	409
rect	253	408	254	409
rect	254	408	255	409
rect	255	408	256	409
rect	256	408	257	409
rect	257	408	258	409
rect	258	408	259	409
rect	259	408	260	409
rect	260	408	261	409
rect	261	408	262	409
rect	262	408	263	409
rect	263	408	264	409
rect	264	408	265	409
rect	265	408	266	409
rect	266	408	267	409
rect	267	408	268	409
rect	268	408	269	409
rect	269	408	270	409
rect	270	408	271	409
rect	271	408	272	409
rect	272	408	273	409
rect	273	408	274	409
rect	274	408	275	409
rect	275	408	276	409
rect	276	408	277	409
rect	277	408	278	409
rect	278	408	279	409
rect	279	408	280	409
rect	280	408	281	409
rect	281	408	282	409
rect	282	408	283	409
rect	283	408	284	409
rect	284	408	285	409
rect	285	408	286	409
rect	286	408	287	409
rect	287	408	288	409
rect	288	408	289	409
rect	289	408	290	409
rect	290	408	291	409
rect	291	408	292	409
rect	292	408	293	409
rect	293	408	294	409
rect	294	408	295	409
rect	296	408	297	409
rect	297	408	298	409
rect	298	408	299	409
rect	299	408	300	409
rect	300	408	301	409
rect	301	408	302	409
rect	302	408	303	409
rect	303	408	304	409
rect	304	408	305	409
rect	305	408	306	409
rect	306	408	307	409
rect	307	408	308	409
rect	308	408	309	409
rect	309	408	310	409
rect	310	408	311	409
rect	311	408	312	409
rect	312	408	313	409
rect	313	408	314	409
rect	314	408	315	409
rect	315	408	316	409
rect	316	408	317	409
rect	317	408	318	409
rect	318	408	319	409
rect	319	408	320	409
rect	321	408	322	409
rect	322	408	323	409
rect	323	408	324	409
rect	324	408	325	409
rect	325	408	326	409
rect	326	408	327	409
rect	327	408	328	409
rect	328	408	329	409
rect	329	408	330	409
rect	330	408	331	409
rect	331	408	332	409
rect	332	408	333	409
rect	0	409	1	410
rect	1	409	2	410
rect	2	409	3	410
rect	3	409	4	410
rect	4	409	5	410
rect	5	409	6	410
rect	7	409	8	410
rect	8	409	9	410
rect	9	409	10	410
rect	10	409	11	410
rect	11	409	12	410
rect	12	409	13	410
rect	14	409	15	410
rect	15	409	16	410
rect	16	409	17	410
rect	17	409	18	410
rect	18	409	19	410
rect	19	409	20	410
rect	21	409	22	410
rect	22	409	23	410
rect	23	409	24	410
rect	24	409	25	410
rect	25	409	26	410
rect	26	409	27	410
rect	28	409	29	410
rect	29	409	30	410
rect	30	409	31	410
rect	31	409	32	410
rect	32	409	33	410
rect	33	409	34	410
rect	35	409	36	410
rect	36	409	37	410
rect	37	409	38	410
rect	38	409	39	410
rect	39	409	40	410
rect	40	409	41	410
rect	42	409	43	410
rect	43	409	44	410
rect	44	409	45	410
rect	45	409	46	410
rect	46	409	47	410
rect	47	409	48	410
rect	49	409	50	410
rect	50	409	51	410
rect	51	409	52	410
rect	52	409	53	410
rect	53	409	54	410
rect	54	409	55	410
rect	56	409	57	410
rect	57	409	58	410
rect	58	409	59	410
rect	59	409	60	410
rect	60	409	61	410
rect	61	409	62	410
rect	62	409	63	410
rect	63	409	64	410
rect	64	409	65	410
rect	65	409	66	410
rect	66	409	67	410
rect	67	409	68	410
rect	68	409	69	410
rect	69	409	70	410
rect	70	409	71	410
rect	71	409	72	410
rect	72	409	73	410
rect	73	409	74	410
rect	74	409	75	410
rect	75	409	76	410
rect	76	409	77	410
rect	77	409	78	410
rect	78	409	79	410
rect	79	409	80	410
rect	80	409	81	410
rect	81	409	82	410
rect	82	409	83	410
rect	83	409	84	410
rect	84	409	85	410
rect	85	409	86	410
rect	86	409	87	410
rect	87	409	88	410
rect	88	409	89	410
rect	90	409	91	410
rect	91	409	92	410
rect	92	409	93	410
rect	93	409	94	410
rect	94	409	95	410
rect	95	409	96	410
rect	96	409	97	410
rect	97	409	98	410
rect	98	409	99	410
rect	99	409	100	410
rect	100	409	101	410
rect	101	409	102	410
rect	102	409	103	410
rect	103	409	104	410
rect	104	409	105	410
rect	105	409	106	410
rect	106	409	107	410
rect	107	409	108	410
rect	108	409	109	410
rect	109	409	110	410
rect	110	409	111	410
rect	111	409	112	410
rect	112	409	113	410
rect	113	409	114	410
rect	114	409	115	410
rect	115	409	116	410
rect	116	409	117	410
rect	117	409	118	410
rect	118	409	119	410
rect	119	409	120	410
rect	120	409	121	410
rect	121	409	122	410
rect	122	409	123	410
rect	123	409	124	410
rect	124	409	125	410
rect	125	409	126	410
rect	126	409	127	410
rect	127	409	128	410
rect	128	409	129	410
rect	129	409	130	410
rect	130	409	131	410
rect	131	409	132	410
rect	132	409	133	410
rect	133	409	134	410
rect	134	409	135	410
rect	135	409	136	410
rect	136	409	137	410
rect	137	409	138	410
rect	139	409	140	410
rect	140	409	141	410
rect	141	409	142	410
rect	142	409	143	410
rect	143	409	144	410
rect	144	409	145	410
rect	145	409	146	410
rect	146	409	147	410
rect	147	409	148	410
rect	148	409	149	410
rect	149	409	150	410
rect	150	409	151	410
rect	151	409	152	410
rect	152	409	153	410
rect	153	409	154	410
rect	155	409	156	410
rect	156	409	157	410
rect	157	409	158	410
rect	158	409	159	410
rect	159	409	160	410
rect	160	409	161	410
rect	162	409	163	410
rect	163	409	164	410
rect	164	409	165	410
rect	165	409	166	410
rect	166	409	167	410
rect	167	409	168	410
rect	169	409	170	410
rect	170	409	171	410
rect	171	409	172	410
rect	172	409	173	410
rect	173	409	174	410
rect	174	409	175	410
rect	176	409	177	410
rect	177	409	178	410
rect	178	409	179	410
rect	179	409	180	410
rect	180	409	181	410
rect	181	409	182	410
rect	183	409	184	410
rect	184	409	185	410
rect	185	409	186	410
rect	186	409	187	410
rect	187	409	188	410
rect	188	409	189	410
rect	190	409	191	410
rect	191	409	192	410
rect	192	409	193	410
rect	193	409	194	410
rect	194	409	195	410
rect	195	409	196	410
rect	196	409	197	410
rect	197	409	198	410
rect	198	409	199	410
rect	199	409	200	410
rect	200	409	201	410
rect	201	409	202	410
rect	202	409	203	410
rect	203	409	204	410
rect	204	409	205	410
rect	205	409	206	410
rect	206	409	207	410
rect	207	409	208	410
rect	208	409	209	410
rect	209	409	210	410
rect	210	409	211	410
rect	211	409	212	410
rect	212	409	213	410
rect	213	409	214	410
rect	214	409	215	410
rect	215	409	216	410
rect	216	409	217	410
rect	217	409	218	410
rect	218	409	219	410
rect	219	409	220	410
rect	220	409	221	410
rect	221	409	222	410
rect	222	409	223	410
rect	223	409	224	410
rect	224	409	225	410
rect	225	409	226	410
rect	226	409	227	410
rect	227	409	228	410
rect	228	409	229	410
rect	229	409	230	410
rect	230	409	231	410
rect	231	409	232	410
rect	232	409	233	410
rect	233	409	234	410
rect	234	409	235	410
rect	235	409	236	410
rect	236	409	237	410
rect	237	409	238	410
rect	238	409	239	410
rect	239	409	240	410
rect	240	409	241	410
rect	241	409	242	410
rect	242	409	243	410
rect	243	409	244	410
rect	244	409	245	410
rect	245	409	246	410
rect	246	409	247	410
rect	247	409	248	410
rect	248	409	249	410
rect	249	409	250	410
rect	250	409	251	410
rect	251	409	252	410
rect	252	409	253	410
rect	253	409	254	410
rect	254	409	255	410
rect	255	409	256	410
rect	256	409	257	410
rect	257	409	258	410
rect	258	409	259	410
rect	259	409	260	410
rect	260	409	261	410
rect	261	409	262	410
rect	262	409	263	410
rect	263	409	264	410
rect	264	409	265	410
rect	265	409	266	410
rect	266	409	267	410
rect	267	409	268	410
rect	268	409	269	410
rect	269	409	270	410
rect	270	409	271	410
rect	271	409	272	410
rect	272	409	273	410
rect	273	409	274	410
rect	274	409	275	410
rect	275	409	276	410
rect	276	409	277	410
rect	277	409	278	410
rect	278	409	279	410
rect	279	409	280	410
rect	280	409	281	410
rect	281	409	282	410
rect	282	409	283	410
rect	283	409	284	410
rect	284	409	285	410
rect	285	409	286	410
rect	286	409	287	410
rect	287	409	288	410
rect	288	409	289	410
rect	289	409	290	410
rect	290	409	291	410
rect	291	409	292	410
rect	292	409	293	410
rect	293	409	294	410
rect	294	409	295	410
rect	296	409	297	410
rect	297	409	298	410
rect	298	409	299	410
rect	299	409	300	410
rect	300	409	301	410
rect	301	409	302	410
rect	302	409	303	410
rect	303	409	304	410
rect	304	409	305	410
rect	305	409	306	410
rect	306	409	307	410
rect	307	409	308	410
rect	308	409	309	410
rect	309	409	310	410
rect	310	409	311	410
rect	311	409	312	410
rect	312	409	313	410
rect	313	409	314	410
rect	314	409	315	410
rect	315	409	316	410
rect	316	409	317	410
rect	317	409	318	410
rect	318	409	319	410
rect	319	409	320	410
rect	321	409	322	410
rect	322	409	323	410
rect	323	409	324	410
rect	324	409	325	410
rect	325	409	326	410
rect	326	409	327	410
rect	327	409	328	410
rect	328	409	329	410
rect	329	409	330	410
rect	330	409	331	410
rect	331	409	332	410
rect	332	409	333	410
rect	0	410	1	411
rect	1	410	2	411
rect	2	410	3	411
rect	3	410	4	411
rect	4	410	5	411
rect	5	410	6	411
rect	7	410	8	411
rect	8	410	9	411
rect	9	410	10	411
rect	10	410	11	411
rect	11	410	12	411
rect	12	410	13	411
rect	14	410	15	411
rect	15	410	16	411
rect	16	410	17	411
rect	17	410	18	411
rect	18	410	19	411
rect	19	410	20	411
rect	21	410	22	411
rect	22	410	23	411
rect	23	410	24	411
rect	24	410	25	411
rect	25	410	26	411
rect	26	410	27	411
rect	28	410	29	411
rect	29	410	30	411
rect	30	410	31	411
rect	31	410	32	411
rect	32	410	33	411
rect	33	410	34	411
rect	35	410	36	411
rect	36	410	37	411
rect	37	410	38	411
rect	38	410	39	411
rect	39	410	40	411
rect	40	410	41	411
rect	42	410	43	411
rect	43	410	44	411
rect	44	410	45	411
rect	45	410	46	411
rect	46	410	47	411
rect	47	410	48	411
rect	49	410	50	411
rect	50	410	51	411
rect	51	410	52	411
rect	52	410	53	411
rect	53	410	54	411
rect	54	410	55	411
rect	56	410	57	411
rect	57	410	58	411
rect	58	410	59	411
rect	59	410	60	411
rect	60	410	61	411
rect	61	410	62	411
rect	62	410	63	411
rect	63	410	64	411
rect	64	410	65	411
rect	65	410	66	411
rect	66	410	67	411
rect	67	410	68	411
rect	68	410	69	411
rect	69	410	70	411
rect	70	410	71	411
rect	71	410	72	411
rect	72	410	73	411
rect	73	410	74	411
rect	74	410	75	411
rect	75	410	76	411
rect	76	410	77	411
rect	77	410	78	411
rect	78	410	79	411
rect	79	410	80	411
rect	80	410	81	411
rect	81	410	82	411
rect	82	410	83	411
rect	83	410	84	411
rect	84	410	85	411
rect	85	410	86	411
rect	86	410	87	411
rect	87	410	88	411
rect	88	410	89	411
rect	90	410	91	411
rect	91	410	92	411
rect	92	410	93	411
rect	93	410	94	411
rect	94	410	95	411
rect	95	410	96	411
rect	96	410	97	411
rect	97	410	98	411
rect	98	410	99	411
rect	99	410	100	411
rect	100	410	101	411
rect	101	410	102	411
rect	102	410	103	411
rect	103	410	104	411
rect	104	410	105	411
rect	105	410	106	411
rect	106	410	107	411
rect	107	410	108	411
rect	108	410	109	411
rect	109	410	110	411
rect	110	410	111	411
rect	111	410	112	411
rect	112	410	113	411
rect	113	410	114	411
rect	114	410	115	411
rect	115	410	116	411
rect	116	410	117	411
rect	117	410	118	411
rect	118	410	119	411
rect	119	410	120	411
rect	120	410	121	411
rect	121	410	122	411
rect	122	410	123	411
rect	123	410	124	411
rect	124	410	125	411
rect	125	410	126	411
rect	126	410	127	411
rect	127	410	128	411
rect	128	410	129	411
rect	129	410	130	411
rect	130	410	131	411
rect	131	410	132	411
rect	132	410	133	411
rect	133	410	134	411
rect	134	410	135	411
rect	135	410	136	411
rect	136	410	137	411
rect	137	410	138	411
rect	139	410	140	411
rect	140	410	141	411
rect	141	410	142	411
rect	142	410	143	411
rect	143	410	144	411
rect	144	410	145	411
rect	145	410	146	411
rect	146	410	147	411
rect	147	410	148	411
rect	148	410	149	411
rect	149	410	150	411
rect	150	410	151	411
rect	151	410	152	411
rect	152	410	153	411
rect	153	410	154	411
rect	155	410	156	411
rect	156	410	157	411
rect	157	410	158	411
rect	158	410	159	411
rect	159	410	160	411
rect	160	410	161	411
rect	162	410	163	411
rect	163	410	164	411
rect	164	410	165	411
rect	165	410	166	411
rect	166	410	167	411
rect	167	410	168	411
rect	169	410	170	411
rect	170	410	171	411
rect	171	410	172	411
rect	172	410	173	411
rect	173	410	174	411
rect	174	410	175	411
rect	176	410	177	411
rect	177	410	178	411
rect	178	410	179	411
rect	179	410	180	411
rect	180	410	181	411
rect	181	410	182	411
rect	183	410	184	411
rect	184	410	185	411
rect	185	410	186	411
rect	186	410	187	411
rect	187	410	188	411
rect	188	410	189	411
rect	190	410	191	411
rect	191	410	192	411
rect	192	410	193	411
rect	193	410	194	411
rect	194	410	195	411
rect	195	410	196	411
rect	196	410	197	411
rect	197	410	198	411
rect	198	410	199	411
rect	199	410	200	411
rect	200	410	201	411
rect	201	410	202	411
rect	202	410	203	411
rect	203	410	204	411
rect	204	410	205	411
rect	205	410	206	411
rect	206	410	207	411
rect	207	410	208	411
rect	208	410	209	411
rect	209	410	210	411
rect	210	410	211	411
rect	211	410	212	411
rect	212	410	213	411
rect	213	410	214	411
rect	214	410	215	411
rect	215	410	216	411
rect	216	410	217	411
rect	217	410	218	411
rect	218	410	219	411
rect	219	410	220	411
rect	220	410	221	411
rect	221	410	222	411
rect	222	410	223	411
rect	223	410	224	411
rect	224	410	225	411
rect	225	410	226	411
rect	226	410	227	411
rect	227	410	228	411
rect	228	410	229	411
rect	229	410	230	411
rect	230	410	231	411
rect	231	410	232	411
rect	232	410	233	411
rect	233	410	234	411
rect	234	410	235	411
rect	235	410	236	411
rect	236	410	237	411
rect	237	410	238	411
rect	238	410	239	411
rect	239	410	240	411
rect	240	410	241	411
rect	241	410	242	411
rect	242	410	243	411
rect	243	410	244	411
rect	244	410	245	411
rect	245	410	246	411
rect	246	410	247	411
rect	247	410	248	411
rect	248	410	249	411
rect	249	410	250	411
rect	250	410	251	411
rect	251	410	252	411
rect	252	410	253	411
rect	253	410	254	411
rect	254	410	255	411
rect	255	410	256	411
rect	256	410	257	411
rect	257	410	258	411
rect	258	410	259	411
rect	259	410	260	411
rect	260	410	261	411
rect	261	410	262	411
rect	262	410	263	411
rect	263	410	264	411
rect	264	410	265	411
rect	265	410	266	411
rect	266	410	267	411
rect	267	410	268	411
rect	268	410	269	411
rect	269	410	270	411
rect	270	410	271	411
rect	271	410	272	411
rect	272	410	273	411
rect	273	410	274	411
rect	274	410	275	411
rect	275	410	276	411
rect	276	410	277	411
rect	277	410	278	411
rect	278	410	279	411
rect	279	410	280	411
rect	280	410	281	411
rect	281	410	282	411
rect	282	410	283	411
rect	283	410	284	411
rect	284	410	285	411
rect	285	410	286	411
rect	286	410	287	411
rect	287	410	288	411
rect	288	410	289	411
rect	289	410	290	411
rect	290	410	291	411
rect	291	410	292	411
rect	292	410	293	411
rect	293	410	294	411
rect	294	410	295	411
rect	296	410	297	411
rect	297	410	298	411
rect	298	410	299	411
rect	299	410	300	411
rect	300	410	301	411
rect	301	410	302	411
rect	302	410	303	411
rect	303	410	304	411
rect	304	410	305	411
rect	305	410	306	411
rect	306	410	307	411
rect	307	410	308	411
rect	308	410	309	411
rect	309	410	310	411
rect	310	410	311	411
rect	311	410	312	411
rect	312	410	313	411
rect	313	410	314	411
rect	314	410	315	411
rect	315	410	316	411
rect	316	410	317	411
rect	317	410	318	411
rect	318	410	319	411
rect	319	410	320	411
rect	321	410	322	411
rect	322	410	323	411
rect	323	410	324	411
rect	324	410	325	411
rect	325	410	326	411
rect	326	410	327	411
rect	327	410	328	411
rect	328	410	329	411
rect	329	410	330	411
rect	330	410	331	411
rect	331	410	332	411
rect	332	410	333	411
rect	0	411	1	412
rect	1	411	2	412
rect	2	411	3	412
rect	3	411	4	412
rect	4	411	5	412
rect	5	411	6	412
rect	7	411	8	412
rect	8	411	9	412
rect	9	411	10	412
rect	10	411	11	412
rect	11	411	12	412
rect	12	411	13	412
rect	14	411	15	412
rect	15	411	16	412
rect	16	411	17	412
rect	17	411	18	412
rect	18	411	19	412
rect	19	411	20	412
rect	21	411	22	412
rect	22	411	23	412
rect	23	411	24	412
rect	24	411	25	412
rect	25	411	26	412
rect	26	411	27	412
rect	28	411	29	412
rect	29	411	30	412
rect	30	411	31	412
rect	31	411	32	412
rect	32	411	33	412
rect	33	411	34	412
rect	35	411	36	412
rect	36	411	37	412
rect	37	411	38	412
rect	38	411	39	412
rect	39	411	40	412
rect	40	411	41	412
rect	42	411	43	412
rect	43	411	44	412
rect	44	411	45	412
rect	45	411	46	412
rect	46	411	47	412
rect	47	411	48	412
rect	49	411	50	412
rect	50	411	51	412
rect	51	411	52	412
rect	52	411	53	412
rect	53	411	54	412
rect	54	411	55	412
rect	56	411	57	412
rect	57	411	58	412
rect	58	411	59	412
rect	59	411	60	412
rect	60	411	61	412
rect	61	411	62	412
rect	62	411	63	412
rect	63	411	64	412
rect	64	411	65	412
rect	65	411	66	412
rect	66	411	67	412
rect	67	411	68	412
rect	68	411	69	412
rect	69	411	70	412
rect	70	411	71	412
rect	71	411	72	412
rect	72	411	73	412
rect	73	411	74	412
rect	74	411	75	412
rect	75	411	76	412
rect	76	411	77	412
rect	77	411	78	412
rect	78	411	79	412
rect	79	411	80	412
rect	80	411	81	412
rect	81	411	82	412
rect	82	411	83	412
rect	83	411	84	412
rect	84	411	85	412
rect	85	411	86	412
rect	86	411	87	412
rect	87	411	88	412
rect	88	411	89	412
rect	90	411	91	412
rect	91	411	92	412
rect	92	411	93	412
rect	93	411	94	412
rect	94	411	95	412
rect	95	411	96	412
rect	96	411	97	412
rect	97	411	98	412
rect	98	411	99	412
rect	99	411	100	412
rect	100	411	101	412
rect	101	411	102	412
rect	102	411	103	412
rect	103	411	104	412
rect	104	411	105	412
rect	105	411	106	412
rect	106	411	107	412
rect	107	411	108	412
rect	108	411	109	412
rect	109	411	110	412
rect	110	411	111	412
rect	111	411	112	412
rect	112	411	113	412
rect	113	411	114	412
rect	114	411	115	412
rect	115	411	116	412
rect	116	411	117	412
rect	117	411	118	412
rect	118	411	119	412
rect	119	411	120	412
rect	120	411	121	412
rect	121	411	122	412
rect	122	411	123	412
rect	123	411	124	412
rect	124	411	125	412
rect	125	411	126	412
rect	126	411	127	412
rect	127	411	128	412
rect	128	411	129	412
rect	129	411	130	412
rect	130	411	131	412
rect	131	411	132	412
rect	132	411	133	412
rect	133	411	134	412
rect	134	411	135	412
rect	135	411	136	412
rect	136	411	137	412
rect	137	411	138	412
rect	139	411	140	412
rect	140	411	141	412
rect	141	411	142	412
rect	142	411	143	412
rect	143	411	144	412
rect	144	411	145	412
rect	145	411	146	412
rect	146	411	147	412
rect	147	411	148	412
rect	148	411	149	412
rect	149	411	150	412
rect	150	411	151	412
rect	151	411	152	412
rect	152	411	153	412
rect	153	411	154	412
rect	155	411	156	412
rect	156	411	157	412
rect	157	411	158	412
rect	158	411	159	412
rect	159	411	160	412
rect	160	411	161	412
rect	162	411	163	412
rect	163	411	164	412
rect	164	411	165	412
rect	165	411	166	412
rect	166	411	167	412
rect	167	411	168	412
rect	169	411	170	412
rect	170	411	171	412
rect	171	411	172	412
rect	172	411	173	412
rect	173	411	174	412
rect	174	411	175	412
rect	176	411	177	412
rect	177	411	178	412
rect	178	411	179	412
rect	179	411	180	412
rect	180	411	181	412
rect	181	411	182	412
rect	183	411	184	412
rect	184	411	185	412
rect	185	411	186	412
rect	186	411	187	412
rect	187	411	188	412
rect	188	411	189	412
rect	190	411	191	412
rect	191	411	192	412
rect	192	411	193	412
rect	193	411	194	412
rect	194	411	195	412
rect	195	411	196	412
rect	196	411	197	412
rect	197	411	198	412
rect	198	411	199	412
rect	199	411	200	412
rect	200	411	201	412
rect	201	411	202	412
rect	202	411	203	412
rect	203	411	204	412
rect	204	411	205	412
rect	205	411	206	412
rect	206	411	207	412
rect	207	411	208	412
rect	208	411	209	412
rect	209	411	210	412
rect	210	411	211	412
rect	211	411	212	412
rect	212	411	213	412
rect	213	411	214	412
rect	214	411	215	412
rect	215	411	216	412
rect	216	411	217	412
rect	217	411	218	412
rect	218	411	219	412
rect	219	411	220	412
rect	220	411	221	412
rect	221	411	222	412
rect	222	411	223	412
rect	223	411	224	412
rect	224	411	225	412
rect	225	411	226	412
rect	226	411	227	412
rect	227	411	228	412
rect	228	411	229	412
rect	229	411	230	412
rect	230	411	231	412
rect	231	411	232	412
rect	232	411	233	412
rect	233	411	234	412
rect	234	411	235	412
rect	235	411	236	412
rect	236	411	237	412
rect	237	411	238	412
rect	238	411	239	412
rect	239	411	240	412
rect	240	411	241	412
rect	241	411	242	412
rect	242	411	243	412
rect	243	411	244	412
rect	244	411	245	412
rect	245	411	246	412
rect	246	411	247	412
rect	247	411	248	412
rect	248	411	249	412
rect	249	411	250	412
rect	250	411	251	412
rect	251	411	252	412
rect	252	411	253	412
rect	253	411	254	412
rect	254	411	255	412
rect	255	411	256	412
rect	256	411	257	412
rect	257	411	258	412
rect	258	411	259	412
rect	259	411	260	412
rect	260	411	261	412
rect	261	411	262	412
rect	262	411	263	412
rect	263	411	264	412
rect	264	411	265	412
rect	265	411	266	412
rect	266	411	267	412
rect	267	411	268	412
rect	268	411	269	412
rect	269	411	270	412
rect	270	411	271	412
rect	271	411	272	412
rect	272	411	273	412
rect	273	411	274	412
rect	274	411	275	412
rect	275	411	276	412
rect	276	411	277	412
rect	277	411	278	412
rect	278	411	279	412
rect	279	411	280	412
rect	280	411	281	412
rect	281	411	282	412
rect	282	411	283	412
rect	283	411	284	412
rect	284	411	285	412
rect	285	411	286	412
rect	286	411	287	412
rect	287	411	288	412
rect	288	411	289	412
rect	289	411	290	412
rect	290	411	291	412
rect	291	411	292	412
rect	292	411	293	412
rect	293	411	294	412
rect	294	411	295	412
rect	296	411	297	412
rect	297	411	298	412
rect	298	411	299	412
rect	299	411	300	412
rect	300	411	301	412
rect	301	411	302	412
rect	302	411	303	412
rect	303	411	304	412
rect	304	411	305	412
rect	305	411	306	412
rect	306	411	307	412
rect	307	411	308	412
rect	308	411	309	412
rect	309	411	310	412
rect	310	411	311	412
rect	311	411	312	412
rect	312	411	313	412
rect	313	411	314	412
rect	314	411	315	412
rect	315	411	316	412
rect	316	411	317	412
rect	317	411	318	412
rect	318	411	319	412
rect	319	411	320	412
rect	321	411	322	412
rect	322	411	323	412
rect	323	411	324	412
rect	324	411	325	412
rect	325	411	326	412
rect	326	411	327	412
rect	327	411	328	412
rect	328	411	329	412
rect	329	411	330	412
rect	330	411	331	412
rect	331	411	332	412
rect	332	411	333	412
rect	0	429	1	430
rect	1	429	2	430
rect	2	429	3	430
rect	3	429	4	430
rect	4	429	5	430
rect	5	429	6	430
rect	7	429	8	430
rect	8	429	9	430
rect	9	429	10	430
rect	10	429	11	430
rect	11	429	12	430
rect	12	429	13	430
rect	14	429	15	430
rect	15	429	16	430
rect	16	429	17	430
rect	17	429	18	430
rect	18	429	19	430
rect	19	429	20	430
rect	21	429	22	430
rect	22	429	23	430
rect	23	429	24	430
rect	24	429	25	430
rect	25	429	26	430
rect	26	429	27	430
rect	28	429	29	430
rect	29	429	30	430
rect	30	429	31	430
rect	31	429	32	430
rect	32	429	33	430
rect	33	429	34	430
rect	35	429	36	430
rect	36	429	37	430
rect	37	429	38	430
rect	38	429	39	430
rect	39	429	40	430
rect	40	429	41	430
rect	42	429	43	430
rect	43	429	44	430
rect	44	429	45	430
rect	45	429	46	430
rect	46	429	47	430
rect	47	429	48	430
rect	49	429	50	430
rect	50	429	51	430
rect	51	429	52	430
rect	52	429	53	430
rect	53	429	54	430
rect	54	429	55	430
rect	56	429	57	430
rect	57	429	58	430
rect	58	429	59	430
rect	59	429	60	430
rect	60	429	61	430
rect	61	429	62	430
rect	63	429	64	430
rect	64	429	65	430
rect	65	429	66	430
rect	66	429	67	430
rect	67	429	68	430
rect	68	429	69	430
rect	70	429	71	430
rect	71	429	72	430
rect	72	429	73	430
rect	73	429	74	430
rect	74	429	75	430
rect	75	429	76	430
rect	76	429	77	430
rect	77	429	78	430
rect	78	429	79	430
rect	79	429	80	430
rect	80	429	81	430
rect	81	429	82	430
rect	82	429	83	430
rect	83	429	84	430
rect	84	429	85	430
rect	85	429	86	430
rect	86	429	87	430
rect	87	429	88	430
rect	88	429	89	430
rect	89	429	90	430
rect	90	429	91	430
rect	91	429	92	430
rect	92	429	93	430
rect	93	429	94	430
rect	94	429	95	430
rect	95	429	96	430
rect	96	429	97	430
rect	97	429	98	430
rect	98	429	99	430
rect	99	429	100	430
rect	100	429	101	430
rect	101	429	102	430
rect	102	429	103	430
rect	103	429	104	430
rect	104	429	105	430
rect	105	429	106	430
rect	106	429	107	430
rect	107	429	108	430
rect	108	429	109	430
rect	109	429	110	430
rect	110	429	111	430
rect	111	429	112	430
rect	112	429	113	430
rect	113	429	114	430
rect	114	429	115	430
rect	115	429	116	430
rect	116	429	117	430
rect	117	429	118	430
rect	119	429	120	430
rect	120	429	121	430
rect	121	429	122	430
rect	122	429	123	430
rect	123	429	124	430
rect	124	429	125	430
rect	126	429	127	430
rect	127	429	128	430
rect	128	429	129	430
rect	129	429	130	430
rect	130	429	131	430
rect	131	429	132	430
rect	133	429	134	430
rect	134	429	135	430
rect	135	429	136	430
rect	136	429	137	430
rect	137	429	138	430
rect	138	429	139	430
rect	140	429	141	430
rect	141	429	142	430
rect	142	429	143	430
rect	143	429	144	430
rect	144	429	145	430
rect	145	429	146	430
rect	147	429	148	430
rect	148	429	149	430
rect	149	429	150	430
rect	150	429	151	430
rect	151	429	152	430
rect	152	429	153	430
rect	154	429	155	430
rect	155	429	156	430
rect	156	429	157	430
rect	157	429	158	430
rect	158	429	159	430
rect	159	429	160	430
rect	161	429	162	430
rect	162	429	163	430
rect	163	429	164	430
rect	164	429	165	430
rect	165	429	166	430
rect	166	429	167	430
rect	168	429	169	430
rect	169	429	170	430
rect	170	429	171	430
rect	171	429	172	430
rect	172	429	173	430
rect	173	429	174	430
rect	175	429	176	430
rect	176	429	177	430
rect	177	429	178	430
rect	178	429	179	430
rect	179	429	180	430
rect	180	429	181	430
rect	182	429	183	430
rect	183	429	184	430
rect	184	429	185	430
rect	185	429	186	430
rect	186	429	187	430
rect	187	429	188	430
rect	189	429	190	430
rect	190	429	191	430
rect	191	429	192	430
rect	192	429	193	430
rect	193	429	194	430
rect	194	429	195	430
rect	195	429	196	430
rect	196	429	197	430
rect	197	429	198	430
rect	198	429	199	430
rect	199	429	200	430
rect	200	429	201	430
rect	201	429	202	430
rect	202	429	203	430
rect	203	429	204	430
rect	204	429	205	430
rect	205	429	206	430
rect	206	429	207	430
rect	207	429	208	430
rect	208	429	209	430
rect	209	429	210	430
rect	210	429	211	430
rect	211	429	212	430
rect	212	429	213	430
rect	214	429	215	430
rect	215	429	216	430
rect	216	429	217	430
rect	217	429	218	430
rect	218	429	219	430
rect	219	429	220	430
rect	220	429	221	430
rect	221	429	222	430
rect	222	429	223	430
rect	223	429	224	430
rect	224	429	225	430
rect	225	429	226	430
rect	226	429	227	430
rect	227	429	228	430
rect	228	429	229	430
rect	230	429	231	430
rect	231	429	232	430
rect	232	429	233	430
rect	233	429	234	430
rect	234	429	235	430
rect	235	429	236	430
rect	236	429	237	430
rect	237	429	238	430
rect	238	429	239	430
rect	239	429	240	430
rect	240	429	241	430
rect	241	429	242	430
rect	242	429	243	430
rect	243	429	244	430
rect	244	429	245	430
rect	246	429	247	430
rect	247	429	248	430
rect	248	429	249	430
rect	249	429	250	430
rect	250	429	251	430
rect	251	429	252	430
rect	252	429	253	430
rect	253	429	254	430
rect	254	429	255	430
rect	255	429	256	430
rect	256	429	257	430
rect	257	429	258	430
rect	258	429	259	430
rect	259	429	260	430
rect	260	429	261	430
rect	261	429	262	430
rect	262	429	263	430
rect	263	429	264	430
rect	264	429	265	430
rect	265	429	266	430
rect	266	429	267	430
rect	267	429	268	430
rect	268	429	269	430
rect	269	429	270	430
rect	270	429	271	430
rect	271	429	272	430
rect	272	429	273	430
rect	274	429	275	430
rect	275	429	276	430
rect	276	429	277	430
rect	277	429	278	430
rect	278	429	279	430
rect	279	429	280	430
rect	280	429	281	430
rect	281	429	282	430
rect	282	429	283	430
rect	0	430	1	431
rect	1	430	2	431
rect	2	430	3	431
rect	3	430	4	431
rect	4	430	5	431
rect	5	430	6	431
rect	7	430	8	431
rect	8	430	9	431
rect	9	430	10	431
rect	10	430	11	431
rect	11	430	12	431
rect	12	430	13	431
rect	14	430	15	431
rect	15	430	16	431
rect	16	430	17	431
rect	17	430	18	431
rect	18	430	19	431
rect	19	430	20	431
rect	21	430	22	431
rect	22	430	23	431
rect	23	430	24	431
rect	24	430	25	431
rect	25	430	26	431
rect	26	430	27	431
rect	28	430	29	431
rect	29	430	30	431
rect	30	430	31	431
rect	31	430	32	431
rect	32	430	33	431
rect	33	430	34	431
rect	35	430	36	431
rect	36	430	37	431
rect	37	430	38	431
rect	38	430	39	431
rect	39	430	40	431
rect	40	430	41	431
rect	42	430	43	431
rect	43	430	44	431
rect	44	430	45	431
rect	45	430	46	431
rect	46	430	47	431
rect	47	430	48	431
rect	49	430	50	431
rect	50	430	51	431
rect	51	430	52	431
rect	52	430	53	431
rect	53	430	54	431
rect	54	430	55	431
rect	56	430	57	431
rect	57	430	58	431
rect	58	430	59	431
rect	59	430	60	431
rect	60	430	61	431
rect	61	430	62	431
rect	63	430	64	431
rect	64	430	65	431
rect	65	430	66	431
rect	66	430	67	431
rect	67	430	68	431
rect	68	430	69	431
rect	70	430	71	431
rect	71	430	72	431
rect	72	430	73	431
rect	73	430	74	431
rect	74	430	75	431
rect	75	430	76	431
rect	76	430	77	431
rect	77	430	78	431
rect	78	430	79	431
rect	79	430	80	431
rect	80	430	81	431
rect	81	430	82	431
rect	82	430	83	431
rect	83	430	84	431
rect	84	430	85	431
rect	85	430	86	431
rect	86	430	87	431
rect	87	430	88	431
rect	88	430	89	431
rect	89	430	90	431
rect	90	430	91	431
rect	91	430	92	431
rect	92	430	93	431
rect	93	430	94	431
rect	94	430	95	431
rect	95	430	96	431
rect	96	430	97	431
rect	97	430	98	431
rect	98	430	99	431
rect	99	430	100	431
rect	100	430	101	431
rect	101	430	102	431
rect	102	430	103	431
rect	103	430	104	431
rect	104	430	105	431
rect	105	430	106	431
rect	106	430	107	431
rect	107	430	108	431
rect	108	430	109	431
rect	109	430	110	431
rect	110	430	111	431
rect	111	430	112	431
rect	112	430	113	431
rect	113	430	114	431
rect	114	430	115	431
rect	115	430	116	431
rect	116	430	117	431
rect	117	430	118	431
rect	119	430	120	431
rect	120	430	121	431
rect	121	430	122	431
rect	122	430	123	431
rect	123	430	124	431
rect	124	430	125	431
rect	126	430	127	431
rect	127	430	128	431
rect	128	430	129	431
rect	129	430	130	431
rect	130	430	131	431
rect	131	430	132	431
rect	133	430	134	431
rect	134	430	135	431
rect	135	430	136	431
rect	136	430	137	431
rect	137	430	138	431
rect	138	430	139	431
rect	140	430	141	431
rect	141	430	142	431
rect	142	430	143	431
rect	143	430	144	431
rect	144	430	145	431
rect	145	430	146	431
rect	147	430	148	431
rect	148	430	149	431
rect	149	430	150	431
rect	150	430	151	431
rect	151	430	152	431
rect	152	430	153	431
rect	154	430	155	431
rect	155	430	156	431
rect	156	430	157	431
rect	157	430	158	431
rect	158	430	159	431
rect	159	430	160	431
rect	161	430	162	431
rect	162	430	163	431
rect	163	430	164	431
rect	164	430	165	431
rect	165	430	166	431
rect	166	430	167	431
rect	168	430	169	431
rect	169	430	170	431
rect	170	430	171	431
rect	171	430	172	431
rect	172	430	173	431
rect	173	430	174	431
rect	175	430	176	431
rect	176	430	177	431
rect	177	430	178	431
rect	178	430	179	431
rect	179	430	180	431
rect	180	430	181	431
rect	182	430	183	431
rect	183	430	184	431
rect	184	430	185	431
rect	185	430	186	431
rect	186	430	187	431
rect	187	430	188	431
rect	189	430	190	431
rect	190	430	191	431
rect	191	430	192	431
rect	192	430	193	431
rect	193	430	194	431
rect	194	430	195	431
rect	195	430	196	431
rect	196	430	197	431
rect	197	430	198	431
rect	198	430	199	431
rect	199	430	200	431
rect	200	430	201	431
rect	201	430	202	431
rect	202	430	203	431
rect	203	430	204	431
rect	204	430	205	431
rect	205	430	206	431
rect	206	430	207	431
rect	207	430	208	431
rect	208	430	209	431
rect	209	430	210	431
rect	210	430	211	431
rect	211	430	212	431
rect	212	430	213	431
rect	214	430	215	431
rect	215	430	216	431
rect	216	430	217	431
rect	217	430	218	431
rect	218	430	219	431
rect	219	430	220	431
rect	220	430	221	431
rect	221	430	222	431
rect	222	430	223	431
rect	223	430	224	431
rect	224	430	225	431
rect	225	430	226	431
rect	226	430	227	431
rect	227	430	228	431
rect	228	430	229	431
rect	230	430	231	431
rect	231	430	232	431
rect	232	430	233	431
rect	233	430	234	431
rect	234	430	235	431
rect	235	430	236	431
rect	236	430	237	431
rect	237	430	238	431
rect	238	430	239	431
rect	239	430	240	431
rect	240	430	241	431
rect	241	430	242	431
rect	242	430	243	431
rect	243	430	244	431
rect	244	430	245	431
rect	246	430	247	431
rect	247	430	248	431
rect	248	430	249	431
rect	249	430	250	431
rect	250	430	251	431
rect	251	430	252	431
rect	252	430	253	431
rect	253	430	254	431
rect	254	430	255	431
rect	255	430	256	431
rect	256	430	257	431
rect	257	430	258	431
rect	258	430	259	431
rect	259	430	260	431
rect	260	430	261	431
rect	261	430	262	431
rect	262	430	263	431
rect	263	430	264	431
rect	264	430	265	431
rect	265	430	266	431
rect	266	430	267	431
rect	267	430	268	431
rect	268	430	269	431
rect	269	430	270	431
rect	270	430	271	431
rect	271	430	272	431
rect	272	430	273	431
rect	274	430	275	431
rect	275	430	276	431
rect	276	430	277	431
rect	277	430	278	431
rect	278	430	279	431
rect	279	430	280	431
rect	280	430	281	431
rect	281	430	282	431
rect	282	430	283	431
rect	0	431	1	432
rect	1	431	2	432
rect	2	431	3	432
rect	3	431	4	432
rect	4	431	5	432
rect	5	431	6	432
rect	7	431	8	432
rect	8	431	9	432
rect	9	431	10	432
rect	10	431	11	432
rect	11	431	12	432
rect	12	431	13	432
rect	14	431	15	432
rect	15	431	16	432
rect	16	431	17	432
rect	17	431	18	432
rect	18	431	19	432
rect	19	431	20	432
rect	21	431	22	432
rect	22	431	23	432
rect	23	431	24	432
rect	24	431	25	432
rect	25	431	26	432
rect	26	431	27	432
rect	28	431	29	432
rect	29	431	30	432
rect	30	431	31	432
rect	31	431	32	432
rect	32	431	33	432
rect	33	431	34	432
rect	35	431	36	432
rect	36	431	37	432
rect	37	431	38	432
rect	38	431	39	432
rect	39	431	40	432
rect	40	431	41	432
rect	42	431	43	432
rect	43	431	44	432
rect	44	431	45	432
rect	45	431	46	432
rect	46	431	47	432
rect	47	431	48	432
rect	49	431	50	432
rect	50	431	51	432
rect	51	431	52	432
rect	52	431	53	432
rect	53	431	54	432
rect	54	431	55	432
rect	56	431	57	432
rect	57	431	58	432
rect	58	431	59	432
rect	59	431	60	432
rect	60	431	61	432
rect	61	431	62	432
rect	63	431	64	432
rect	64	431	65	432
rect	65	431	66	432
rect	66	431	67	432
rect	67	431	68	432
rect	68	431	69	432
rect	70	431	71	432
rect	71	431	72	432
rect	72	431	73	432
rect	73	431	74	432
rect	74	431	75	432
rect	75	431	76	432
rect	76	431	77	432
rect	77	431	78	432
rect	78	431	79	432
rect	79	431	80	432
rect	80	431	81	432
rect	81	431	82	432
rect	82	431	83	432
rect	83	431	84	432
rect	84	431	85	432
rect	85	431	86	432
rect	86	431	87	432
rect	87	431	88	432
rect	88	431	89	432
rect	89	431	90	432
rect	90	431	91	432
rect	91	431	92	432
rect	92	431	93	432
rect	93	431	94	432
rect	94	431	95	432
rect	95	431	96	432
rect	96	431	97	432
rect	97	431	98	432
rect	98	431	99	432
rect	99	431	100	432
rect	100	431	101	432
rect	101	431	102	432
rect	102	431	103	432
rect	103	431	104	432
rect	104	431	105	432
rect	105	431	106	432
rect	106	431	107	432
rect	107	431	108	432
rect	108	431	109	432
rect	109	431	110	432
rect	110	431	111	432
rect	111	431	112	432
rect	112	431	113	432
rect	113	431	114	432
rect	114	431	115	432
rect	115	431	116	432
rect	116	431	117	432
rect	117	431	118	432
rect	119	431	120	432
rect	120	431	121	432
rect	121	431	122	432
rect	122	431	123	432
rect	123	431	124	432
rect	124	431	125	432
rect	126	431	127	432
rect	127	431	128	432
rect	128	431	129	432
rect	129	431	130	432
rect	130	431	131	432
rect	131	431	132	432
rect	133	431	134	432
rect	134	431	135	432
rect	135	431	136	432
rect	136	431	137	432
rect	137	431	138	432
rect	138	431	139	432
rect	140	431	141	432
rect	141	431	142	432
rect	142	431	143	432
rect	143	431	144	432
rect	144	431	145	432
rect	145	431	146	432
rect	147	431	148	432
rect	148	431	149	432
rect	149	431	150	432
rect	150	431	151	432
rect	151	431	152	432
rect	152	431	153	432
rect	154	431	155	432
rect	155	431	156	432
rect	156	431	157	432
rect	157	431	158	432
rect	158	431	159	432
rect	159	431	160	432
rect	161	431	162	432
rect	162	431	163	432
rect	163	431	164	432
rect	164	431	165	432
rect	165	431	166	432
rect	166	431	167	432
rect	168	431	169	432
rect	169	431	170	432
rect	170	431	171	432
rect	171	431	172	432
rect	172	431	173	432
rect	173	431	174	432
rect	175	431	176	432
rect	176	431	177	432
rect	177	431	178	432
rect	178	431	179	432
rect	179	431	180	432
rect	180	431	181	432
rect	182	431	183	432
rect	183	431	184	432
rect	184	431	185	432
rect	185	431	186	432
rect	186	431	187	432
rect	187	431	188	432
rect	189	431	190	432
rect	190	431	191	432
rect	191	431	192	432
rect	192	431	193	432
rect	193	431	194	432
rect	194	431	195	432
rect	195	431	196	432
rect	196	431	197	432
rect	197	431	198	432
rect	198	431	199	432
rect	199	431	200	432
rect	200	431	201	432
rect	201	431	202	432
rect	202	431	203	432
rect	203	431	204	432
rect	204	431	205	432
rect	205	431	206	432
rect	206	431	207	432
rect	207	431	208	432
rect	208	431	209	432
rect	209	431	210	432
rect	210	431	211	432
rect	211	431	212	432
rect	212	431	213	432
rect	214	431	215	432
rect	215	431	216	432
rect	216	431	217	432
rect	217	431	218	432
rect	218	431	219	432
rect	219	431	220	432
rect	220	431	221	432
rect	221	431	222	432
rect	222	431	223	432
rect	223	431	224	432
rect	224	431	225	432
rect	225	431	226	432
rect	226	431	227	432
rect	227	431	228	432
rect	228	431	229	432
rect	230	431	231	432
rect	231	431	232	432
rect	232	431	233	432
rect	233	431	234	432
rect	234	431	235	432
rect	235	431	236	432
rect	236	431	237	432
rect	237	431	238	432
rect	238	431	239	432
rect	239	431	240	432
rect	240	431	241	432
rect	241	431	242	432
rect	242	431	243	432
rect	243	431	244	432
rect	244	431	245	432
rect	246	431	247	432
rect	247	431	248	432
rect	248	431	249	432
rect	249	431	250	432
rect	250	431	251	432
rect	251	431	252	432
rect	252	431	253	432
rect	253	431	254	432
rect	254	431	255	432
rect	255	431	256	432
rect	256	431	257	432
rect	257	431	258	432
rect	258	431	259	432
rect	259	431	260	432
rect	260	431	261	432
rect	261	431	262	432
rect	262	431	263	432
rect	263	431	264	432
rect	264	431	265	432
rect	265	431	266	432
rect	266	431	267	432
rect	267	431	268	432
rect	268	431	269	432
rect	269	431	270	432
rect	270	431	271	432
rect	271	431	272	432
rect	272	431	273	432
rect	274	431	275	432
rect	275	431	276	432
rect	276	431	277	432
rect	277	431	278	432
rect	278	431	279	432
rect	279	431	280	432
rect	280	431	281	432
rect	281	431	282	432
rect	282	431	283	432
rect	0	432	1	433
rect	1	432	2	433
rect	2	432	3	433
rect	3	432	4	433
rect	4	432	5	433
rect	5	432	6	433
rect	7	432	8	433
rect	8	432	9	433
rect	9	432	10	433
rect	10	432	11	433
rect	11	432	12	433
rect	12	432	13	433
rect	14	432	15	433
rect	15	432	16	433
rect	16	432	17	433
rect	17	432	18	433
rect	18	432	19	433
rect	19	432	20	433
rect	21	432	22	433
rect	22	432	23	433
rect	23	432	24	433
rect	24	432	25	433
rect	25	432	26	433
rect	26	432	27	433
rect	28	432	29	433
rect	29	432	30	433
rect	30	432	31	433
rect	31	432	32	433
rect	32	432	33	433
rect	33	432	34	433
rect	35	432	36	433
rect	36	432	37	433
rect	37	432	38	433
rect	38	432	39	433
rect	39	432	40	433
rect	40	432	41	433
rect	42	432	43	433
rect	43	432	44	433
rect	44	432	45	433
rect	45	432	46	433
rect	46	432	47	433
rect	47	432	48	433
rect	49	432	50	433
rect	50	432	51	433
rect	51	432	52	433
rect	52	432	53	433
rect	53	432	54	433
rect	54	432	55	433
rect	56	432	57	433
rect	57	432	58	433
rect	58	432	59	433
rect	59	432	60	433
rect	60	432	61	433
rect	61	432	62	433
rect	63	432	64	433
rect	64	432	65	433
rect	65	432	66	433
rect	66	432	67	433
rect	67	432	68	433
rect	68	432	69	433
rect	70	432	71	433
rect	71	432	72	433
rect	72	432	73	433
rect	73	432	74	433
rect	74	432	75	433
rect	75	432	76	433
rect	76	432	77	433
rect	77	432	78	433
rect	78	432	79	433
rect	79	432	80	433
rect	80	432	81	433
rect	81	432	82	433
rect	82	432	83	433
rect	83	432	84	433
rect	84	432	85	433
rect	85	432	86	433
rect	86	432	87	433
rect	87	432	88	433
rect	88	432	89	433
rect	89	432	90	433
rect	90	432	91	433
rect	91	432	92	433
rect	92	432	93	433
rect	93	432	94	433
rect	94	432	95	433
rect	95	432	96	433
rect	96	432	97	433
rect	97	432	98	433
rect	98	432	99	433
rect	99	432	100	433
rect	100	432	101	433
rect	101	432	102	433
rect	102	432	103	433
rect	103	432	104	433
rect	104	432	105	433
rect	105	432	106	433
rect	106	432	107	433
rect	107	432	108	433
rect	108	432	109	433
rect	109	432	110	433
rect	110	432	111	433
rect	111	432	112	433
rect	112	432	113	433
rect	113	432	114	433
rect	114	432	115	433
rect	115	432	116	433
rect	116	432	117	433
rect	117	432	118	433
rect	119	432	120	433
rect	120	432	121	433
rect	121	432	122	433
rect	122	432	123	433
rect	123	432	124	433
rect	124	432	125	433
rect	126	432	127	433
rect	127	432	128	433
rect	128	432	129	433
rect	129	432	130	433
rect	130	432	131	433
rect	131	432	132	433
rect	133	432	134	433
rect	134	432	135	433
rect	135	432	136	433
rect	136	432	137	433
rect	137	432	138	433
rect	138	432	139	433
rect	140	432	141	433
rect	141	432	142	433
rect	142	432	143	433
rect	143	432	144	433
rect	144	432	145	433
rect	145	432	146	433
rect	147	432	148	433
rect	148	432	149	433
rect	149	432	150	433
rect	150	432	151	433
rect	151	432	152	433
rect	152	432	153	433
rect	154	432	155	433
rect	155	432	156	433
rect	156	432	157	433
rect	157	432	158	433
rect	158	432	159	433
rect	159	432	160	433
rect	161	432	162	433
rect	162	432	163	433
rect	163	432	164	433
rect	164	432	165	433
rect	165	432	166	433
rect	166	432	167	433
rect	168	432	169	433
rect	169	432	170	433
rect	170	432	171	433
rect	171	432	172	433
rect	172	432	173	433
rect	173	432	174	433
rect	175	432	176	433
rect	176	432	177	433
rect	177	432	178	433
rect	178	432	179	433
rect	179	432	180	433
rect	180	432	181	433
rect	182	432	183	433
rect	183	432	184	433
rect	184	432	185	433
rect	185	432	186	433
rect	186	432	187	433
rect	187	432	188	433
rect	189	432	190	433
rect	190	432	191	433
rect	191	432	192	433
rect	192	432	193	433
rect	193	432	194	433
rect	194	432	195	433
rect	195	432	196	433
rect	196	432	197	433
rect	197	432	198	433
rect	198	432	199	433
rect	199	432	200	433
rect	200	432	201	433
rect	201	432	202	433
rect	202	432	203	433
rect	203	432	204	433
rect	204	432	205	433
rect	205	432	206	433
rect	206	432	207	433
rect	207	432	208	433
rect	208	432	209	433
rect	209	432	210	433
rect	210	432	211	433
rect	211	432	212	433
rect	212	432	213	433
rect	214	432	215	433
rect	215	432	216	433
rect	216	432	217	433
rect	217	432	218	433
rect	218	432	219	433
rect	219	432	220	433
rect	220	432	221	433
rect	221	432	222	433
rect	222	432	223	433
rect	223	432	224	433
rect	224	432	225	433
rect	225	432	226	433
rect	226	432	227	433
rect	227	432	228	433
rect	228	432	229	433
rect	230	432	231	433
rect	231	432	232	433
rect	232	432	233	433
rect	233	432	234	433
rect	234	432	235	433
rect	235	432	236	433
rect	236	432	237	433
rect	237	432	238	433
rect	238	432	239	433
rect	239	432	240	433
rect	240	432	241	433
rect	241	432	242	433
rect	242	432	243	433
rect	243	432	244	433
rect	244	432	245	433
rect	246	432	247	433
rect	247	432	248	433
rect	248	432	249	433
rect	249	432	250	433
rect	250	432	251	433
rect	251	432	252	433
rect	252	432	253	433
rect	253	432	254	433
rect	254	432	255	433
rect	255	432	256	433
rect	256	432	257	433
rect	257	432	258	433
rect	258	432	259	433
rect	259	432	260	433
rect	260	432	261	433
rect	261	432	262	433
rect	262	432	263	433
rect	263	432	264	433
rect	264	432	265	433
rect	265	432	266	433
rect	266	432	267	433
rect	267	432	268	433
rect	268	432	269	433
rect	269	432	270	433
rect	270	432	271	433
rect	271	432	272	433
rect	272	432	273	433
rect	274	432	275	433
rect	275	432	276	433
rect	276	432	277	433
rect	277	432	278	433
rect	278	432	279	433
rect	279	432	280	433
rect	280	432	281	433
rect	281	432	282	433
rect	282	432	283	433
rect	0	433	1	434
rect	1	433	2	434
rect	2	433	3	434
rect	3	433	4	434
rect	4	433	5	434
rect	5	433	6	434
rect	7	433	8	434
rect	8	433	9	434
rect	9	433	10	434
rect	10	433	11	434
rect	11	433	12	434
rect	12	433	13	434
rect	14	433	15	434
rect	15	433	16	434
rect	16	433	17	434
rect	17	433	18	434
rect	18	433	19	434
rect	19	433	20	434
rect	21	433	22	434
rect	22	433	23	434
rect	23	433	24	434
rect	24	433	25	434
rect	25	433	26	434
rect	26	433	27	434
rect	28	433	29	434
rect	29	433	30	434
rect	30	433	31	434
rect	31	433	32	434
rect	32	433	33	434
rect	33	433	34	434
rect	35	433	36	434
rect	36	433	37	434
rect	37	433	38	434
rect	38	433	39	434
rect	39	433	40	434
rect	40	433	41	434
rect	42	433	43	434
rect	43	433	44	434
rect	44	433	45	434
rect	45	433	46	434
rect	46	433	47	434
rect	47	433	48	434
rect	49	433	50	434
rect	50	433	51	434
rect	51	433	52	434
rect	52	433	53	434
rect	53	433	54	434
rect	54	433	55	434
rect	56	433	57	434
rect	57	433	58	434
rect	58	433	59	434
rect	59	433	60	434
rect	60	433	61	434
rect	61	433	62	434
rect	63	433	64	434
rect	64	433	65	434
rect	65	433	66	434
rect	66	433	67	434
rect	67	433	68	434
rect	68	433	69	434
rect	70	433	71	434
rect	71	433	72	434
rect	72	433	73	434
rect	73	433	74	434
rect	74	433	75	434
rect	75	433	76	434
rect	76	433	77	434
rect	77	433	78	434
rect	78	433	79	434
rect	79	433	80	434
rect	80	433	81	434
rect	81	433	82	434
rect	82	433	83	434
rect	83	433	84	434
rect	84	433	85	434
rect	85	433	86	434
rect	86	433	87	434
rect	87	433	88	434
rect	88	433	89	434
rect	89	433	90	434
rect	90	433	91	434
rect	91	433	92	434
rect	92	433	93	434
rect	93	433	94	434
rect	94	433	95	434
rect	95	433	96	434
rect	96	433	97	434
rect	97	433	98	434
rect	98	433	99	434
rect	99	433	100	434
rect	100	433	101	434
rect	101	433	102	434
rect	102	433	103	434
rect	103	433	104	434
rect	104	433	105	434
rect	105	433	106	434
rect	106	433	107	434
rect	107	433	108	434
rect	108	433	109	434
rect	109	433	110	434
rect	110	433	111	434
rect	111	433	112	434
rect	112	433	113	434
rect	113	433	114	434
rect	114	433	115	434
rect	115	433	116	434
rect	116	433	117	434
rect	117	433	118	434
rect	119	433	120	434
rect	120	433	121	434
rect	121	433	122	434
rect	122	433	123	434
rect	123	433	124	434
rect	124	433	125	434
rect	126	433	127	434
rect	127	433	128	434
rect	128	433	129	434
rect	129	433	130	434
rect	130	433	131	434
rect	131	433	132	434
rect	133	433	134	434
rect	134	433	135	434
rect	135	433	136	434
rect	136	433	137	434
rect	137	433	138	434
rect	138	433	139	434
rect	140	433	141	434
rect	141	433	142	434
rect	142	433	143	434
rect	143	433	144	434
rect	144	433	145	434
rect	145	433	146	434
rect	147	433	148	434
rect	148	433	149	434
rect	149	433	150	434
rect	150	433	151	434
rect	151	433	152	434
rect	152	433	153	434
rect	154	433	155	434
rect	155	433	156	434
rect	156	433	157	434
rect	157	433	158	434
rect	158	433	159	434
rect	159	433	160	434
rect	161	433	162	434
rect	162	433	163	434
rect	163	433	164	434
rect	164	433	165	434
rect	165	433	166	434
rect	166	433	167	434
rect	168	433	169	434
rect	169	433	170	434
rect	170	433	171	434
rect	171	433	172	434
rect	172	433	173	434
rect	173	433	174	434
rect	175	433	176	434
rect	176	433	177	434
rect	177	433	178	434
rect	178	433	179	434
rect	179	433	180	434
rect	180	433	181	434
rect	182	433	183	434
rect	183	433	184	434
rect	184	433	185	434
rect	185	433	186	434
rect	186	433	187	434
rect	187	433	188	434
rect	189	433	190	434
rect	190	433	191	434
rect	191	433	192	434
rect	192	433	193	434
rect	193	433	194	434
rect	194	433	195	434
rect	195	433	196	434
rect	196	433	197	434
rect	197	433	198	434
rect	198	433	199	434
rect	199	433	200	434
rect	200	433	201	434
rect	201	433	202	434
rect	202	433	203	434
rect	203	433	204	434
rect	204	433	205	434
rect	205	433	206	434
rect	206	433	207	434
rect	207	433	208	434
rect	208	433	209	434
rect	209	433	210	434
rect	210	433	211	434
rect	211	433	212	434
rect	212	433	213	434
rect	214	433	215	434
rect	215	433	216	434
rect	216	433	217	434
rect	217	433	218	434
rect	218	433	219	434
rect	219	433	220	434
rect	220	433	221	434
rect	221	433	222	434
rect	222	433	223	434
rect	223	433	224	434
rect	224	433	225	434
rect	225	433	226	434
rect	226	433	227	434
rect	227	433	228	434
rect	228	433	229	434
rect	230	433	231	434
rect	231	433	232	434
rect	232	433	233	434
rect	233	433	234	434
rect	234	433	235	434
rect	235	433	236	434
rect	236	433	237	434
rect	237	433	238	434
rect	238	433	239	434
rect	239	433	240	434
rect	240	433	241	434
rect	241	433	242	434
rect	242	433	243	434
rect	243	433	244	434
rect	244	433	245	434
rect	246	433	247	434
rect	247	433	248	434
rect	248	433	249	434
rect	249	433	250	434
rect	250	433	251	434
rect	251	433	252	434
rect	252	433	253	434
rect	253	433	254	434
rect	254	433	255	434
rect	255	433	256	434
rect	256	433	257	434
rect	257	433	258	434
rect	258	433	259	434
rect	259	433	260	434
rect	260	433	261	434
rect	261	433	262	434
rect	262	433	263	434
rect	263	433	264	434
rect	264	433	265	434
rect	265	433	266	434
rect	266	433	267	434
rect	267	433	268	434
rect	268	433	269	434
rect	269	433	270	434
rect	270	433	271	434
rect	271	433	272	434
rect	272	433	273	434
rect	274	433	275	434
rect	275	433	276	434
rect	276	433	277	434
rect	277	433	278	434
rect	278	433	279	434
rect	279	433	280	434
rect	280	433	281	434
rect	281	433	282	434
rect	282	433	283	434
rect	0	434	1	435
rect	1	434	2	435
rect	2	434	3	435
rect	3	434	4	435
rect	4	434	5	435
rect	5	434	6	435
rect	7	434	8	435
rect	8	434	9	435
rect	9	434	10	435
rect	10	434	11	435
rect	11	434	12	435
rect	12	434	13	435
rect	14	434	15	435
rect	15	434	16	435
rect	16	434	17	435
rect	17	434	18	435
rect	18	434	19	435
rect	19	434	20	435
rect	21	434	22	435
rect	22	434	23	435
rect	23	434	24	435
rect	24	434	25	435
rect	25	434	26	435
rect	26	434	27	435
rect	28	434	29	435
rect	29	434	30	435
rect	30	434	31	435
rect	31	434	32	435
rect	32	434	33	435
rect	33	434	34	435
rect	35	434	36	435
rect	36	434	37	435
rect	37	434	38	435
rect	38	434	39	435
rect	39	434	40	435
rect	40	434	41	435
rect	42	434	43	435
rect	43	434	44	435
rect	44	434	45	435
rect	45	434	46	435
rect	46	434	47	435
rect	47	434	48	435
rect	49	434	50	435
rect	50	434	51	435
rect	51	434	52	435
rect	52	434	53	435
rect	53	434	54	435
rect	54	434	55	435
rect	56	434	57	435
rect	57	434	58	435
rect	58	434	59	435
rect	59	434	60	435
rect	60	434	61	435
rect	61	434	62	435
rect	63	434	64	435
rect	64	434	65	435
rect	65	434	66	435
rect	66	434	67	435
rect	67	434	68	435
rect	68	434	69	435
rect	70	434	71	435
rect	71	434	72	435
rect	72	434	73	435
rect	73	434	74	435
rect	74	434	75	435
rect	75	434	76	435
rect	76	434	77	435
rect	77	434	78	435
rect	78	434	79	435
rect	79	434	80	435
rect	80	434	81	435
rect	81	434	82	435
rect	82	434	83	435
rect	83	434	84	435
rect	84	434	85	435
rect	85	434	86	435
rect	86	434	87	435
rect	87	434	88	435
rect	88	434	89	435
rect	89	434	90	435
rect	90	434	91	435
rect	91	434	92	435
rect	92	434	93	435
rect	93	434	94	435
rect	94	434	95	435
rect	95	434	96	435
rect	96	434	97	435
rect	97	434	98	435
rect	98	434	99	435
rect	99	434	100	435
rect	100	434	101	435
rect	101	434	102	435
rect	102	434	103	435
rect	103	434	104	435
rect	104	434	105	435
rect	105	434	106	435
rect	106	434	107	435
rect	107	434	108	435
rect	108	434	109	435
rect	109	434	110	435
rect	110	434	111	435
rect	111	434	112	435
rect	112	434	113	435
rect	113	434	114	435
rect	114	434	115	435
rect	115	434	116	435
rect	116	434	117	435
rect	117	434	118	435
rect	119	434	120	435
rect	120	434	121	435
rect	121	434	122	435
rect	122	434	123	435
rect	123	434	124	435
rect	124	434	125	435
rect	126	434	127	435
rect	127	434	128	435
rect	128	434	129	435
rect	129	434	130	435
rect	130	434	131	435
rect	131	434	132	435
rect	133	434	134	435
rect	134	434	135	435
rect	135	434	136	435
rect	136	434	137	435
rect	137	434	138	435
rect	138	434	139	435
rect	140	434	141	435
rect	141	434	142	435
rect	142	434	143	435
rect	143	434	144	435
rect	144	434	145	435
rect	145	434	146	435
rect	147	434	148	435
rect	148	434	149	435
rect	149	434	150	435
rect	150	434	151	435
rect	151	434	152	435
rect	152	434	153	435
rect	154	434	155	435
rect	155	434	156	435
rect	156	434	157	435
rect	157	434	158	435
rect	158	434	159	435
rect	159	434	160	435
rect	161	434	162	435
rect	162	434	163	435
rect	163	434	164	435
rect	164	434	165	435
rect	165	434	166	435
rect	166	434	167	435
rect	168	434	169	435
rect	169	434	170	435
rect	170	434	171	435
rect	171	434	172	435
rect	172	434	173	435
rect	173	434	174	435
rect	175	434	176	435
rect	176	434	177	435
rect	177	434	178	435
rect	178	434	179	435
rect	179	434	180	435
rect	180	434	181	435
rect	182	434	183	435
rect	183	434	184	435
rect	184	434	185	435
rect	185	434	186	435
rect	186	434	187	435
rect	187	434	188	435
rect	189	434	190	435
rect	190	434	191	435
rect	191	434	192	435
rect	192	434	193	435
rect	193	434	194	435
rect	194	434	195	435
rect	195	434	196	435
rect	196	434	197	435
rect	197	434	198	435
rect	198	434	199	435
rect	199	434	200	435
rect	200	434	201	435
rect	201	434	202	435
rect	202	434	203	435
rect	203	434	204	435
rect	204	434	205	435
rect	205	434	206	435
rect	206	434	207	435
rect	207	434	208	435
rect	208	434	209	435
rect	209	434	210	435
rect	210	434	211	435
rect	211	434	212	435
rect	212	434	213	435
rect	214	434	215	435
rect	215	434	216	435
rect	216	434	217	435
rect	217	434	218	435
rect	218	434	219	435
rect	219	434	220	435
rect	220	434	221	435
rect	221	434	222	435
rect	222	434	223	435
rect	223	434	224	435
rect	224	434	225	435
rect	225	434	226	435
rect	226	434	227	435
rect	227	434	228	435
rect	228	434	229	435
rect	230	434	231	435
rect	231	434	232	435
rect	232	434	233	435
rect	233	434	234	435
rect	234	434	235	435
rect	235	434	236	435
rect	236	434	237	435
rect	237	434	238	435
rect	238	434	239	435
rect	239	434	240	435
rect	240	434	241	435
rect	241	434	242	435
rect	242	434	243	435
rect	243	434	244	435
rect	244	434	245	435
rect	246	434	247	435
rect	247	434	248	435
rect	248	434	249	435
rect	249	434	250	435
rect	250	434	251	435
rect	251	434	252	435
rect	252	434	253	435
rect	253	434	254	435
rect	254	434	255	435
rect	255	434	256	435
rect	256	434	257	435
rect	257	434	258	435
rect	258	434	259	435
rect	259	434	260	435
rect	260	434	261	435
rect	261	434	262	435
rect	262	434	263	435
rect	263	434	264	435
rect	264	434	265	435
rect	265	434	266	435
rect	266	434	267	435
rect	267	434	268	435
rect	268	434	269	435
rect	269	434	270	435
rect	270	434	271	435
rect	271	434	272	435
rect	272	434	273	435
rect	274	434	275	435
rect	275	434	276	435
rect	276	434	277	435
rect	277	434	278	435
rect	278	434	279	435
rect	279	434	280	435
rect	280	434	281	435
rect	281	434	282	435
rect	282	434	283	435
rect	0	446	1	447
rect	1	446	2	447
rect	2	446	3	447
rect	3	446	4	447
rect	4	446	5	447
rect	5	446	6	447
rect	7	446	8	447
rect	8	446	9	447
rect	9	446	10	447
rect	10	446	11	447
rect	11	446	12	447
rect	12	446	13	447
rect	14	446	15	447
rect	15	446	16	447
rect	16	446	17	447
rect	17	446	18	447
rect	18	446	19	447
rect	19	446	20	447
rect	21	446	22	447
rect	22	446	23	447
rect	23	446	24	447
rect	24	446	25	447
rect	25	446	26	447
rect	26	446	27	447
rect	28	446	29	447
rect	29	446	30	447
rect	30	446	31	447
rect	31	446	32	447
rect	32	446	33	447
rect	33	446	34	447
rect	35	446	36	447
rect	36	446	37	447
rect	37	446	38	447
rect	38	446	39	447
rect	39	446	40	447
rect	40	446	41	447
rect	42	446	43	447
rect	43	446	44	447
rect	44	446	45	447
rect	45	446	46	447
rect	46	446	47	447
rect	47	446	48	447
rect	49	446	50	447
rect	50	446	51	447
rect	51	446	52	447
rect	52	446	53	447
rect	53	446	54	447
rect	54	446	55	447
rect	56	446	57	447
rect	57	446	58	447
rect	58	446	59	447
rect	59	446	60	447
rect	60	446	61	447
rect	61	446	62	447
rect	63	446	64	447
rect	64	446	65	447
rect	65	446	66	447
rect	66	446	67	447
rect	67	446	68	447
rect	68	446	69	447
rect	70	446	71	447
rect	71	446	72	447
rect	72	446	73	447
rect	73	446	74	447
rect	74	446	75	447
rect	75	446	76	447
rect	77	446	78	447
rect	78	446	79	447
rect	79	446	80	447
rect	80	446	81	447
rect	81	446	82	447
rect	82	446	83	447
rect	84	446	85	447
rect	85	446	86	447
rect	86	446	87	447
rect	87	446	88	447
rect	88	446	89	447
rect	89	446	90	447
rect	91	446	92	447
rect	92	446	93	447
rect	93	446	94	447
rect	94	446	95	447
rect	95	446	96	447
rect	96	446	97	447
rect	97	446	98	447
rect	98	446	99	447
rect	99	446	100	447
rect	100	446	101	447
rect	101	446	102	447
rect	102	446	103	447
rect	103	446	104	447
rect	104	446	105	447
rect	105	446	106	447
rect	106	446	107	447
rect	107	446	108	447
rect	108	446	109	447
rect	110	446	111	447
rect	111	446	112	447
rect	112	446	113	447
rect	113	446	114	447
rect	114	446	115	447
rect	115	446	116	447
rect	117	446	118	447
rect	118	446	119	447
rect	119	446	120	447
rect	120	446	121	447
rect	121	446	122	447
rect	122	446	123	447
rect	124	446	125	447
rect	125	446	126	447
rect	126	446	127	447
rect	127	446	128	447
rect	128	446	129	447
rect	129	446	130	447
rect	131	446	132	447
rect	132	446	133	447
rect	133	446	134	447
rect	134	446	135	447
rect	135	446	136	447
rect	136	446	137	447
rect	138	446	139	447
rect	139	446	140	447
rect	140	446	141	447
rect	141	446	142	447
rect	142	446	143	447
rect	143	446	144	447
rect	145	446	146	447
rect	146	446	147	447
rect	147	446	148	447
rect	148	446	149	447
rect	149	446	150	447
rect	150	446	151	447
rect	152	446	153	447
rect	153	446	154	447
rect	154	446	155	447
rect	155	446	156	447
rect	156	446	157	447
rect	157	446	158	447
rect	159	446	160	447
rect	160	446	161	447
rect	161	446	162	447
rect	162	446	163	447
rect	163	446	164	447
rect	164	446	165	447
rect	166	446	167	447
rect	167	446	168	447
rect	168	446	169	447
rect	169	446	170	447
rect	170	446	171	447
rect	171	446	172	447
rect	0	447	1	448
rect	1	447	2	448
rect	2	447	3	448
rect	3	447	4	448
rect	4	447	5	448
rect	5	447	6	448
rect	7	447	8	448
rect	8	447	9	448
rect	9	447	10	448
rect	10	447	11	448
rect	11	447	12	448
rect	12	447	13	448
rect	14	447	15	448
rect	15	447	16	448
rect	16	447	17	448
rect	17	447	18	448
rect	18	447	19	448
rect	19	447	20	448
rect	21	447	22	448
rect	22	447	23	448
rect	23	447	24	448
rect	24	447	25	448
rect	25	447	26	448
rect	26	447	27	448
rect	28	447	29	448
rect	29	447	30	448
rect	30	447	31	448
rect	31	447	32	448
rect	32	447	33	448
rect	33	447	34	448
rect	35	447	36	448
rect	36	447	37	448
rect	37	447	38	448
rect	38	447	39	448
rect	39	447	40	448
rect	40	447	41	448
rect	42	447	43	448
rect	43	447	44	448
rect	44	447	45	448
rect	45	447	46	448
rect	46	447	47	448
rect	47	447	48	448
rect	49	447	50	448
rect	50	447	51	448
rect	51	447	52	448
rect	52	447	53	448
rect	53	447	54	448
rect	54	447	55	448
rect	56	447	57	448
rect	57	447	58	448
rect	58	447	59	448
rect	59	447	60	448
rect	60	447	61	448
rect	61	447	62	448
rect	63	447	64	448
rect	64	447	65	448
rect	65	447	66	448
rect	66	447	67	448
rect	67	447	68	448
rect	68	447	69	448
rect	70	447	71	448
rect	71	447	72	448
rect	72	447	73	448
rect	73	447	74	448
rect	74	447	75	448
rect	75	447	76	448
rect	77	447	78	448
rect	78	447	79	448
rect	79	447	80	448
rect	80	447	81	448
rect	81	447	82	448
rect	82	447	83	448
rect	84	447	85	448
rect	85	447	86	448
rect	86	447	87	448
rect	87	447	88	448
rect	88	447	89	448
rect	89	447	90	448
rect	91	447	92	448
rect	92	447	93	448
rect	93	447	94	448
rect	94	447	95	448
rect	95	447	96	448
rect	96	447	97	448
rect	97	447	98	448
rect	98	447	99	448
rect	99	447	100	448
rect	100	447	101	448
rect	101	447	102	448
rect	102	447	103	448
rect	103	447	104	448
rect	104	447	105	448
rect	105	447	106	448
rect	106	447	107	448
rect	107	447	108	448
rect	108	447	109	448
rect	110	447	111	448
rect	111	447	112	448
rect	112	447	113	448
rect	113	447	114	448
rect	114	447	115	448
rect	115	447	116	448
rect	117	447	118	448
rect	118	447	119	448
rect	119	447	120	448
rect	120	447	121	448
rect	121	447	122	448
rect	122	447	123	448
rect	124	447	125	448
rect	125	447	126	448
rect	126	447	127	448
rect	127	447	128	448
rect	128	447	129	448
rect	129	447	130	448
rect	131	447	132	448
rect	132	447	133	448
rect	133	447	134	448
rect	134	447	135	448
rect	135	447	136	448
rect	136	447	137	448
rect	138	447	139	448
rect	139	447	140	448
rect	140	447	141	448
rect	141	447	142	448
rect	142	447	143	448
rect	143	447	144	448
rect	145	447	146	448
rect	146	447	147	448
rect	147	447	148	448
rect	148	447	149	448
rect	149	447	150	448
rect	150	447	151	448
rect	152	447	153	448
rect	153	447	154	448
rect	154	447	155	448
rect	155	447	156	448
rect	156	447	157	448
rect	157	447	158	448
rect	159	447	160	448
rect	160	447	161	448
rect	161	447	162	448
rect	162	447	163	448
rect	163	447	164	448
rect	164	447	165	448
rect	166	447	167	448
rect	167	447	168	448
rect	168	447	169	448
rect	169	447	170	448
rect	170	447	171	448
rect	171	447	172	448
rect	0	448	1	449
rect	1	448	2	449
rect	2	448	3	449
rect	3	448	4	449
rect	4	448	5	449
rect	5	448	6	449
rect	7	448	8	449
rect	8	448	9	449
rect	9	448	10	449
rect	10	448	11	449
rect	11	448	12	449
rect	12	448	13	449
rect	14	448	15	449
rect	15	448	16	449
rect	16	448	17	449
rect	17	448	18	449
rect	18	448	19	449
rect	19	448	20	449
rect	21	448	22	449
rect	22	448	23	449
rect	23	448	24	449
rect	24	448	25	449
rect	25	448	26	449
rect	26	448	27	449
rect	28	448	29	449
rect	29	448	30	449
rect	30	448	31	449
rect	31	448	32	449
rect	32	448	33	449
rect	33	448	34	449
rect	35	448	36	449
rect	36	448	37	449
rect	37	448	38	449
rect	38	448	39	449
rect	39	448	40	449
rect	40	448	41	449
rect	42	448	43	449
rect	43	448	44	449
rect	44	448	45	449
rect	45	448	46	449
rect	46	448	47	449
rect	47	448	48	449
rect	49	448	50	449
rect	50	448	51	449
rect	51	448	52	449
rect	52	448	53	449
rect	53	448	54	449
rect	54	448	55	449
rect	56	448	57	449
rect	57	448	58	449
rect	58	448	59	449
rect	59	448	60	449
rect	60	448	61	449
rect	61	448	62	449
rect	63	448	64	449
rect	64	448	65	449
rect	65	448	66	449
rect	66	448	67	449
rect	67	448	68	449
rect	68	448	69	449
rect	70	448	71	449
rect	71	448	72	449
rect	72	448	73	449
rect	73	448	74	449
rect	74	448	75	449
rect	75	448	76	449
rect	77	448	78	449
rect	78	448	79	449
rect	79	448	80	449
rect	80	448	81	449
rect	81	448	82	449
rect	82	448	83	449
rect	84	448	85	449
rect	85	448	86	449
rect	86	448	87	449
rect	87	448	88	449
rect	88	448	89	449
rect	89	448	90	449
rect	91	448	92	449
rect	92	448	93	449
rect	93	448	94	449
rect	94	448	95	449
rect	95	448	96	449
rect	96	448	97	449
rect	97	448	98	449
rect	98	448	99	449
rect	99	448	100	449
rect	100	448	101	449
rect	101	448	102	449
rect	102	448	103	449
rect	103	448	104	449
rect	104	448	105	449
rect	105	448	106	449
rect	106	448	107	449
rect	107	448	108	449
rect	108	448	109	449
rect	110	448	111	449
rect	111	448	112	449
rect	112	448	113	449
rect	113	448	114	449
rect	114	448	115	449
rect	115	448	116	449
rect	117	448	118	449
rect	118	448	119	449
rect	119	448	120	449
rect	120	448	121	449
rect	121	448	122	449
rect	122	448	123	449
rect	124	448	125	449
rect	125	448	126	449
rect	126	448	127	449
rect	127	448	128	449
rect	128	448	129	449
rect	129	448	130	449
rect	131	448	132	449
rect	132	448	133	449
rect	133	448	134	449
rect	134	448	135	449
rect	135	448	136	449
rect	136	448	137	449
rect	138	448	139	449
rect	139	448	140	449
rect	140	448	141	449
rect	141	448	142	449
rect	142	448	143	449
rect	143	448	144	449
rect	145	448	146	449
rect	146	448	147	449
rect	147	448	148	449
rect	148	448	149	449
rect	149	448	150	449
rect	150	448	151	449
rect	152	448	153	449
rect	153	448	154	449
rect	154	448	155	449
rect	155	448	156	449
rect	156	448	157	449
rect	157	448	158	449
rect	159	448	160	449
rect	160	448	161	449
rect	161	448	162	449
rect	162	448	163	449
rect	163	448	164	449
rect	164	448	165	449
rect	166	448	167	449
rect	167	448	168	449
rect	168	448	169	449
rect	169	448	170	449
rect	170	448	171	449
rect	171	448	172	449
rect	0	449	1	450
rect	1	449	2	450
rect	2	449	3	450
rect	3	449	4	450
rect	4	449	5	450
rect	5	449	6	450
rect	7	449	8	450
rect	8	449	9	450
rect	9	449	10	450
rect	10	449	11	450
rect	11	449	12	450
rect	12	449	13	450
rect	14	449	15	450
rect	15	449	16	450
rect	16	449	17	450
rect	17	449	18	450
rect	18	449	19	450
rect	19	449	20	450
rect	21	449	22	450
rect	22	449	23	450
rect	23	449	24	450
rect	24	449	25	450
rect	25	449	26	450
rect	26	449	27	450
rect	28	449	29	450
rect	29	449	30	450
rect	30	449	31	450
rect	31	449	32	450
rect	32	449	33	450
rect	33	449	34	450
rect	35	449	36	450
rect	36	449	37	450
rect	37	449	38	450
rect	38	449	39	450
rect	39	449	40	450
rect	40	449	41	450
rect	42	449	43	450
rect	43	449	44	450
rect	44	449	45	450
rect	45	449	46	450
rect	46	449	47	450
rect	47	449	48	450
rect	49	449	50	450
rect	50	449	51	450
rect	51	449	52	450
rect	52	449	53	450
rect	53	449	54	450
rect	54	449	55	450
rect	56	449	57	450
rect	57	449	58	450
rect	58	449	59	450
rect	59	449	60	450
rect	60	449	61	450
rect	61	449	62	450
rect	63	449	64	450
rect	64	449	65	450
rect	65	449	66	450
rect	66	449	67	450
rect	67	449	68	450
rect	68	449	69	450
rect	70	449	71	450
rect	71	449	72	450
rect	72	449	73	450
rect	73	449	74	450
rect	74	449	75	450
rect	75	449	76	450
rect	77	449	78	450
rect	78	449	79	450
rect	79	449	80	450
rect	80	449	81	450
rect	81	449	82	450
rect	82	449	83	450
rect	84	449	85	450
rect	85	449	86	450
rect	86	449	87	450
rect	87	449	88	450
rect	88	449	89	450
rect	89	449	90	450
rect	91	449	92	450
rect	92	449	93	450
rect	93	449	94	450
rect	94	449	95	450
rect	95	449	96	450
rect	96	449	97	450
rect	97	449	98	450
rect	98	449	99	450
rect	99	449	100	450
rect	100	449	101	450
rect	101	449	102	450
rect	102	449	103	450
rect	103	449	104	450
rect	104	449	105	450
rect	105	449	106	450
rect	106	449	107	450
rect	107	449	108	450
rect	108	449	109	450
rect	110	449	111	450
rect	111	449	112	450
rect	112	449	113	450
rect	113	449	114	450
rect	114	449	115	450
rect	115	449	116	450
rect	117	449	118	450
rect	118	449	119	450
rect	119	449	120	450
rect	120	449	121	450
rect	121	449	122	450
rect	122	449	123	450
rect	124	449	125	450
rect	125	449	126	450
rect	126	449	127	450
rect	127	449	128	450
rect	128	449	129	450
rect	129	449	130	450
rect	131	449	132	450
rect	132	449	133	450
rect	133	449	134	450
rect	134	449	135	450
rect	135	449	136	450
rect	136	449	137	450
rect	138	449	139	450
rect	139	449	140	450
rect	140	449	141	450
rect	141	449	142	450
rect	142	449	143	450
rect	143	449	144	450
rect	145	449	146	450
rect	146	449	147	450
rect	147	449	148	450
rect	148	449	149	450
rect	149	449	150	450
rect	150	449	151	450
rect	152	449	153	450
rect	153	449	154	450
rect	154	449	155	450
rect	155	449	156	450
rect	156	449	157	450
rect	157	449	158	450
rect	159	449	160	450
rect	160	449	161	450
rect	161	449	162	450
rect	162	449	163	450
rect	163	449	164	450
rect	164	449	165	450
rect	166	449	167	450
rect	167	449	168	450
rect	168	449	169	450
rect	169	449	170	450
rect	170	449	171	450
rect	171	449	172	450
rect	0	450	1	451
rect	1	450	2	451
rect	2	450	3	451
rect	3	450	4	451
rect	4	450	5	451
rect	5	450	6	451
rect	7	450	8	451
rect	8	450	9	451
rect	9	450	10	451
rect	10	450	11	451
rect	11	450	12	451
rect	12	450	13	451
rect	14	450	15	451
rect	15	450	16	451
rect	16	450	17	451
rect	17	450	18	451
rect	18	450	19	451
rect	19	450	20	451
rect	21	450	22	451
rect	22	450	23	451
rect	23	450	24	451
rect	24	450	25	451
rect	25	450	26	451
rect	26	450	27	451
rect	28	450	29	451
rect	29	450	30	451
rect	30	450	31	451
rect	31	450	32	451
rect	32	450	33	451
rect	33	450	34	451
rect	35	450	36	451
rect	36	450	37	451
rect	37	450	38	451
rect	38	450	39	451
rect	39	450	40	451
rect	40	450	41	451
rect	42	450	43	451
rect	43	450	44	451
rect	44	450	45	451
rect	45	450	46	451
rect	46	450	47	451
rect	47	450	48	451
rect	49	450	50	451
rect	50	450	51	451
rect	51	450	52	451
rect	52	450	53	451
rect	53	450	54	451
rect	54	450	55	451
rect	56	450	57	451
rect	57	450	58	451
rect	58	450	59	451
rect	59	450	60	451
rect	60	450	61	451
rect	61	450	62	451
rect	63	450	64	451
rect	64	450	65	451
rect	65	450	66	451
rect	66	450	67	451
rect	67	450	68	451
rect	68	450	69	451
rect	70	450	71	451
rect	71	450	72	451
rect	72	450	73	451
rect	73	450	74	451
rect	74	450	75	451
rect	75	450	76	451
rect	77	450	78	451
rect	78	450	79	451
rect	79	450	80	451
rect	80	450	81	451
rect	81	450	82	451
rect	82	450	83	451
rect	84	450	85	451
rect	85	450	86	451
rect	86	450	87	451
rect	87	450	88	451
rect	88	450	89	451
rect	89	450	90	451
rect	91	450	92	451
rect	92	450	93	451
rect	93	450	94	451
rect	94	450	95	451
rect	95	450	96	451
rect	96	450	97	451
rect	97	450	98	451
rect	98	450	99	451
rect	99	450	100	451
rect	100	450	101	451
rect	101	450	102	451
rect	102	450	103	451
rect	103	450	104	451
rect	104	450	105	451
rect	105	450	106	451
rect	106	450	107	451
rect	107	450	108	451
rect	108	450	109	451
rect	110	450	111	451
rect	111	450	112	451
rect	112	450	113	451
rect	113	450	114	451
rect	114	450	115	451
rect	115	450	116	451
rect	117	450	118	451
rect	118	450	119	451
rect	119	450	120	451
rect	120	450	121	451
rect	121	450	122	451
rect	122	450	123	451
rect	124	450	125	451
rect	125	450	126	451
rect	126	450	127	451
rect	127	450	128	451
rect	128	450	129	451
rect	129	450	130	451
rect	131	450	132	451
rect	132	450	133	451
rect	133	450	134	451
rect	134	450	135	451
rect	135	450	136	451
rect	136	450	137	451
rect	138	450	139	451
rect	139	450	140	451
rect	140	450	141	451
rect	141	450	142	451
rect	142	450	143	451
rect	143	450	144	451
rect	145	450	146	451
rect	146	450	147	451
rect	147	450	148	451
rect	148	450	149	451
rect	149	450	150	451
rect	150	450	151	451
rect	152	450	153	451
rect	153	450	154	451
rect	154	450	155	451
rect	155	450	156	451
rect	156	450	157	451
rect	157	450	158	451
rect	159	450	160	451
rect	160	450	161	451
rect	161	450	162	451
rect	162	450	163	451
rect	163	450	164	451
rect	164	450	165	451
rect	166	450	167	451
rect	167	450	168	451
rect	168	450	169	451
rect	169	450	170	451
rect	170	450	171	451
rect	171	450	172	451
rect	0	451	1	452
rect	1	451	2	452
rect	2	451	3	452
rect	3	451	4	452
rect	4	451	5	452
rect	5	451	6	452
rect	7	451	8	452
rect	8	451	9	452
rect	9	451	10	452
rect	10	451	11	452
rect	11	451	12	452
rect	12	451	13	452
rect	14	451	15	452
rect	15	451	16	452
rect	16	451	17	452
rect	17	451	18	452
rect	18	451	19	452
rect	19	451	20	452
rect	21	451	22	452
rect	22	451	23	452
rect	23	451	24	452
rect	24	451	25	452
rect	25	451	26	452
rect	26	451	27	452
rect	28	451	29	452
rect	29	451	30	452
rect	30	451	31	452
rect	31	451	32	452
rect	32	451	33	452
rect	33	451	34	452
rect	35	451	36	452
rect	36	451	37	452
rect	37	451	38	452
rect	38	451	39	452
rect	39	451	40	452
rect	40	451	41	452
rect	42	451	43	452
rect	43	451	44	452
rect	44	451	45	452
rect	45	451	46	452
rect	46	451	47	452
rect	47	451	48	452
rect	49	451	50	452
rect	50	451	51	452
rect	51	451	52	452
rect	52	451	53	452
rect	53	451	54	452
rect	54	451	55	452
rect	56	451	57	452
rect	57	451	58	452
rect	58	451	59	452
rect	59	451	60	452
rect	60	451	61	452
rect	61	451	62	452
rect	63	451	64	452
rect	64	451	65	452
rect	65	451	66	452
rect	66	451	67	452
rect	67	451	68	452
rect	68	451	69	452
rect	70	451	71	452
rect	71	451	72	452
rect	72	451	73	452
rect	73	451	74	452
rect	74	451	75	452
rect	75	451	76	452
rect	77	451	78	452
rect	78	451	79	452
rect	79	451	80	452
rect	80	451	81	452
rect	81	451	82	452
rect	82	451	83	452
rect	84	451	85	452
rect	85	451	86	452
rect	86	451	87	452
rect	87	451	88	452
rect	88	451	89	452
rect	89	451	90	452
rect	91	451	92	452
rect	92	451	93	452
rect	93	451	94	452
rect	94	451	95	452
rect	95	451	96	452
rect	96	451	97	452
rect	97	451	98	452
rect	98	451	99	452
rect	99	451	100	452
rect	100	451	101	452
rect	101	451	102	452
rect	102	451	103	452
rect	103	451	104	452
rect	104	451	105	452
rect	105	451	106	452
rect	106	451	107	452
rect	107	451	108	452
rect	108	451	109	452
rect	110	451	111	452
rect	111	451	112	452
rect	112	451	113	452
rect	113	451	114	452
rect	114	451	115	452
rect	115	451	116	452
rect	117	451	118	452
rect	118	451	119	452
rect	119	451	120	452
rect	120	451	121	452
rect	121	451	122	452
rect	122	451	123	452
rect	124	451	125	452
rect	125	451	126	452
rect	126	451	127	452
rect	127	451	128	452
rect	128	451	129	452
rect	129	451	130	452
rect	131	451	132	452
rect	132	451	133	452
rect	133	451	134	452
rect	134	451	135	452
rect	135	451	136	452
rect	136	451	137	452
rect	138	451	139	452
rect	139	451	140	452
rect	140	451	141	452
rect	141	451	142	452
rect	142	451	143	452
rect	143	451	144	452
rect	145	451	146	452
rect	146	451	147	452
rect	147	451	148	452
rect	148	451	149	452
rect	149	451	150	452
rect	150	451	151	452
rect	152	451	153	452
rect	153	451	154	452
rect	154	451	155	452
rect	155	451	156	452
rect	156	451	157	452
rect	157	451	158	452
rect	159	451	160	452
rect	160	451	161	452
rect	161	451	162	452
rect	162	451	163	452
rect	163	451	164	452
rect	164	451	165	452
rect	166	451	167	452
rect	167	451	168	452
rect	168	451	169	452
rect	169	451	170	452
rect	170	451	171	452
rect	171	451	172	452
<< metal1 >>
rect	70	0	71	1
rect	71	0	72	1
rect	57	2	58	3
rect	58	2	59	3
rect	59	2	60	3
rect	60	2	61	3
rect	61	2	62	3
rect	62	2	63	3
rect	63	2	64	3
rect	64	2	65	3
rect	65	2	66	3
rect	66	2	67	3
rect	67	2	68	3
rect	68	2	69	3
rect	70	2	71	3
rect	71	2	72	3
rect	73	2	74	3
rect	74	2	75	3
rect	75	2	76	3
rect	76	2	77	3
rect	77	2	78	3
rect	78	2	79	3
rect	79	2	80	3
rect	80	2	81	3
rect	81	2	82	3
rect	82	2	83	3
rect	83	2	84	3
rect	84	2	85	3
rect	85	2	86	3
rect	86	2	87	3
rect	87	2	88	3
rect	88	2	89	3
rect	89	2	90	3
rect	90	2	91	3
rect	91	2	92	3
rect	92	2	93	3
rect	93	2	94	3
rect	94	2	95	3
rect	95	2	96	3
rect	96	2	97	3
rect	97	2	98	3
rect	98	2	99	3
rect	99	2	100	3
rect	100	2	101	3
rect	101	2	102	3
rect	102	2	103	3
rect	103	2	104	3
rect	104	2	105	3
rect	105	2	106	3
rect	106	2	107	3
rect	107	2	108	3
rect	108	2	109	3
rect	109	2	110	3
rect	110	2	111	3
rect	111	2	112	3
rect	112	2	113	3
rect	113	2	114	3
rect	114	2	115	3
rect	115	2	116	3
rect	116	2	117	3
rect	117	2	118	3
rect	118	2	119	3
rect	119	2	120	3
rect	120	2	121	3
rect	121	2	122	3
rect	122	2	123	3
rect	123	2	124	3
rect	124	2	125	3
rect	125	2	126	3
rect	126	2	127	3
rect	127	2	128	3
rect	128	2	129	3
rect	129	2	130	3
rect	130	2	131	3
rect	191	2	192	3
rect	192	2	193	3
rect	44	4	45	5
rect	45	4	46	5
rect	46	4	47	5
rect	47	4	48	5
rect	48	4	49	5
rect	49	4	50	5
rect	50	4	51	5
rect	51	4	52	5
rect	52	4	53	5
rect	53	4	54	5
rect	54	4	55	5
rect	55	4	56	5
rect	57	4	58	5
rect	58	4	59	5
rect	59	4	60	5
rect	60	4	61	5
rect	61	4	62	5
rect	62	4	63	5
rect	63	4	64	5
rect	64	4	65	5
rect	65	4	66	5
rect	66	4	67	5
rect	67	4	68	5
rect	68	4	69	5
rect	70	4	71	5
rect	71	4	72	5
rect	73	4	74	5
rect	74	4	75	5
rect	75	4	76	5
rect	76	4	77	5
rect	77	4	78	5
rect	78	4	79	5
rect	79	4	80	5
rect	80	4	81	5
rect	81	4	82	5
rect	82	4	83	5
rect	83	4	84	5
rect	84	4	85	5
rect	85	4	86	5
rect	86	4	87	5
rect	87	4	88	5
rect	88	4	89	5
rect	89	4	90	5
rect	90	4	91	5
rect	91	4	92	5
rect	92	4	93	5
rect	93	4	94	5
rect	94	4	95	5
rect	95	4	96	5
rect	96	4	97	5
rect	97	4	98	5
rect	98	4	99	5
rect	99	4	100	5
rect	100	4	101	5
rect	101	4	102	5
rect	102	4	103	5
rect	103	4	104	5
rect	104	4	105	5
rect	105	4	106	5
rect	106	4	107	5
rect	107	4	108	5
rect	108	4	109	5
rect	119	4	120	5
rect	120	4	121	5
rect	121	4	122	5
rect	122	4	123	5
rect	123	4	124	5
rect	174	4	175	5
rect	175	4	176	5
rect	176	4	177	5
rect	177	4	178	5
rect	178	4	179	5
rect	179	4	180	5
rect	180	4	181	5
rect	181	4	182	5
rect	182	4	183	5
rect	183	4	184	5
rect	184	4	185	5
rect	185	4	186	5
rect	186	4	187	5
rect	187	4	188	5
rect	188	4	189	5
rect	189	4	190	5
rect	191	4	192	5
rect	192	4	193	5
rect	194	4	195	5
rect	195	4	196	5
rect	196	4	197	5
rect	197	4	198	5
rect	198	4	199	5
rect	199	4	200	5
rect	200	4	201	5
rect	201	4	202	5
rect	202	4	203	5
rect	203	4	204	5
rect	204	4	205	5
rect	205	4	206	5
rect	206	4	207	5
rect	207	4	208	5
rect	208	4	209	5
rect	209	4	210	5
rect	210	4	211	5
rect	211	4	212	5
rect	212	4	213	5
rect	213	4	214	5
rect	214	4	215	5
rect	215	4	216	5
rect	216	4	217	5
rect	217	4	218	5
rect	218	4	219	5
rect	219	4	220	5
rect	238	4	239	5
rect	239	4	240	5
rect	240	4	241	5
rect	241	4	242	5
rect	242	4	243	5
rect	247	4	248	5
rect	248	4	249	5
rect	249	4	250	5
rect	250	4	251	5
rect	251	4	252	5
rect	263	4	264	5
rect	264	4	265	5
rect	33	13	34	14
rect	34	13	35	14
rect	35	13	36	14
rect	36	13	37	14
rect	37	13	38	14
rect	38	13	39	14
rect	39	13	40	14
rect	40	13	41	14
rect	41	13	42	14
rect	42	13	43	14
rect	43	13	44	14
rect	44	13	45	14
rect	45	13	46	14
rect	46	13	47	14
rect	47	13	48	14
rect	48	13	49	14
rect	49	13	50	14
rect	50	13	51	14
rect	51	13	52	14
rect	52	13	53	14
rect	54	13	55	14
rect	55	13	56	14
rect	57	13	58	14
rect	58	13	59	14
rect	59	13	60	14
rect	60	13	61	14
rect	61	13	62	14
rect	62	13	63	14
rect	63	13	64	14
rect	64	13	65	14
rect	65	13	66	14
rect	66	13	67	14
rect	67	13	68	14
rect	68	13	69	14
rect	69	13	70	14
rect	70	13	71	14
rect	71	13	72	14
rect	73	13	74	14
rect	74	13	75	14
rect	75	13	76	14
rect	76	13	77	14
rect	77	13	78	14
rect	78	13	79	14
rect	79	13	80	14
rect	80	13	81	14
rect	81	13	82	14
rect	82	13	83	14
rect	83	13	84	14
rect	84	13	85	14
rect	86	13	87	14
rect	87	13	88	14
rect	88	13	89	14
rect	89	13	90	14
rect	90	13	91	14
rect	91	13	92	14
rect	92	13	93	14
rect	93	13	94	14
rect	94	13	95	14
rect	95	13	96	14
rect	96	13	97	14
rect	97	13	98	14
rect	98	13	99	14
rect	99	13	100	14
rect	100	13	101	14
rect	101	13	102	14
rect	102	13	103	14
rect	103	13	104	14
rect	104	13	105	14
rect	105	13	106	14
rect	106	13	107	14
rect	107	13	108	14
rect	108	13	109	14
rect	110	13	111	14
rect	111	13	112	14
rect	112	13	113	14
rect	113	13	114	14
rect	114	13	115	14
rect	115	13	116	14
rect	116	13	117	14
rect	117	13	118	14
rect	119	13	120	14
rect	120	13	121	14
rect	121	13	122	14
rect	122	13	123	14
rect	123	13	124	14
rect	124	13	125	14
rect	125	13	126	14
rect	126	13	127	14
rect	127	13	128	14
rect	128	13	129	14
rect	129	13	130	14
rect	130	13	131	14
rect	132	13	133	14
rect	133	13	134	14
rect	134	13	135	14
rect	135	13	136	14
rect	136	13	137	14
rect	137	13	138	14
rect	138	13	139	14
rect	139	13	140	14
rect	140	13	141	14
rect	141	13	142	14
rect	143	13	144	14
rect	144	13	145	14
rect	145	13	146	14
rect	146	13	147	14
rect	147	13	148	14
rect	148	13	149	14
rect	149	13	150	14
rect	150	13	151	14
rect	151	13	152	14
rect	152	13	153	14
rect	153	13	154	14
rect	154	13	155	14
rect	155	13	156	14
rect	156	13	157	14
rect	157	13	158	14
rect	158	13	159	14
rect	159	13	160	14
rect	160	13	161	14
rect	161	13	162	14
rect	162	13	163	14
rect	164	13	165	14
rect	165	13	166	14
rect	166	13	167	14
rect	167	13	168	14
rect	168	13	169	14
rect	169	13	170	14
rect	171	13	172	14
rect	172	13	173	14
rect	173	13	174	14
rect	174	13	175	14
rect	175	13	176	14
rect	176	13	177	14
rect	178	13	179	14
rect	179	13	180	14
rect	181	13	182	14
rect	182	13	183	14
rect	183	13	184	14
rect	184	13	185	14
rect	185	13	186	14
rect	186	13	187	14
rect	187	13	188	14
rect	188	13	189	14
rect	189	13	190	14
rect	191	13	192	14
rect	192	13	193	14
rect	193	13	194	14
rect	194	13	195	14
rect	195	13	196	14
rect	196	13	197	14
rect	197	13	198	14
rect	198	13	199	14
rect	199	13	200	14
rect	201	13	202	14
rect	202	13	203	14
rect	203	13	204	14
rect	204	13	205	14
rect	205	13	206	14
rect	206	13	207	14
rect	207	13	208	14
rect	208	13	209	14
rect	209	13	210	14
rect	210	13	211	14
rect	211	13	212	14
rect	212	13	213	14
rect	213	13	214	14
rect	215	13	216	14
rect	216	13	217	14
rect	217	13	218	14
rect	218	13	219	14
rect	219	13	220	14
rect	221	13	222	14
rect	222	13	223	14
rect	223	13	224	14
rect	224	13	225	14
rect	225	13	226	14
rect	226	13	227	14
rect	227	13	228	14
rect	228	13	229	14
rect	229	13	230	14
rect	230	13	231	14
rect	231	13	232	14
rect	232	13	233	14
rect	233	13	234	14
rect	234	13	235	14
rect	235	13	236	14
rect	236	13	237	14
rect	237	13	238	14
rect	238	13	239	14
rect	239	13	240	14
rect	240	13	241	14
rect	241	13	242	14
rect	242	13	243	14
rect	244	13	245	14
rect	245	13	246	14
rect	247	13	248	14
rect	248	13	249	14
rect	249	13	250	14
rect	250	13	251	14
rect	251	13	252	14
rect	181	15	182	16
rect	247	15	248	16
rect	248	15	249	16
rect	249	15	250	16
rect	250	15	251	16
rect	251	15	252	16
rect	252	15	253	16
rect	180	17	181	18
rect	181	17	182	18
rect	183	17	184	18
rect	184	17	185	18
rect	185	17	186	18
rect	186	17	187	18
rect	187	17	188	18
rect	188	17	189	18
rect	189	17	190	18
rect	190	17	191	18
rect	192	17	193	18
rect	193	17	194	18
rect	194	17	195	18
rect	195	17	196	18
rect	196	17	197	18
rect	197	17	198	18
rect	198	17	199	18
rect	199	17	200	18
rect	244	17	245	18
rect	245	17	246	18
rect	246	17	247	18
rect	247	17	248	18
rect	248	17	249	18
rect	249	17	250	18
rect	250	17	251	18
rect	251	17	252	18
rect	252	17	253	18
rect	254	17	255	18
rect	255	17	256	18
rect	256	17	257	18
rect	257	17	258	18
rect	258	17	259	18
rect	259	17	260	18
rect	260	17	261	18
rect	261	17	262	18
rect	263	17	264	18
rect	264	17	265	18
rect	96	19	97	20
rect	97	19	98	20
rect	98	19	99	20
rect	99	19	100	20
rect	100	19	101	20
rect	101	19	102	20
rect	102	19	103	20
rect	103	19	104	20
rect	104	19	105	20
rect	105	19	106	20
rect	106	19	107	20
rect	107	19	108	20
rect	109	19	110	20
rect	110	19	111	20
rect	111	19	112	20
rect	112	19	113	20
rect	113	19	114	20
rect	114	19	115	20
rect	115	19	116	20
rect	116	19	117	20
rect	117	19	118	20
rect	168	19	169	20
rect	169	19	170	20
rect	178	19	179	20
rect	180	19	181	20
rect	181	19	182	20
rect	183	19	184	20
rect	184	19	185	20
rect	185	19	186	20
rect	186	19	187	20
rect	187	19	188	20
rect	188	19	189	20
rect	189	19	190	20
rect	190	19	191	20
rect	192	19	193	20
rect	193	19	194	20
rect	194	19	195	20
rect	195	19	196	20
rect	196	19	197	20
rect	197	19	198	20
rect	198	19	199	20
rect	199	19	200	20
rect	210	19	211	20
rect	211	19	212	20
rect	212	19	213	20
rect	213	19	214	20
rect	215	19	216	20
rect	216	19	217	20
rect	217	19	218	20
rect	218	19	219	20
rect	219	19	220	20
rect	220	19	221	20
rect	222	19	223	20
rect	223	19	224	20
rect	224	19	225	20
rect	225	19	226	20
rect	226	19	227	20
rect	227	19	228	20
rect	228	19	229	20
rect	229	19	230	20
rect	230	19	231	20
rect	231	19	232	20
rect	232	19	233	20
rect	233	19	234	20
rect	234	19	235	20
rect	235	19	236	20
rect	236	19	237	20
rect	237	19	238	20
rect	238	19	239	20
rect	239	19	240	20
rect	240	19	241	20
rect	241	19	242	20
rect	242	19	243	20
rect	243	19	244	20
rect	244	19	245	20
rect	245	19	246	20
rect	246	19	247	20
rect	247	19	248	20
rect	248	19	249	20
rect	249	19	250	20
rect	250	19	251	20
rect	251	19	252	20
rect	252	19	253	20
rect	254	19	255	20
rect	255	19	256	20
rect	256	19	257	20
rect	257	19	258	20
rect	258	19	259	20
rect	259	19	260	20
rect	260	19	261	20
rect	261	19	262	20
rect	263	19	264	20
rect	264	19	265	20
rect	266	19	267	20
rect	267	19	268	20
rect	268	19	269	20
rect	269	19	270	20
rect	270	19	271	20
rect	271	19	272	20
rect	272	19	273	20
rect	273	19	274	20
rect	274	19	275	20
rect	275	19	276	20
rect	276	19	277	20
rect	277	19	278	20
rect	54	21	55	22
rect	55	21	56	22
rect	86	21	87	22
rect	87	21	88	22
rect	88	21	89	22
rect	89	21	90	22
rect	90	21	91	22
rect	91	21	92	22
rect	92	21	93	22
rect	93	21	94	22
rect	94	21	95	22
rect	96	21	97	22
rect	97	21	98	22
rect	98	21	99	22
rect	99	21	100	22
rect	100	21	101	22
rect	101	21	102	22
rect	102	21	103	22
rect	103	21	104	22
rect	104	21	105	22
rect	105	21	106	22
rect	106	21	107	22
rect	107	21	108	22
rect	109	21	110	22
rect	110	21	111	22
rect	111	21	112	22
rect	112	21	113	22
rect	113	21	114	22
rect	114	21	115	22
rect	115	21	116	22
rect	116	21	117	22
rect	117	21	118	22
rect	118	21	119	22
rect	119	21	120	22
rect	120	21	121	22
rect	121	21	122	22
rect	122	21	123	22
rect	123	21	124	22
rect	124	21	125	22
rect	125	21	126	22
rect	126	21	127	22
rect	127	21	128	22
rect	128	21	129	22
rect	129	21	130	22
rect	130	21	131	22
rect	164	21	165	22
rect	165	21	166	22
rect	166	21	167	22
rect	168	21	169	22
rect	169	21	170	22
rect	170	21	171	22
rect	171	21	172	22
rect	172	21	173	22
rect	173	21	174	22
rect	174	21	175	22
rect	175	21	176	22
rect	176	21	177	22
rect	177	21	178	22
rect	178	21	179	22
rect	180	21	181	22
rect	181	21	182	22
rect	183	21	184	22
rect	184	21	185	22
rect	185	21	186	22
rect	186	21	187	22
rect	187	21	188	22
rect	188	21	189	22
rect	189	21	190	22
rect	190	21	191	22
rect	192	21	193	22
rect	193	21	194	22
rect	194	21	195	22
rect	195	21	196	22
rect	196	21	197	22
rect	197	21	198	22
rect	198	21	199	22
rect	199	21	200	22
rect	201	21	202	22
rect	202	21	203	22
rect	203	21	204	22
rect	204	21	205	22
rect	205	21	206	22
rect	206	21	207	22
rect	207	21	208	22
rect	208	21	209	22
rect	210	21	211	22
rect	211	21	212	22
rect	212	21	213	22
rect	213	21	214	22
rect	215	21	216	22
rect	216	21	217	22
rect	217	21	218	22
rect	218	21	219	22
rect	219	21	220	22
rect	220	21	221	22
rect	222	21	223	22
rect	223	21	224	22
rect	224	21	225	22
rect	225	21	226	22
rect	226	21	227	22
rect	227	21	228	22
rect	228	21	229	22
rect	229	21	230	22
rect	230	21	231	22
rect	231	21	232	22
rect	232	21	233	22
rect	233	21	234	22
rect	234	21	235	22
rect	235	21	236	22
rect	236	21	237	22
rect	237	21	238	22
rect	238	21	239	22
rect	239	21	240	22
rect	240	21	241	22
rect	241	21	242	22
rect	242	21	243	22
rect	243	21	244	22
rect	244	21	245	22
rect	245	21	246	22
rect	246	21	247	22
rect	247	21	248	22
rect	248	21	249	22
rect	249	21	250	22
rect	250	21	251	22
rect	251	21	252	22
rect	252	21	253	22
rect	254	21	255	22
rect	255	21	256	22
rect	286	21	287	22
rect	287	21	288	22
rect	288	21	289	22
rect	289	21	290	22
rect	290	21	291	22
rect	291	21	292	22
rect	292	21	293	22
rect	293	21	294	22
rect	294	21	295	22
rect	295	21	296	22
rect	296	21	297	22
rect	297	21	298	22
rect	298	21	299	22
rect	299	21	300	22
rect	300	21	301	22
rect	301	21	302	22
rect	12	23	13	24
rect	13	23	14	24
rect	51	23	52	24
rect	52	23	53	24
rect	63	23	64	24
rect	64	23	65	24
rect	65	23	66	24
rect	66	23	67	24
rect	67	23	68	24
rect	68	23	69	24
rect	69	23	70	24
rect	70	23	71	24
rect	72	23	73	24
rect	73	23	74	24
rect	74	23	75	24
rect	75	23	76	24
rect	76	23	77	24
rect	77	23	78	24
rect	78	23	79	24
rect	79	23	80	24
rect	80	23	81	24
rect	81	23	82	24
rect	82	23	83	24
rect	83	23	84	24
rect	84	23	85	24
rect	85	23	86	24
rect	86	23	87	24
rect	87	23	88	24
rect	88	23	89	24
rect	89	23	90	24
rect	90	23	91	24
rect	91	23	92	24
rect	92	23	93	24
rect	93	23	94	24
rect	94	23	95	24
rect	96	23	97	24
rect	97	23	98	24
rect	98	23	99	24
rect	99	23	100	24
rect	100	23	101	24
rect	101	23	102	24
rect	102	23	103	24
rect	103	23	104	24
rect	104	23	105	24
rect	105	23	106	24
rect	106	23	107	24
rect	107	23	108	24
rect	109	23	110	24
rect	110	23	111	24
rect	111	23	112	24
rect	112	23	113	24
rect	113	23	114	24
rect	114	23	115	24
rect	115	23	116	24
rect	116	23	117	24
rect	117	23	118	24
rect	118	23	119	24
rect	119	23	120	24
rect	120	23	121	24
rect	121	23	122	24
rect	122	23	123	24
rect	123	23	124	24
rect	124	23	125	24
rect	143	23	144	24
rect	144	23	145	24
rect	145	23	146	24
rect	146	23	147	24
rect	147	23	148	24
rect	148	23	149	24
rect	149	23	150	24
rect	150	23	151	24
rect	151	23	152	24
rect	162	23	163	24
rect	163	23	164	24
rect	164	23	165	24
rect	165	23	166	24
rect	166	23	167	24
rect	168	23	169	24
rect	169	23	170	24
rect	170	23	171	24
rect	171	23	172	24
rect	172	23	173	24
rect	173	23	174	24
rect	174	23	175	24
rect	175	23	176	24
rect	176	23	177	24
rect	177	23	178	24
rect	178	23	179	24
rect	180	23	181	24
rect	181	23	182	24
rect	183	23	184	24
rect	184	23	185	24
rect	185	23	186	24
rect	186	23	187	24
rect	187	23	188	24
rect	188	23	189	24
rect	189	23	190	24
rect	190	23	191	24
rect	192	23	193	24
rect	193	23	194	24
rect	194	23	195	24
rect	195	23	196	24
rect	196	23	197	24
rect	197	23	198	24
rect	198	23	199	24
rect	199	23	200	24
rect	201	23	202	24
rect	202	23	203	24
rect	203	23	204	24
rect	204	23	205	24
rect	205	23	206	24
rect	206	23	207	24
rect	207	23	208	24
rect	208	23	209	24
rect	210	23	211	24
rect	211	23	212	24
rect	212	23	213	24
rect	213	23	214	24
rect	219	23	220	24
rect	220	23	221	24
rect	222	23	223	24
rect	223	23	224	24
rect	224	23	225	24
rect	225	23	226	24
rect	226	23	227	24
rect	245	23	246	24
rect	246	23	247	24
rect	263	23	264	24
rect	264	23	265	24
rect	266	23	267	24
rect	267	23	268	24
rect	268	23	269	24
rect	269	23	270	24
rect	270	23	271	24
rect	271	23	272	24
rect	272	23	273	24
rect	273	23	274	24
rect	274	23	275	24
rect	275	23	276	24
rect	276	23	277	24
rect	277	23	278	24
rect	279	23	280	24
rect	280	23	281	24
rect	281	23	282	24
rect	282	23	283	24
rect	283	23	284	24
rect	284	23	285	24
rect	286	23	287	24
rect	287	23	288	24
rect	288	23	289	24
rect	289	23	290	24
rect	290	23	291	24
rect	291	23	292	24
rect	292	23	293	24
rect	293	23	294	24
rect	294	23	295	24
rect	295	23	296	24
rect	12	25	13	26
rect	13	25	14	26
rect	15	25	16	26
rect	16	25	17	26
rect	17	25	18	26
rect	18	25	19	26
rect	19	25	20	26
rect	20	25	21	26
rect	21	25	22	26
rect	22	25	23	26
rect	23	25	24	26
rect	24	25	25	26
rect	25	25	26	26
rect	26	25	27	26
rect	27	25	28	26
rect	28	25	29	26
rect	29	25	30	26
rect	31	25	32	26
rect	32	25	33	26
rect	33	25	34	26
rect	34	25	35	26
rect	35	25	36	26
rect	36	25	37	26
rect	37	25	38	26
rect	38	25	39	26
rect	39	25	40	26
rect	40	25	41	26
rect	41	25	42	26
rect	42	25	43	26
rect	43	25	44	26
rect	44	25	45	26
rect	45	25	46	26
rect	46	25	47	26
rect	47	25	48	26
rect	48	25	49	26
rect	49	25	50	26
rect	51	25	52	26
rect	52	25	53	26
rect	54	25	55	26
rect	55	25	56	26
rect	56	25	57	26
rect	57	25	58	26
rect	58	25	59	26
rect	59	25	60	26
rect	60	25	61	26
rect	61	25	62	26
rect	63	25	64	26
rect	64	25	65	26
rect	65	25	66	26
rect	66	25	67	26
rect	67	25	68	26
rect	68	25	69	26
rect	69	25	70	26
rect	70	25	71	26
rect	72	25	73	26
rect	73	25	74	26
rect	74	25	75	26
rect	75	25	76	26
rect	76	25	77	26
rect	77	25	78	26
rect	78	25	79	26
rect	79	25	80	26
rect	80	25	81	26
rect	81	25	82	26
rect	82	25	83	26
rect	83	25	84	26
rect	84	25	85	26
rect	85	25	86	26
rect	86	25	87	26
rect	87	25	88	26
rect	88	25	89	26
rect	89	25	90	26
rect	90	25	91	26
rect	91	25	92	26
rect	92	25	93	26
rect	93	25	94	26
rect	94	25	95	26
rect	96	25	97	26
rect	97	25	98	26
rect	98	25	99	26
rect	99	25	100	26
rect	100	25	101	26
rect	101	25	102	26
rect	102	25	103	26
rect	103	25	104	26
rect	104	25	105	26
rect	105	25	106	26
rect	106	25	107	26
rect	107	25	108	26
rect	109	25	110	26
rect	110	25	111	26
rect	111	25	112	26
rect	112	25	113	26
rect	113	25	114	26
rect	114	25	115	26
rect	115	25	116	26
rect	116	25	117	26
rect	117	25	118	26
rect	118	25	119	26
rect	119	25	120	26
rect	120	25	121	26
rect	121	25	122	26
rect	122	25	123	26
rect	123	25	124	26
rect	124	25	125	26
rect	126	25	127	26
rect	127	25	128	26
rect	128	25	129	26
rect	129	25	130	26
rect	130	25	131	26
rect	131	25	132	26
rect	132	25	133	26
rect	133	25	134	26
rect	134	25	135	26
rect	135	25	136	26
rect	136	25	137	26
rect	137	25	138	26
rect	138	25	139	26
rect	139	25	140	26
rect	140	25	141	26
rect	141	25	142	26
rect	142	25	143	26
rect	143	25	144	26
rect	144	25	145	26
rect	145	25	146	26
rect	146	25	147	26
rect	147	25	148	26
rect	148	25	149	26
rect	149	25	150	26
rect	150	25	151	26
rect	151	25	152	26
rect	153	25	154	26
rect	154	25	155	26
rect	155	25	156	26
rect	156	25	157	26
rect	157	25	158	26
rect	158	25	159	26
rect	159	25	160	26
rect	160	25	161	26
rect	162	25	163	26
rect	163	25	164	26
rect	171	25	172	26
rect	172	25	173	26
rect	173	25	174	26
rect	174	25	175	26
rect	175	25	176	26
rect	189	25	190	26
rect	190	25	191	26
rect	192	25	193	26
rect	193	25	194	26
rect	194	25	195	26
rect	195	25	196	26
rect	196	25	197	26
rect	197	25	198	26
rect	198	25	199	26
rect	199	25	200	26
rect	201	25	202	26
rect	202	25	203	26
rect	203	25	204	26
rect	204	25	205	26
rect	205	25	206	26
rect	206	25	207	26
rect	207	25	208	26
rect	208	25	209	26
rect	210	25	211	26
rect	211	25	212	26
rect	212	25	213	26
rect	213	25	214	26
rect	214	25	215	26
rect	215	25	216	26
rect	216	25	217	26
rect	217	25	218	26
rect	219	25	220	26
rect	220	25	221	26
rect	222	25	223	26
rect	223	25	224	26
rect	224	25	225	26
rect	225	25	226	26
rect	226	25	227	26
rect	228	25	229	26
rect	229	25	230	26
rect	230	25	231	26
rect	231	25	232	26
rect	232	25	233	26
rect	233	25	234	26
rect	234	25	235	26
rect	235	25	236	26
rect	236	25	237	26
rect	237	25	238	26
rect	238	25	239	26
rect	239	25	240	26
rect	240	25	241	26
rect	241	25	242	26
rect	242	25	243	26
rect	243	25	244	26
rect	245	25	246	26
rect	246	25	247	26
rect	248	25	249	26
rect	249	25	250	26
rect	250	25	251	26
rect	251	25	252	26
rect	252	25	253	26
rect	254	25	255	26
rect	255	25	256	26
rect	257	25	258	26
rect	258	25	259	26
rect	259	25	260	26
rect	260	25	261	26
rect	261	25	262	26
rect	262	25	263	26
rect	263	25	264	26
rect	264	25	265	26
rect	266	25	267	26
rect	267	25	268	26
rect	268	25	269	26
rect	269	25	270	26
rect	270	25	271	26
rect	271	25	272	26
rect	272	25	273	26
rect	273	25	274	26
rect	274	25	275	26
rect	275	25	276	26
rect	276	25	277	26
rect	277	25	278	26
rect	279	25	280	26
rect	280	25	281	26
rect	281	25	282	26
rect	282	25	283	26
rect	283	25	284	26
rect	284	25	285	26
rect	286	25	287	26
rect	287	25	288	26
rect	288	25	289	26
rect	289	25	290	26
rect	290	25	291	26
rect	291	25	292	26
rect	292	25	293	26
rect	293	25	294	26
rect	294	25	295	26
rect	295	25	296	26
rect	297	25	298	26
rect	298	25	299	26
rect	299	25	300	26
rect	300	25	301	26
rect	301	25	302	26
rect	303	25	304	26
rect	304	25	305	26
rect	216	34	217	35
rect	217	34	218	35
rect	204	36	205	37
rect	205	36	206	37
rect	206	36	207	37
rect	207	36	208	37
rect	208	36	209	37
rect	210	36	211	37
rect	211	36	212	37
rect	212	36	213	37
rect	213	36	214	37
rect	214	36	215	37
rect	216	36	217	37
rect	217	36	218	37
rect	201	38	202	39
rect	202	38	203	39
rect	198	40	199	41
rect	199	40	200	41
rect	200	40	201	41
rect	201	40	202	41
rect	202	40	203	41
rect	204	40	205	41
rect	205	40	206	41
rect	206	40	207	41
rect	207	40	208	41
rect	208	40	209	41
rect	210	40	211	41
rect	211	40	212	41
rect	212	40	213	41
rect	213	40	214	41
rect	214	40	215	41
rect	216	40	217	41
rect	217	40	218	41
rect	219	40	220	41
rect	220	40	221	41
rect	222	40	223	41
rect	223	40	224	41
rect	224	40	225	41
rect	225	40	226	41
rect	226	40	227	41
rect	227	40	228	41
rect	228	40	229	41
rect	229	40	230	41
rect	230	40	231	41
rect	232	40	233	41
rect	233	40	234	41
rect	234	40	235	41
rect	235	40	236	41
rect	236	40	237	41
rect	237	40	238	41
rect	238	40	239	41
rect	239	40	240	41
rect	240	40	241	41
rect	241	40	242	41
rect	242	40	243	41
rect	243	40	244	41
rect	245	40	246	41
rect	246	40	247	41
rect	247	40	248	41
rect	248	40	249	41
rect	249	40	250	41
rect	251	40	252	41
rect	252	40	253	41
rect	254	40	255	41
rect	255	40	256	41
rect	257	40	258	41
rect	258	40	259	41
rect	259	40	260	41
rect	260	40	261	41
rect	261	40	262	41
rect	262	40	263	41
rect	263	40	264	41
rect	264	40	265	41
rect	266	40	267	41
rect	267	40	268	41
rect	268	40	269	41
rect	269	40	270	41
rect	270	40	271	41
rect	271	40	272	41
rect	272	40	273	41
rect	273	40	274	41
rect	274	40	275	41
rect	275	40	276	41
rect	276	40	277	41
rect	277	40	278	41
rect	279	40	280	41
rect	280	40	281	41
rect	281	40	282	41
rect	282	40	283	41
rect	283	40	284	41
rect	284	40	285	41
rect	285	40	286	41
rect	286	40	287	41
rect	287	40	288	41
rect	288	40	289	41
rect	289	40	290	41
rect	290	40	291	41
rect	291	40	292	41
rect	292	40	293	41
rect	293	40	294	41
rect	294	40	295	41
rect	295	40	296	41
rect	296	40	297	41
rect	297	40	298	41
rect	298	40	299	41
rect	299	40	300	41
rect	300	40	301	41
rect	301	40	302	41
rect	303	40	304	41
rect	304	40	305	41
rect	306	40	307	41
rect	307	40	308	41
rect	308	40	309	41
rect	177	42	178	43
rect	178	42	179	43
rect	180	42	181	43
rect	181	42	182	43
rect	183	42	184	43
rect	184	42	185	43
rect	185	42	186	43
rect	186	42	187	43
rect	187	42	188	43
rect	188	42	189	43
rect	189	42	190	43
rect	190	42	191	43
rect	192	42	193	43
rect	193	42	194	43
rect	195	42	196	43
rect	196	42	197	43
rect	197	42	198	43
rect	198	42	199	43
rect	199	42	200	43
rect	266	42	267	43
rect	267	42	268	43
rect	268	42	269	43
rect	269	42	270	43
rect	270	42	271	43
rect	271	42	272	43
rect	272	42	273	43
rect	273	42	274	43
rect	274	42	275	43
rect	275	42	276	43
rect	174	44	175	45
rect	175	44	176	45
rect	176	44	177	45
rect	177	44	178	45
rect	178	44	179	45
rect	180	44	181	45
rect	181	44	182	45
rect	183	44	184	45
rect	184	44	185	45
rect	185	44	186	45
rect	186	44	187	45
rect	187	44	188	45
rect	188	44	189	45
rect	189	44	190	45
rect	190	44	191	45
rect	192	44	193	45
rect	193	44	194	45
rect	195	44	196	45
rect	196	44	197	45
rect	262	44	263	45
rect	263	44	264	45
rect	264	44	265	45
rect	265	44	266	45
rect	266	44	267	45
rect	267	44	268	45
rect	268	44	269	45
rect	269	44	270	45
rect	270	44	271	45
rect	271	44	272	45
rect	272	44	273	45
rect	168	46	169	47
rect	169	46	170	47
rect	170	46	171	47
rect	171	46	172	47
rect	172	46	173	47
rect	173	46	174	47
rect	174	46	175	47
rect	175	46	176	47
rect	232	46	233	47
rect	233	46	234	47
rect	234	46	235	47
rect	235	46	236	47
rect	236	46	237	47
rect	237	46	238	47
rect	238	46	239	47
rect	239	46	240	47
rect	240	46	241	47
rect	241	46	242	47
rect	242	46	243	47
rect	243	46	244	47
rect	245	46	246	47
rect	259	46	260	47
rect	260	46	261	47
rect	262	46	263	47
rect	263	46	264	47
rect	264	46	265	47
rect	265	46	266	47
rect	266	46	267	47
rect	267	46	268	47
rect	268	46	269	47
rect	269	46	270	47
rect	165	48	166	49
rect	166	48	167	49
rect	167	48	168	49
rect	168	48	169	49
rect	169	48	170	49
rect	170	48	171	49
rect	171	48	172	49
rect	172	48	173	49
rect	228	48	229	49
rect	229	48	230	49
rect	230	48	231	49
rect	231	48	232	49
rect	232	48	233	49
rect	251	48	252	49
rect	252	48	253	49
rect	254	48	255	49
rect	255	48	256	49
rect	257	48	258	49
rect	259	48	260	49
rect	260	48	261	49
rect	262	48	263	49
rect	263	48	264	49
rect	264	48	265	49
rect	265	48	266	49
rect	266	48	267	49
rect	267	48	268	49
rect	268	48	269	49
rect	269	48	270	49
rect	271	48	272	49
rect	272	48	273	49
rect	274	48	275	49
rect	275	48	276	49
rect	277	48	278	49
rect	279	48	280	49
rect	280	48	281	49
rect	281	48	282	49
rect	282	48	283	49
rect	283	48	284	49
rect	284	48	285	49
rect	285	48	286	49
rect	286	48	287	49
rect	287	48	288	49
rect	288	48	289	49
rect	289	48	290	49
rect	290	48	291	49
rect	291	48	292	49
rect	292	48	293	49
rect	293	48	294	49
rect	294	48	295	49
rect	295	48	296	49
rect	296	48	297	49
rect	297	48	298	49
rect	298	48	299	49
rect	299	48	300	49
rect	120	50	121	51
rect	121	50	122	51
rect	153	50	154	51
rect	154	50	155	51
rect	155	50	156	51
rect	156	50	157	51
rect	157	50	158	51
rect	158	50	159	51
rect	159	50	160	51
rect	160	50	161	51
rect	162	50	163	51
rect	163	50	164	51
rect	164	50	165	51
rect	165	50	166	51
rect	166	50	167	51
rect	171	50	172	51
rect	172	50	173	51
rect	174	50	175	51
rect	175	50	176	51
rect	177	50	178	51
rect	178	50	179	51
rect	180	50	181	51
rect	181	50	182	51
rect	207	50	208	51
rect	208	50	209	51
rect	222	50	223	51
rect	223	50	224	51
rect	224	50	225	51
rect	225	50	226	51
rect	226	50	227	51
rect	228	50	229	51
rect	229	50	230	51
rect	241	50	242	51
rect	242	50	243	51
rect	243	50	244	51
rect	245	50	246	51
rect	247	50	248	51
rect	248	50	249	51
rect	249	50	250	51
rect	250	50	251	51
rect	251	50	252	51
rect	252	50	253	51
rect	254	50	255	51
rect	255	50	256	51
rect	257	50	258	51
rect	259	50	260	51
rect	260	50	261	51
rect	262	50	263	51
rect	263	50	264	51
rect	264	50	265	51
rect	265	50	266	51
rect	266	50	267	51
rect	267	50	268	51
rect	268	50	269	51
rect	269	50	270	51
rect	271	50	272	51
rect	272	50	273	51
rect	274	50	275	51
rect	275	50	276	51
rect	277	50	278	51
rect	279	50	280	51
rect	280	50	281	51
rect	281	50	282	51
rect	282	50	283	51
rect	283	50	284	51
rect	284	50	285	51
rect	285	50	286	51
rect	286	50	287	51
rect	287	50	288	51
rect	306	50	307	51
rect	307	50	308	51
rect	308	50	309	51
rect	310	50	311	51
rect	311	50	312	51
rect	312	50	313	51
rect	313	50	314	51
rect	314	50	315	51
rect	315	50	316	51
rect	316	50	317	51
rect	317	50	318	51
rect	318	50	319	51
rect	319	50	320	51
rect	320	50	321	51
rect	321	50	322	51
rect	322	50	323	51
rect	323	50	324	51
rect	324	50	325	51
rect	325	50	326	51
rect	326	50	327	51
rect	327	50	328	51
rect	328	50	329	51
rect	329	50	330	51
rect	57	52	58	53
rect	58	52	59	53
rect	59	52	60	53
rect	60	52	61	53
rect	61	52	62	53
rect	78	52	79	53
rect	79	52	80	53
rect	80	52	81	53
rect	81	52	82	53
rect	82	52	83	53
rect	83	52	84	53
rect	84	52	85	53
rect	85	52	86	53
rect	86	52	87	53
rect	87	52	88	53
rect	88	52	89	53
rect	89	52	90	53
rect	90	52	91	53
rect	91	52	92	53
rect	92	52	93	53
rect	93	52	94	53
rect	94	52	95	53
rect	95	52	96	53
rect	96	52	97	53
rect	97	52	98	53
rect	98	52	99	53
rect	99	52	100	53
rect	100	52	101	53
rect	101	52	102	53
rect	102	52	103	53
rect	103	52	104	53
rect	104	52	105	53
rect	105	52	106	53
rect	106	52	107	53
rect	107	52	108	53
rect	109	52	110	53
rect	110	52	111	53
rect	111	52	112	53
rect	112	52	113	53
rect	113	52	114	53
rect	115	52	116	53
rect	116	52	117	53
rect	117	52	118	53
rect	118	52	119	53
rect	120	52	121	53
rect	121	52	122	53
rect	123	52	124	53
rect	124	52	125	53
rect	125	52	126	53
rect	126	52	127	53
rect	127	52	128	53
rect	128	52	129	53
rect	129	52	130	53
rect	130	52	131	53
rect	131	52	132	53
rect	132	52	133	53
rect	133	52	134	53
rect	134	52	135	53
rect	135	52	136	53
rect	136	52	137	53
rect	137	52	138	53
rect	138	52	139	53
rect	139	52	140	53
rect	140	52	141	53
rect	141	52	142	53
rect	142	52	143	53
rect	143	52	144	53
rect	144	52	145	53
rect	145	52	146	53
rect	147	52	148	53
rect	148	52	149	53
rect	150	52	151	53
rect	151	52	152	53
rect	152	52	153	53
rect	153	52	154	53
rect	154	52	155	53
rect	155	52	156	53
rect	156	52	157	53
rect	157	52	158	53
rect	158	52	159	53
rect	159	52	160	53
rect	160	52	161	53
rect	162	52	163	53
rect	163	52	164	53
rect	164	52	165	53
rect	165	52	166	53
rect	166	52	167	53
rect	168	52	169	53
rect	169	52	170	53
rect	171	52	172	53
rect	172	52	173	53
rect	174	52	175	53
rect	175	52	176	53
rect	177	52	178	53
rect	178	52	179	53
rect	180	52	181	53
rect	181	52	182	53
rect	182	52	183	53
rect	183	52	184	53
rect	184	52	185	53
rect	185	52	186	53
rect	186	52	187	53
rect	187	52	188	53
rect	188	52	189	53
rect	189	52	190	53
rect	190	52	191	53
rect	192	52	193	53
rect	193	52	194	53
rect	195	52	196	53
rect	196	52	197	53
rect	198	52	199	53
rect	199	52	200	53
rect	201	52	202	53
rect	202	52	203	53
rect	204	52	205	53
rect	205	52	206	53
rect	207	52	208	53
rect	208	52	209	53
rect	209	52	210	53
rect	210	52	211	53
rect	211	52	212	53
rect	212	52	213	53
rect	213	52	214	53
rect	214	52	215	53
rect	216	52	217	53
rect	217	52	218	53
rect	219	52	220	53
rect	220	52	221	53
rect	221	52	222	53
rect	222	52	223	53
rect	223	52	224	53
rect	224	52	225	53
rect	225	52	226	53
rect	226	52	227	53
rect	228	52	229	53
rect	229	52	230	53
rect	231	52	232	53
rect	232	52	233	53
rect	234	52	235	53
rect	235	52	236	53
rect	236	52	237	53
rect	237	52	238	53
rect	238	52	239	53
rect	239	52	240	53
rect	241	52	242	53
rect	242	52	243	53
rect	243	52	244	53
rect	245	52	246	53
rect	247	52	248	53
rect	248	52	249	53
rect	249	52	250	53
rect	250	52	251	53
rect	251	52	252	53
rect	252	52	253	53
rect	254	52	255	53
rect	255	52	256	53
rect	257	52	258	53
rect	259	52	260	53
rect	260	52	261	53
rect	262	52	263	53
rect	263	52	264	53
rect	264	52	265	53
rect	265	52	266	53
rect	266	52	267	53
rect	303	52	304	53
rect	304	52	305	53
rect	305	52	306	53
rect	306	52	307	53
rect	307	52	308	53
rect	308	52	309	53
rect	310	52	311	53
rect	311	52	312	53
rect	312	52	313	53
rect	313	52	314	53
rect	314	52	315	53
rect	315	52	316	53
rect	316	52	317	53
rect	317	52	318	53
rect	318	52	319	53
rect	319	52	320	53
rect	320	52	321	53
rect	321	52	322	53
rect	322	52	323	53
rect	323	52	324	53
rect	324	52	325	53
rect	325	52	326	53
rect	326	52	327	53
rect	327	52	328	53
rect	328	52	329	53
rect	329	52	330	53
rect	331	52	332	53
rect	332	52	333	53
rect	333	52	334	53
rect	334	52	335	53
rect	335	52	336	53
rect	336	52	337	53
rect	337	52	338	53
rect	338	52	339	53
rect	54	54	55	55
rect	55	54	56	55
rect	56	54	57	55
rect	57	54	58	55
rect	58	54	59	55
rect	59	54	60	55
rect	60	54	61	55
rect	61	54	62	55
rect	72	54	73	55
rect	73	54	74	55
rect	74	54	75	55
rect	75	54	76	55
rect	76	54	77	55
rect	77	54	78	55
rect	78	54	79	55
rect	79	54	80	55
rect	109	54	110	55
rect	115	54	116	55
rect	116	54	117	55
rect	117	54	118	55
rect	118	54	119	55
rect	120	54	121	55
rect	121	54	122	55
rect	123	54	124	55
rect	124	54	125	55
rect	125	54	126	55
rect	126	54	127	55
rect	127	54	128	55
rect	150	54	151	55
rect	151	54	152	55
rect	152	54	153	55
rect	153	54	154	55
rect	154	54	155	55
rect	155	54	156	55
rect	156	54	157	55
rect	157	54	158	55
rect	165	54	166	55
rect	166	54	167	55
rect	168	54	169	55
rect	169	54	170	55
rect	171	54	172	55
rect	172	54	173	55
rect	174	54	175	55
rect	175	54	176	55
rect	177	54	178	55
rect	178	54	179	55
rect	189	54	190	55
rect	190	54	191	55
rect	195	54	196	55
rect	196	54	197	55
rect	198	54	199	55
rect	199	54	200	55
rect	201	54	202	55
rect	202	54	203	55
rect	204	54	205	55
rect	205	54	206	55
rect	207	54	208	55
rect	208	54	209	55
rect	209	54	210	55
rect	210	54	211	55
rect	211	54	212	55
rect	212	54	213	55
rect	213	54	214	55
rect	214	54	215	55
rect	216	54	217	55
rect	217	54	218	55
rect	219	54	220	55
rect	220	54	221	55
rect	221	54	222	55
rect	222	54	223	55
rect	223	54	224	55
rect	224	54	225	55
rect	225	54	226	55
rect	226	54	227	55
rect	228	54	229	55
rect	229	54	230	55
rect	231	54	232	55
rect	232	54	233	55
rect	234	54	235	55
rect	235	54	236	55
rect	236	54	237	55
rect	237	54	238	55
rect	238	54	239	55
rect	239	54	240	55
rect	241	54	242	55
rect	242	54	243	55
rect	243	54	244	55
rect	245	54	246	55
rect	247	54	248	55
rect	248	54	249	55
rect	249	54	250	55
rect	250	54	251	55
rect	251	54	252	55
rect	252	54	253	55
rect	254	54	255	55
rect	255	54	256	55
rect	257	54	258	55
rect	259	54	260	55
rect	260	54	261	55
rect	262	54	263	55
rect	263	54	264	55
rect	264	54	265	55
rect	265	54	266	55
rect	266	54	267	55
rect	268	54	269	55
rect	269	54	270	55
rect	271	54	272	55
rect	272	54	273	55
rect	274	54	275	55
rect	275	54	276	55
rect	277	54	278	55
rect	279	54	280	55
rect	280	54	281	55
rect	281	54	282	55
rect	282	54	283	55
rect	283	54	284	55
rect	284	54	285	55
rect	285	54	286	55
rect	286	54	287	55
rect	287	54	288	55
rect	289	54	290	55
rect	290	54	291	55
rect	291	54	292	55
rect	292	54	293	55
rect	293	54	294	55
rect	294	54	295	55
rect	295	54	296	55
rect	296	54	297	55
rect	297	54	298	55
rect	298	54	299	55
rect	299	54	300	55
rect	301	54	302	55
rect	302	54	303	55
rect	303	54	304	55
rect	304	54	305	55
rect	305	54	306	55
rect	306	54	307	55
rect	307	54	308	55
rect	308	54	309	55
rect	310	54	311	55
rect	311	54	312	55
rect	312	54	313	55
rect	313	54	314	55
rect	314	54	315	55
rect	315	54	316	55
rect	316	54	317	55
rect	317	54	318	55
rect	318	54	319	55
rect	319	54	320	55
rect	320	54	321	55
rect	321	54	322	55
rect	322	54	323	55
rect	323	54	324	55
rect	324	54	325	55
rect	325	54	326	55
rect	326	54	327	55
rect	327	54	328	55
rect	328	54	329	55
rect	329	54	330	55
rect	331	54	332	55
rect	332	54	333	55
rect	333	54	334	55
rect	334	54	335	55
rect	335	54	336	55
rect	336	54	337	55
rect	337	54	338	55
rect	338	54	339	55
rect	340	54	341	55
rect	341	54	342	55
rect	342	54	343	55
rect	343	54	344	55
rect	344	54	345	55
rect	345	54	346	55
rect	346	54	347	55
rect	347	54	348	55
rect	348	54	349	55
rect	349	54	350	55
rect	350	54	351	55
rect	351	54	352	55
rect	352	54	353	55
rect	353	54	354	55
rect	354	54	355	55
rect	355	54	356	55
rect	356	54	357	55
rect	35	56	36	57
rect	36	56	37	57
rect	37	56	38	57
rect	38	56	39	57
rect	39	56	40	57
rect	40	56	41	57
rect	41	56	42	57
rect	42	56	43	57
rect	43	56	44	57
rect	44	56	45	57
rect	45	56	46	57
rect	46	56	47	57
rect	48	56	49	57
rect	49	56	50	57
rect	50	56	51	57
rect	51	56	52	57
rect	52	56	53	57
rect	53	56	54	57
rect	54	56	55	57
rect	55	56	56	57
rect	56	56	57	57
rect	57	56	58	57
rect	58	56	59	57
rect	59	56	60	57
rect	60	56	61	57
rect	61	56	62	57
rect	63	56	64	57
rect	64	56	65	57
rect	65	56	66	57
rect	66	56	67	57
rect	67	56	68	57
rect	68	56	69	57
rect	69	56	70	57
rect	70	56	71	57
rect	71	56	72	57
rect	72	56	73	57
rect	73	56	74	57
rect	74	56	75	57
rect	75	56	76	57
rect	76	56	77	57
rect	77	56	78	57
rect	78	56	79	57
rect	79	56	80	57
rect	81	56	82	57
rect	82	56	83	57
rect	83	56	84	57
rect	84	56	85	57
rect	85	56	86	57
rect	86	56	87	57
rect	87	56	88	57
rect	88	56	89	57
rect	89	56	90	57
rect	90	56	91	57
rect	91	56	92	57
rect	92	56	93	57
rect	93	56	94	57
rect	94	56	95	57
rect	95	56	96	57
rect	96	56	97	57
rect	97	56	98	57
rect	98	56	99	57
rect	99	56	100	57
rect	100	56	101	57
rect	101	56	102	57
rect	102	56	103	57
rect	103	56	104	57
rect	104	56	105	57
rect	105	56	106	57
rect	106	56	107	57
rect	107	56	108	57
rect	108	56	109	57
rect	109	56	110	57
rect	111	56	112	57
rect	112	56	113	57
rect	113	56	114	57
rect	114	56	115	57
rect	115	56	116	57
rect	116	56	117	57
rect	117	56	118	57
rect	118	56	119	57
rect	120	56	121	57
rect	121	56	122	57
rect	123	56	124	57
rect	124	56	125	57
rect	125	56	126	57
rect	126	56	127	57
rect	127	56	128	57
rect	129	56	130	57
rect	130	56	131	57
rect	131	56	132	57
rect	132	56	133	57
rect	133	56	134	57
rect	134	56	135	57
rect	135	56	136	57
rect	136	56	137	57
rect	137	56	138	57
rect	138	56	139	57
rect	139	56	140	57
rect	140	56	141	57
rect	141	56	142	57
rect	142	56	143	57
rect	143	56	144	57
rect	144	56	145	57
rect	145	56	146	57
rect	147	56	148	57
rect	148	56	149	57
rect	149	56	150	57
rect	150	56	151	57
rect	151	56	152	57
rect	152	56	153	57
rect	153	56	154	57
rect	154	56	155	57
rect	155	56	156	57
rect	156	56	157	57
rect	157	56	158	57
rect	159	56	160	57
rect	160	56	161	57
rect	162	56	163	57
rect	163	56	164	57
rect	165	56	166	57
rect	166	56	167	57
rect	168	56	169	57
rect	169	56	170	57
rect	171	56	172	57
rect	172	56	173	57
rect	174	56	175	57
rect	175	56	176	57
rect	177	56	178	57
rect	178	56	179	57
rect	192	56	193	57
rect	193	56	194	57
rect	194	56	195	57
rect	195	56	196	57
rect	196	56	197	57
rect	198	56	199	57
rect	199	56	200	57
rect	201	56	202	57
rect	202	56	203	57
rect	204	56	205	57
rect	205	56	206	57
rect	207	56	208	57
rect	208	56	209	57
rect	209	56	210	57
rect	210	56	211	57
rect	211	56	212	57
rect	212	56	213	57
rect	213	56	214	57
rect	214	56	215	57
rect	216	56	217	57
rect	217	56	218	57
rect	219	56	220	57
rect	220	56	221	57
rect	221	56	222	57
rect	222	56	223	57
rect	223	56	224	57
rect	224	56	225	57
rect	225	56	226	57
rect	226	56	227	57
rect	228	56	229	57
rect	229	56	230	57
rect	231	56	232	57
rect	232	56	233	57
rect	234	56	235	57
rect	235	56	236	57
rect	236	56	237	57
rect	237	56	238	57
rect	238	56	239	57
rect	239	56	240	57
rect	241	56	242	57
rect	242	56	243	57
rect	243	56	244	57
rect	250	56	251	57
rect	251	56	252	57
rect	252	56	253	57
rect	257	56	258	57
rect	259	56	260	57
rect	260	56	261	57
rect	262	56	263	57
rect	263	56	264	57
rect	298	56	299	57
rect	299	56	300	57
rect	301	56	302	57
rect	302	56	303	57
rect	303	56	304	57
rect	304	56	305	57
rect	305	56	306	57
rect	15	58	16	59
rect	16	58	17	59
rect	17	58	18	59
rect	18	58	19	59
rect	19	58	20	59
rect	20	58	21	59
rect	31	58	32	59
rect	32	58	33	59
rect	33	58	34	59
rect	35	58	36	59
rect	36	58	37	59
rect	48	58	49	59
rect	49	58	50	59
rect	50	58	51	59
rect	51	58	52	59
rect	52	58	53	59
rect	72	58	73	59
rect	73	58	74	59
rect	74	58	75	59
rect	75	58	76	59
rect	76	58	77	59
rect	77	58	78	59
rect	78	58	79	59
rect	79	58	80	59
rect	81	58	82	59
rect	82	58	83	59
rect	83	58	84	59
rect	84	58	85	59
rect	85	58	86	59
rect	86	58	87	59
rect	87	58	88	59
rect	88	58	89	59
rect	89	58	90	59
rect	90	58	91	59
rect	91	58	92	59
rect	92	58	93	59
rect	93	58	94	59
rect	94	58	95	59
rect	95	58	96	59
rect	96	58	97	59
rect	97	58	98	59
rect	98	58	99	59
rect	99	58	100	59
rect	100	58	101	59
rect	101	58	102	59
rect	102	58	103	59
rect	103	58	104	59
rect	104	58	105	59
rect	105	58	106	59
rect	106	58	107	59
rect	107	58	108	59
rect	108	58	109	59
rect	109	58	110	59
rect	111	58	112	59
rect	112	58	113	59
rect	113	58	114	59
rect	114	58	115	59
rect	115	58	116	59
rect	116	58	117	59
rect	117	58	118	59
rect	118	58	119	59
rect	120	58	121	59
rect	121	58	122	59
rect	123	58	124	59
rect	124	58	125	59
rect	125	58	126	59
rect	126	58	127	59
rect	127	58	128	59
rect	129	58	130	59
rect	130	58	131	59
rect	131	58	132	59
rect	132	58	133	59
rect	133	58	134	59
rect	134	58	135	59
rect	135	58	136	59
rect	136	58	137	59
rect	137	58	138	59
rect	138	58	139	59
rect	139	58	140	59
rect	140	58	141	59
rect	147	58	148	59
rect	148	58	149	59
rect	149	58	150	59
rect	150	58	151	59
rect	151	58	152	59
rect	152	58	153	59
rect	153	58	154	59
rect	154	58	155	59
rect	155	58	156	59
rect	156	58	157	59
rect	157	58	158	59
rect	159	58	160	59
rect	160	58	161	59
rect	162	58	163	59
rect	163	58	164	59
rect	165	58	166	59
rect	166	58	167	59
rect	168	58	169	59
rect	169	58	170	59
rect	171	58	172	59
rect	172	58	173	59
rect	174	58	175	59
rect	175	58	176	59
rect	177	58	178	59
rect	178	58	179	59
rect	180	58	181	59
rect	181	58	182	59
rect	182	58	183	59
rect	183	58	184	59
rect	184	58	185	59
rect	185	58	186	59
rect	186	58	187	59
rect	187	58	188	59
rect	189	58	190	59
rect	190	58	191	59
rect	192	58	193	59
rect	193	58	194	59
rect	194	58	195	59
rect	195	58	196	59
rect	196	58	197	59
rect	198	58	199	59
rect	199	58	200	59
rect	201	58	202	59
rect	202	58	203	59
rect	204	58	205	59
rect	205	58	206	59
rect	207	58	208	59
rect	208	58	209	59
rect	209	58	210	59
rect	210	58	211	59
rect	211	58	212	59
rect	212	58	213	59
rect	213	58	214	59
rect	214	58	215	59
rect	216	58	217	59
rect	217	58	218	59
rect	219	58	220	59
rect	220	58	221	59
rect	221	58	222	59
rect	222	58	223	59
rect	223	58	224	59
rect	224	58	225	59
rect	225	58	226	59
rect	226	58	227	59
rect	228	58	229	59
rect	229	58	230	59
rect	231	58	232	59
rect	232	58	233	59
rect	234	58	235	59
rect	235	58	236	59
rect	236	58	237	59
rect	237	58	238	59
rect	238	58	239	59
rect	239	58	240	59
rect	241	58	242	59
rect	242	58	243	59
rect	243	58	244	59
rect	244	58	245	59
rect	245	58	246	59
rect	247	58	248	59
rect	248	58	249	59
rect	250	58	251	59
rect	251	58	252	59
rect	252	58	253	59
rect	253	58	254	59
rect	254	58	255	59
rect	255	58	256	59
rect	256	58	257	59
rect	257	58	258	59
rect	259	58	260	59
rect	260	58	261	59
rect	262	58	263	59
rect	263	58	264	59
rect	265	58	266	59
rect	266	58	267	59
rect	268	58	269	59
rect	269	58	270	59
rect	271	58	272	59
rect	272	58	273	59
rect	274	58	275	59
rect	275	58	276	59
rect	277	58	278	59
rect	278	58	279	59
rect	280	58	281	59
rect	281	58	282	59
rect	282	58	283	59
rect	283	58	284	59
rect	284	58	285	59
rect	285	58	286	59
rect	286	58	287	59
rect	287	58	288	59
rect	289	58	290	59
rect	290	58	291	59
rect	291	58	292	59
rect	292	58	293	59
rect	293	58	294	59
rect	294	58	295	59
rect	295	58	296	59
rect	296	58	297	59
rect	298	58	299	59
rect	299	58	300	59
rect	301	58	302	59
rect	302	58	303	59
rect	303	58	304	59
rect	304	58	305	59
rect	305	58	306	59
rect	307	58	308	59
rect	308	58	309	59
rect	310	58	311	59
rect	311	58	312	59
rect	312	58	313	59
rect	313	58	314	59
rect	314	58	315	59
rect	315	58	316	59
rect	316	58	317	59
rect	317	58	318	59
rect	322	58	323	59
rect	323	58	324	59
rect	324	58	325	59
rect	325	58	326	59
rect	326	58	327	59
rect	327	58	328	59
rect	328	58	329	59
rect	329	58	330	59
rect	331	58	332	59
rect	332	58	333	59
rect	349	58	350	59
rect	350	58	351	59
rect	351	58	352	59
rect	352	58	353	59
rect	353	58	354	59
rect	358	67	359	68
rect	359	67	360	68
rect	360	67	361	68
rect	361	67	362	68
rect	362	67	363	68
rect	363	67	364	68
rect	364	67	365	68
rect	365	67	366	68
rect	366	67	367	68
rect	367	67	368	68
rect	368	67	369	68
rect	369	67	370	68
rect	370	67	371	68
rect	371	67	372	68
rect	372	67	373	68
rect	373	67	374	68
rect	374	67	375	68
rect	375	67	376	68
rect	376	67	377	68
rect	377	67	378	68
rect	378	67	379	68
rect	379	67	380	68
rect	380	67	381	68
rect	381	67	382	68
rect	382	67	383	68
rect	383	67	384	68
rect	384	67	385	68
rect	385	67	386	68
rect	386	67	387	68
rect	387	67	388	68
rect	388	67	389	68
rect	389	67	390	68
rect	390	67	391	68
rect	391	67	392	68
rect	392	67	393	68
rect	393	67	394	68
rect	394	67	395	68
rect	395	67	396	68
rect	340	69	341	70
rect	341	69	342	70
rect	342	69	343	70
rect	343	69	344	70
rect	344	69	345	70
rect	345	69	346	70
rect	346	69	347	70
rect	347	69	348	70
rect	349	69	350	70
rect	350	69	351	70
rect	351	69	352	70
rect	352	69	353	70
rect	353	69	354	70
rect	354	69	355	70
rect	355	69	356	70
rect	356	69	357	70
rect	331	71	332	72
rect	332	71	333	72
rect	333	71	334	72
rect	334	71	335	72
rect	335	71	336	72
rect	336	71	337	72
rect	337	71	338	72
rect	338	71	339	72
rect	295	73	296	74
rect	296	73	297	74
rect	298	73	299	74
rect	299	73	300	74
rect	301	73	302	74
rect	302	73	303	74
rect	303	73	304	74
rect	304	73	305	74
rect	305	73	306	74
rect	306	73	307	74
rect	307	73	308	74
rect	308	73	309	74
rect	310	73	311	74
rect	311	73	312	74
rect	312	73	313	74
rect	313	73	314	74
rect	314	73	315	74
rect	315	73	316	74
rect	316	73	317	74
rect	317	73	318	74
rect	319	73	320	74
rect	320	73	321	74
rect	322	73	323	74
rect	323	73	324	74
rect	324	73	325	74
rect	325	73	326	74
rect	326	73	327	74
rect	327	73	328	74
rect	328	73	329	74
rect	329	73	330	74
rect	289	75	290	76
rect	290	75	291	76
rect	291	75	292	76
rect	292	75	293	76
rect	293	75	294	76
rect	294	75	295	76
rect	295	75	296	76
rect	296	75	297	76
rect	298	75	299	76
rect	299	75	300	76
rect	301	75	302	76
rect	302	75	303	76
rect	303	75	304	76
rect	304	75	305	76
rect	305	75	306	76
rect	306	75	307	76
rect	307	75	308	76
rect	308	75	309	76
rect	310	75	311	76
rect	311	75	312	76
rect	312	75	313	76
rect	313	75	314	76
rect	314	75	315	76
rect	201	77	202	78
rect	202	77	203	78
rect	204	77	205	78
rect	205	77	206	78
rect	207	77	208	78
rect	208	77	209	78
rect	210	77	211	78
rect	211	77	212	78
rect	212	77	213	78
rect	213	77	214	78
rect	214	77	215	78
rect	216	77	217	78
rect	217	77	218	78
rect	219	77	220	78
rect	220	77	221	78
rect	221	77	222	78
rect	222	77	223	78
rect	223	77	224	78
rect	224	77	225	78
rect	225	77	226	78
rect	226	77	227	78
rect	228	77	229	78
rect	229	77	230	78
rect	231	77	232	78
rect	232	77	233	78
rect	233	77	234	78
rect	234	77	235	78
rect	235	77	236	78
rect	236	77	237	78
rect	237	77	238	78
rect	238	77	239	78
rect	239	77	240	78
rect	240	77	241	78
rect	241	77	242	78
rect	242	77	243	78
rect	243	77	244	78
rect	244	77	245	78
rect	245	77	246	78
rect	247	77	248	78
rect	248	77	249	78
rect	250	77	251	78
rect	251	77	252	78
rect	252	77	253	78
rect	253	77	254	78
rect	254	77	255	78
rect	256	77	257	78
rect	257	77	258	78
rect	259	77	260	78
rect	260	77	261	78
rect	262	77	263	78
rect	263	77	264	78
rect	265	77	266	78
rect	266	77	267	78
rect	268	77	269	78
rect	269	77	270	78
rect	270	77	271	78
rect	271	77	272	78
rect	272	77	273	78
rect	273	77	274	78
rect	274	77	275	78
rect	275	77	276	78
rect	277	77	278	78
rect	278	77	279	78
rect	280	77	281	78
rect	281	77	282	78
rect	282	77	283	78
rect	283	77	284	78
rect	284	77	285	78
rect	285	77	286	78
rect	286	77	287	78
rect	287	77	288	78
rect	288	77	289	78
rect	289	77	290	78
rect	290	77	291	78
rect	291	77	292	78
rect	292	77	293	78
rect	293	77	294	78
rect	294	77	295	78
rect	295	77	296	78
rect	296	77	297	78
rect	298	77	299	78
rect	299	77	300	78
rect	301	77	302	78
rect	302	77	303	78
rect	303	77	304	78
rect	304	77	305	78
rect	305	77	306	78
rect	306	77	307	78
rect	307	77	308	78
rect	308	77	309	78
rect	310	77	311	78
rect	311	77	312	78
rect	312	77	313	78
rect	313	77	314	78
rect	314	77	315	78
rect	316	77	317	78
rect	317	77	318	78
rect	319	77	320	78
rect	320	77	321	78
rect	322	77	323	78
rect	323	77	324	78
rect	168	79	169	80
rect	169	79	170	80
rect	171	79	172	80
rect	172	79	173	80
rect	174	79	175	80
rect	175	79	176	80
rect	177	79	178	80
rect	178	79	179	80
rect	180	79	181	80
rect	181	79	182	80
rect	182	79	183	80
rect	183	79	184	80
rect	184	79	185	80
rect	185	79	186	80
rect	186	79	187	80
rect	187	79	188	80
rect	189	79	190	80
rect	190	79	191	80
rect	191	79	192	80
rect	192	79	193	80
rect	193	79	194	80
rect	195	79	196	80
rect	196	79	197	80
rect	198	79	199	80
rect	199	79	200	80
rect	250	79	251	80
rect	251	79	252	80
rect	265	79	266	80
rect	266	79	267	80
rect	268	79	269	80
rect	269	79	270	80
rect	270	79	271	80
rect	271	79	272	80
rect	272	79	273	80
rect	273	79	274	80
rect	274	79	275	80
rect	275	79	276	80
rect	277	79	278	80
rect	278	79	279	80
rect	280	79	281	80
rect	281	79	282	80
rect	282	79	283	80
rect	283	79	284	80
rect	284	79	285	80
rect	285	79	286	80
rect	286	79	287	80
rect	287	79	288	80
rect	288	79	289	80
rect	289	79	290	80
rect	290	79	291	80
rect	291	79	292	80
rect	292	79	293	80
rect	293	79	294	80
rect	149	81	150	82
rect	150	81	151	82
rect	151	81	152	82
rect	152	81	153	82
rect	153	81	154	82
rect	154	81	155	82
rect	156	81	157	82
rect	157	81	158	82
rect	159	81	160	82
rect	160	81	161	82
rect	162	81	163	82
rect	163	81	164	82
rect	165	81	166	82
rect	166	81	167	82
rect	167	81	168	82
rect	168	81	169	82
rect	169	81	170	82
rect	171	81	172	82
rect	172	81	173	82
rect	174	81	175	82
rect	175	81	176	82
rect	177	81	178	82
rect	178	81	179	82
rect	180	81	181	82
rect	181	81	182	82
rect	182	81	183	82
rect	183	81	184	82
rect	184	81	185	82
rect	185	81	186	82
rect	186	81	187	82
rect	187	81	188	82
rect	228	81	229	82
rect	229	81	230	82
rect	231	81	232	82
rect	232	81	233	82
rect	233	81	234	82
rect	234	81	235	82
rect	235	81	236	82
rect	236	81	237	82
rect	237	81	238	82
rect	238	81	239	82
rect	239	81	240	82
rect	240	81	241	82
rect	241	81	242	82
rect	242	81	243	82
rect	243	81	244	82
rect	244	81	245	82
rect	245	81	246	82
rect	247	81	248	82
rect	248	81	249	82
rect	262	81	263	82
rect	263	81	264	82
rect	264	81	265	82
rect	265	81	266	82
rect	266	81	267	82
rect	268	81	269	82
rect	269	81	270	82
rect	270	81	271	82
rect	271	81	272	82
rect	272	81	273	82
rect	273	81	274	82
rect	274	81	275	82
rect	275	81	276	82
rect	277	81	278	82
rect	278	81	279	82
rect	280	81	281	82
rect	281	81	282	82
rect	282	81	283	82
rect	283	81	284	82
rect	284	81	285	82
rect	285	81	286	82
rect	286	81	287	82
rect	287	81	288	82
rect	288	81	289	82
rect	289	81	290	82
rect	290	81	291	82
rect	165	83	166	84
rect	166	83	167	84
rect	167	83	168	84
rect	168	83	169	84
rect	169	83	170	84
rect	171	83	172	84
rect	172	83	173	84
rect	174	83	175	84
rect	175	83	176	84
rect	177	83	178	84
rect	178	83	179	84
rect	180	83	181	84
rect	181	83	182	84
rect	182	83	183	84
rect	183	83	184	84
rect	184	83	185	84
rect	185	83	186	84
rect	186	83	187	84
rect	187	83	188	84
rect	219	83	220	84
rect	220	83	221	84
rect	221	83	222	84
rect	222	83	223	84
rect	223	83	224	84
rect	224	83	225	84
rect	225	83	226	84
rect	226	83	227	84
rect	227	83	228	84
rect	259	83	260	84
rect	260	83	261	84
rect	261	83	262	84
rect	262	83	263	84
rect	263	83	264	84
rect	264	83	265	84
rect	265	83	266	84
rect	266	83	267	84
rect	268	83	269	84
rect	269	83	270	84
rect	270	83	271	84
rect	271	83	272	84
rect	272	83	273	84
rect	273	83	274	84
rect	274	83	275	84
rect	275	83	276	84
rect	277	83	278	84
rect	278	83	279	84
rect	280	83	281	84
rect	281	83	282	84
rect	282	83	283	84
rect	283	83	284	84
rect	284	83	285	84
rect	285	83	286	84
rect	286	83	287	84
rect	287	83	288	84
rect	162	85	163	86
rect	163	85	164	86
rect	168	85	169	86
rect	169	85	170	86
rect	195	85	196	86
rect	196	85	197	86
rect	198	85	199	86
rect	199	85	200	86
rect	201	85	202	86
rect	202	85	203	86
rect	204	85	205	86
rect	205	85	206	86
rect	207	85	208	86
rect	208	85	209	86
rect	210	85	211	86
rect	211	85	212	86
rect	212	85	213	86
rect	213	85	214	86
rect	214	85	215	86
rect	216	85	217	86
rect	217	85	218	86
rect	218	85	219	86
rect	219	85	220	86
rect	220	85	221	86
rect	221	85	222	86
rect	222	85	223	86
rect	223	85	224	86
rect	224	85	225	86
rect	225	85	226	86
rect	226	85	227	86
rect	227	85	228	86
rect	229	85	230	86
rect	231	85	232	86
rect	232	85	233	86
rect	233	85	234	86
rect	234	85	235	86
rect	235	85	236	86
rect	236	85	237	86
rect	237	85	238	86
rect	238	85	239	86
rect	239	85	240	86
rect	240	85	241	86
rect	241	85	242	86
rect	242	85	243	86
rect	243	85	244	86
rect	244	85	245	86
rect	245	85	246	86
rect	247	85	248	86
rect	248	85	249	86
rect	250	85	251	86
rect	251	85	252	86
rect	253	85	254	86
rect	254	85	255	86
rect	256	85	257	86
rect	257	85	258	86
rect	258	85	259	86
rect	259	85	260	86
rect	260	85	261	86
rect	261	85	262	86
rect	262	85	263	86
rect	263	85	264	86
rect	264	85	265	86
rect	265	85	266	86
rect	266	85	267	86
rect	268	85	269	86
rect	269	85	270	86
rect	298	85	299	86
rect	299	85	300	86
rect	301	85	302	86
rect	302	85	303	86
rect	303	85	304	86
rect	304	85	305	86
rect	305	85	306	86
rect	306	85	307	86
rect	307	85	308	86
rect	308	85	309	86
rect	310	85	311	86
rect	311	85	312	86
rect	312	85	313	86
rect	313	85	314	86
rect	314	85	315	86
rect	316	85	317	86
rect	317	85	318	86
rect	319	85	320	86
rect	320	85	321	86
rect	322	85	323	86
rect	323	85	324	86
rect	325	85	326	86
rect	326	85	327	86
rect	327	85	328	86
rect	328	85	329	86
rect	329	85	330	86
rect	331	85	332	86
rect	332	85	333	86
rect	349	85	350	86
rect	350	85	351	86
rect	351	85	352	86
rect	352	85	353	86
rect	353	85	354	86
rect	354	85	355	86
rect	355	85	356	86
rect	356	85	357	86
rect	358	85	359	86
rect	359	85	360	86
rect	360	85	361	86
rect	361	85	362	86
rect	362	85	363	86
rect	363	85	364	86
rect	364	85	365	86
rect	365	85	366	86
rect	366	85	367	86
rect	367	85	368	86
rect	368	85	369	86
rect	54	87	55	88
rect	55	87	56	88
rect	56	87	57	88
rect	57	87	58	88
rect	58	87	59	88
rect	69	87	70	88
rect	70	87	71	88
rect	78	87	79	88
rect	79	87	80	88
rect	81	87	82	88
rect	82	87	83	88
rect	83	87	84	88
rect	84	87	85	88
rect	85	87	86	88
rect	86	87	87	88
rect	87	87	88	88
rect	88	87	89	88
rect	89	87	90	88
rect	90	87	91	88
rect	91	87	92	88
rect	92	87	93	88
rect	93	87	94	88
rect	94	87	95	88
rect	95	87	96	88
rect	96	87	97	88
rect	97	87	98	88
rect	98	87	99	88
rect	99	87	100	88
rect	100	87	101	88
rect	101	87	102	88
rect	102	87	103	88
rect	103	87	104	88
rect	104	87	105	88
rect	105	87	106	88
rect	106	87	107	88
rect	107	87	108	88
rect	108	87	109	88
rect	109	87	110	88
rect	111	87	112	88
rect	139	87	140	88
rect	140	87	141	88
rect	141	87	142	88
rect	142	87	143	88
rect	143	87	144	88
rect	144	87	145	88
rect	145	87	146	88
rect	146	87	147	88
rect	147	87	148	88
rect	159	87	160	88
rect	160	87	161	88
rect	161	87	162	88
rect	162	87	163	88
rect	163	87	164	88
rect	165	87	166	88
rect	166	87	167	88
rect	168	87	169	88
rect	169	87	170	88
rect	170	87	171	88
rect	171	87	172	88
rect	172	87	173	88
rect	174	87	175	88
rect	175	87	176	88
rect	177	87	178	88
rect	178	87	179	88
rect	180	87	181	88
rect	181	87	182	88
rect	182	87	183	88
rect	183	87	184	88
rect	184	87	185	88
rect	185	87	186	88
rect	186	87	187	88
rect	187	87	188	88
rect	189	87	190	88
rect	190	87	191	88
rect	191	87	192	88
rect	192	87	193	88
rect	193	87	194	88
rect	204	87	205	88
rect	205	87	206	88
rect	207	87	208	88
rect	208	87	209	88
rect	210	87	211	88
rect	211	87	212	88
rect	212	87	213	88
rect	213	87	214	88
rect	214	87	215	88
rect	216	87	217	88
rect	217	87	218	88
rect	218	87	219	88
rect	219	87	220	88
rect	220	87	221	88
rect	221	87	222	88
rect	222	87	223	88
rect	223	87	224	88
rect	224	87	225	88
rect	256	87	257	88
rect	257	87	258	88
rect	258	87	259	88
rect	259	87	260	88
rect	260	87	261	88
rect	261	87	262	88
rect	262	87	263	88
rect	263	87	264	88
rect	264	87	265	88
rect	265	87	266	88
rect	266	87	267	88
rect	268	87	269	88
rect	269	87	270	88
rect	271	87	272	88
rect	272	87	273	88
rect	273	87	274	88
rect	274	87	275	88
rect	275	87	276	88
rect	277	87	278	88
rect	278	87	279	88
rect	280	87	281	88
rect	281	87	282	88
rect	282	87	283	88
rect	283	87	284	88
rect	284	87	285	88
rect	285	87	286	88
rect	286	87	287	88
rect	287	87	288	88
rect	289	87	290	88
rect	290	87	291	88
rect	292	87	293	88
rect	293	87	294	88
rect	295	87	296	88
rect	296	87	297	88
rect	297	87	298	88
rect	298	87	299	88
rect	299	87	300	88
rect	301	87	302	88
rect	302	87	303	88
rect	303	87	304	88
rect	304	87	305	88
rect	305	87	306	88
rect	319	87	320	88
rect	320	87	321	88
rect	322	87	323	88
rect	323	87	324	88
rect	325	87	326	88
rect	326	87	327	88
rect	327	87	328	88
rect	328	87	329	88
rect	329	87	330	88
rect	331	87	332	88
rect	332	87	333	88
rect	334	87	335	88
rect	335	87	336	88
rect	336	87	337	88
rect	337	87	338	88
rect	338	87	339	88
rect	340	87	341	88
rect	341	87	342	88
rect	342	87	343	88
rect	343	87	344	88
rect	344	87	345	88
rect	345	87	346	88
rect	346	87	347	88
rect	347	87	348	88
rect	38	89	39	90
rect	39	89	40	90
rect	51	89	52	90
rect	52	89	53	90
rect	53	89	54	90
rect	54	89	55	90
rect	55	89	56	90
rect	56	89	57	90
rect	57	89	58	90
rect	58	89	59	90
rect	60	89	61	90
rect	61	89	62	90
rect	63	89	64	90
rect	64	89	65	90
rect	65	89	66	90
rect	66	89	67	90
rect	67	89	68	90
rect	69	89	70	90
rect	70	89	71	90
rect	71	89	72	90
rect	72	89	73	90
rect	73	89	74	90
rect	74	89	75	90
rect	75	89	76	90
rect	76	89	77	90
rect	77	89	78	90
rect	78	89	79	90
rect	79	89	80	90
rect	81	89	82	90
rect	82	89	83	90
rect	83	89	84	90
rect	84	89	85	90
rect	85	89	86	90
rect	86	89	87	90
rect	87	89	88	90
rect	88	89	89	90
rect	89	89	90	90
rect	90	89	91	90
rect	91	89	92	90
rect	92	89	93	90
rect	93	89	94	90
rect	94	89	95	90
rect	95	89	96	90
rect	96	89	97	90
rect	97	89	98	90
rect	98	89	99	90
rect	99	89	100	90
rect	100	89	101	90
rect	101	89	102	90
rect	102	89	103	90
rect	103	89	104	90
rect	104	89	105	90
rect	105	89	106	90
rect	106	89	107	90
rect	107	89	108	90
rect	108	89	109	90
rect	109	89	110	90
rect	111	89	112	90
rect	113	89	114	90
rect	114	89	115	90
rect	115	89	116	90
rect	116	89	117	90
rect	117	89	118	90
rect	118	89	119	90
rect	120	89	121	90
rect	121	89	122	90
rect	122	89	123	90
rect	123	89	124	90
rect	124	89	125	90
rect	125	89	126	90
rect	126	89	127	90
rect	127	89	128	90
rect	129	89	130	90
rect	130	89	131	90
rect	131	89	132	90
rect	132	89	133	90
rect	133	89	134	90
rect	134	89	135	90
rect	135	89	136	90
rect	136	89	137	90
rect	137	89	138	90
rect	138	89	139	90
rect	139	89	140	90
rect	140	89	141	90
rect	141	89	142	90
rect	142	89	143	90
rect	143	89	144	90
rect	144	89	145	90
rect	145	89	146	90
rect	146	89	147	90
rect	147	89	148	90
rect	149	89	150	90
rect	150	89	151	90
rect	151	89	152	90
rect	152	89	153	90
rect	153	89	154	90
rect	154	89	155	90
rect	156	89	157	90
rect	157	89	158	90
rect	158	89	159	90
rect	159	89	160	90
rect	160	89	161	90
rect	161	89	162	90
rect	162	89	163	90
rect	163	89	164	90
rect	165	89	166	90
rect	166	89	167	90
rect	168	89	169	90
rect	169	89	170	90
rect	170	89	171	90
rect	171	89	172	90
rect	172	89	173	90
rect	174	89	175	90
rect	175	89	176	90
rect	177	89	178	90
rect	178	89	179	90
rect	180	89	181	90
rect	181	89	182	90
rect	182	89	183	90
rect	183	89	184	90
rect	184	89	185	90
rect	185	89	186	90
rect	186	89	187	90
rect	187	89	188	90
rect	189	89	190	90
rect	190	89	191	90
rect	191	89	192	90
rect	192	89	193	90
rect	193	89	194	90
rect	195	89	196	90
rect	196	89	197	90
rect	198	89	199	90
rect	199	89	200	90
rect	201	89	202	90
rect	202	89	203	90
rect	216	89	217	90
rect	217	89	218	90
rect	218	89	219	90
rect	231	89	232	90
rect	232	89	233	90
rect	233	89	234	90
rect	234	89	235	90
rect	235	89	236	90
rect	236	89	237	90
rect	237	89	238	90
rect	238	89	239	90
rect	239	89	240	90
rect	240	89	241	90
rect	241	89	242	90
rect	242	89	243	90
rect	243	89	244	90
rect	244	89	245	90
rect	245	89	246	90
rect	247	89	248	90
rect	248	89	249	90
rect	250	89	251	90
rect	251	89	252	90
rect	253	89	254	90
rect	254	89	255	90
rect	255	89	256	90
rect	256	89	257	90
rect	257	89	258	90
rect	258	89	259	90
rect	259	89	260	90
rect	260	89	261	90
rect	261	89	262	90
rect	262	89	263	90
rect	263	89	264	90
rect	277	89	278	90
rect	278	89	279	90
rect	280	89	281	90
rect	281	89	282	90
rect	282	89	283	90
rect	283	89	284	90
rect	284	89	285	90
rect	285	89	286	90
rect	286	89	287	90
rect	287	89	288	90
rect	289	89	290	90
rect	290	89	291	90
rect	292	89	293	90
rect	293	89	294	90
rect	295	89	296	90
rect	296	89	297	90
rect	319	89	320	90
rect	320	89	321	90
rect	35	91	36	92
rect	36	91	37	92
rect	51	91	52	92
rect	52	91	53	92
rect	53	91	54	92
rect	54	91	55	92
rect	55	91	56	92
rect	63	91	64	92
rect	64	91	65	92
rect	65	91	66	92
rect	66	91	67	92
rect	67	91	68	92
rect	69	91	70	92
rect	70	91	71	92
rect	71	91	72	92
rect	72	91	73	92
rect	73	91	74	92
rect	74	91	75	92
rect	75	91	76	92
rect	76	91	77	92
rect	81	91	82	92
rect	82	91	83	92
rect	83	91	84	92
rect	84	91	85	92
rect	85	91	86	92
rect	120	91	121	92
rect	121	91	122	92
rect	122	91	123	92
rect	123	91	124	92
rect	124	91	125	92
rect	125	91	126	92
rect	126	91	127	92
rect	127	91	128	92
rect	129	91	130	92
rect	137	91	138	92
rect	138	91	139	92
rect	143	91	144	92
rect	144	91	145	92
rect	145	91	146	92
rect	146	91	147	92
rect	147	91	148	92
rect	149	91	150	92
rect	150	91	151	92
rect	151	91	152	92
rect	152	91	153	92
rect	153	91	154	92
rect	154	91	155	92
rect	156	91	157	92
rect	157	91	158	92
rect	158	91	159	92
rect	159	91	160	92
rect	160	91	161	92
rect	161	91	162	92
rect	162	91	163	92
rect	163	91	164	92
rect	165	91	166	92
rect	166	91	167	92
rect	168	91	169	92
rect	169	91	170	92
rect	170	91	171	92
rect	171	91	172	92
rect	172	91	173	92
rect	174	91	175	92
rect	175	91	176	92
rect	177	91	178	92
rect	178	91	179	92
rect	180	91	181	92
rect	181	91	182	92
rect	182	91	183	92
rect	183	91	184	92
rect	184	91	185	92
rect	185	91	186	92
rect	186	91	187	92
rect	187	91	188	92
rect	189	91	190	92
rect	190	91	191	92
rect	191	91	192	92
rect	192	91	193	92
rect	193	91	194	92
rect	195	91	196	92
rect	196	91	197	92
rect	198	91	199	92
rect	199	91	200	92
rect	201	91	202	92
rect	202	91	203	92
rect	204	91	205	92
rect	205	91	206	92
rect	207	91	208	92
rect	208	91	209	92
rect	210	91	211	92
rect	211	91	212	92
rect	212	91	213	92
rect	213	91	214	92
rect	214	91	215	92
rect	215	91	216	92
rect	216	91	217	92
rect	217	91	218	92
rect	218	91	219	92
rect	220	91	221	92
rect	221	91	222	92
rect	222	91	223	92
rect	223	91	224	92
rect	224	91	225	92
rect	226	91	227	92
rect	227	91	228	92
rect	229	91	230	92
rect	230	91	231	92
rect	231	91	232	92
rect	232	91	233	92
rect	233	91	234	92
rect	234	91	235	92
rect	235	91	236	92
rect	236	91	237	92
rect	237	91	238	92
rect	238	91	239	92
rect	239	91	240	92
rect	240	91	241	92
rect	241	91	242	92
rect	242	91	243	92
rect	243	91	244	92
rect	244	91	245	92
rect	245	91	246	92
rect	247	91	248	92
rect	248	91	249	92
rect	250	91	251	92
rect	251	91	252	92
rect	253	91	254	92
rect	254	91	255	92
rect	255	91	256	92
rect	256	91	257	92
rect	257	91	258	92
rect	258	91	259	92
rect	259	91	260	92
rect	260	91	261	92
rect	261	91	262	92
rect	262	91	263	92
rect	263	91	264	92
rect	265	91	266	92
rect	266	91	267	92
rect	268	91	269	92
rect	269	91	270	92
rect	271	91	272	92
rect	272	91	273	92
rect	273	91	274	92
rect	274	91	275	92
rect	275	91	276	92
rect	276	91	277	92
rect	277	91	278	92
rect	278	91	279	92
rect	280	91	281	92
rect	281	91	282	92
rect	282	91	283	92
rect	283	91	284	92
rect	284	91	285	92
rect	285	91	286	92
rect	286	91	287	92
rect	287	91	288	92
rect	289	91	290	92
rect	290	91	291	92
rect	292	91	293	92
rect	293	91	294	92
rect	295	91	296	92
rect	296	91	297	92
rect	298	91	299	92
rect	299	91	300	92
rect	301	91	302	92
rect	302	91	303	92
rect	303	91	304	92
rect	304	91	305	92
rect	305	91	306	92
rect	307	91	308	92
rect	308	91	309	92
rect	310	91	311	92
rect	311	91	312	92
rect	312	91	313	92
rect	313	91	314	92
rect	314	91	315	92
rect	316	91	317	92
rect	317	91	318	92
rect	319	91	320	92
rect	320	91	321	92
rect	321	91	322	92
rect	322	91	323	92
rect	323	91	324	92
rect	325	91	326	92
rect	326	91	327	92
rect	327	91	328	92
rect	328	91	329	92
rect	329	91	330	92
rect	331	91	332	92
rect	332	91	333	92
rect	334	91	335	92
rect	335	91	336	92
rect	336	91	337	92
rect	337	91	338	92
rect	338	91	339	92
rect	340	91	341	92
rect	341	91	342	92
rect	342	91	343	92
rect	343	91	344	92
rect	344	91	345	92
rect	345	91	346	92
rect	346	91	347	92
rect	347	91	348	92
rect	349	91	350	92
rect	350	91	351	92
rect	351	91	352	92
rect	352	91	353	92
rect	353	91	354	92
rect	354	91	355	92
rect	355	91	356	92
rect	356	91	357	92
rect	358	91	359	92
rect	359	91	360	92
rect	22	93	23	94
rect	23	93	24	94
rect	24	93	25	94
rect	25	93	26	94
rect	26	93	27	94
rect	27	93	28	94
rect	32	93	33	94
rect	33	93	34	94
rect	35	93	36	94
rect	36	93	37	94
rect	38	93	39	94
rect	39	93	40	94
rect	41	93	42	94
rect	42	93	43	94
rect	43	93	44	94
rect	44	93	45	94
rect	45	93	46	94
rect	46	93	47	94
rect	47	93	48	94
rect	48	93	49	94
rect	49	93	50	94
rect	51	93	52	94
rect	52	93	53	94
rect	53	93	54	94
rect	54	93	55	94
rect	55	93	56	94
rect	57	93	58	94
rect	58	93	59	94
rect	60	93	61	94
rect	61	93	62	94
rect	62	93	63	94
rect	63	93	64	94
rect	64	93	65	94
rect	65	93	66	94
rect	66	93	67	94
rect	67	93	68	94
rect	69	93	70	94
rect	70	93	71	94
rect	71	93	72	94
rect	72	93	73	94
rect	73	93	74	94
rect	74	93	75	94
rect	75	93	76	94
rect	76	93	77	94
rect	78	93	79	94
rect	79	93	80	94
rect	80	93	81	94
rect	81	93	82	94
rect	82	93	83	94
rect	83	93	84	94
rect	84	93	85	94
rect	85	93	86	94
rect	87	93	88	94
rect	88	93	89	94
rect	111	93	112	94
rect	113	93	114	94
rect	114	93	115	94
rect	115	93	116	94
rect	116	93	117	94
rect	117	93	118	94
rect	118	93	119	94
rect	119	93	120	94
rect	120	93	121	94
rect	129	93	130	94
rect	131	93	132	94
rect	132	93	133	94
rect	133	93	134	94
rect	134	93	135	94
rect	135	93	136	94
rect	137	93	138	94
rect	138	93	139	94
rect	140	93	141	94
rect	141	93	142	94
rect	143	93	144	94
rect	144	93	145	94
rect	145	93	146	94
rect	146	93	147	94
rect	147	93	148	94
rect	149	93	150	94
rect	150	93	151	94
rect	156	93	157	94
rect	157	93	158	94
rect	158	93	159	94
rect	159	93	160	94
rect	160	93	161	94
rect	161	93	162	94
rect	162	93	163	94
rect	163	93	164	94
rect	165	93	166	94
rect	166	93	167	94
rect	168	93	169	94
rect	169	93	170	94
rect	170	93	171	94
rect	171	93	172	94
rect	172	93	173	94
rect	174	93	175	94
rect	175	93	176	94
rect	177	93	178	94
rect	178	93	179	94
rect	180	93	181	94
rect	181	93	182	94
rect	182	93	183	94
rect	183	93	184	94
rect	184	93	185	94
rect	185	93	186	94
rect	186	93	187	94
rect	187	93	188	94
rect	189	93	190	94
rect	190	93	191	94
rect	198	93	199	94
rect	199	93	200	94
rect	201	93	202	94
rect	202	93	203	94
rect	204	93	205	94
rect	205	93	206	94
rect	207	93	208	94
rect	208	93	209	94
rect	210	93	211	94
rect	211	93	212	94
rect	212	93	213	94
rect	213	93	214	94
rect	214	93	215	94
rect	215	93	216	94
rect	216	93	217	94
rect	217	93	218	94
rect	218	93	219	94
rect	220	93	221	94
rect	221	93	222	94
rect	232	93	233	94
rect	233	93	234	94
rect	234	93	235	94
rect	235	93	236	94
rect	236	93	237	94
rect	237	93	238	94
rect	238	93	239	94
rect	239	93	240	94
rect	240	93	241	94
rect	241	93	242	94
rect	242	93	243	94
rect	243	93	244	94
rect	244	93	245	94
rect	245	93	246	94
rect	247	93	248	94
rect	248	93	249	94
rect	250	93	251	94
rect	251	93	252	94
rect	253	93	254	94
rect	254	93	255	94
rect	259	93	260	94
rect	260	93	261	94
rect	268	93	269	94
rect	269	93	270	94
rect	271	93	272	94
rect	272	93	273	94
rect	277	93	278	94
rect	278	93	279	94
rect	310	93	311	94
rect	311	93	312	94
rect	312	93	313	94
rect	313	93	314	94
rect	314	93	315	94
rect	316	93	317	94
rect	317	93	318	94
rect	319	93	320	94
rect	320	93	321	94
rect	12	95	13	96
rect	13	95	14	96
rect	14	95	15	96
rect	15	95	16	96
rect	16	95	17	96
rect	17	95	18	96
rect	18	95	19	96
rect	19	95	20	96
rect	20	95	21	96
rect	21	95	22	96
rect	22	95	23	96
rect	23	95	24	96
rect	24	95	25	96
rect	25	95	26	96
rect	26	95	27	96
rect	27	95	28	96
rect	29	95	30	96
rect	30	95	31	96
rect	32	95	33	96
rect	33	95	34	96
rect	35	95	36	96
rect	36	95	37	96
rect	38	95	39	96
rect	39	95	40	96
rect	41	95	42	96
rect	42	95	43	96
rect	43	95	44	96
rect	44	95	45	96
rect	45	95	46	96
rect	46	95	47	96
rect	47	95	48	96
rect	48	95	49	96
rect	49	95	50	96
rect	51	95	52	96
rect	52	95	53	96
rect	53	95	54	96
rect	54	95	55	96
rect	55	95	56	96
rect	57	95	58	96
rect	58	95	59	96
rect	60	95	61	96
rect	61	95	62	96
rect	62	95	63	96
rect	63	95	64	96
rect	64	95	65	96
rect	65	95	66	96
rect	66	95	67	96
rect	67	95	68	96
rect	69	95	70	96
rect	70	95	71	96
rect	71	95	72	96
rect	72	95	73	96
rect	73	95	74	96
rect	74	95	75	96
rect	75	95	76	96
rect	76	95	77	96
rect	78	95	79	96
rect	79	95	80	96
rect	80	95	81	96
rect	81	95	82	96
rect	82	95	83	96
rect	83	95	84	96
rect	84	95	85	96
rect	85	95	86	96
rect	87	95	88	96
rect	88	95	89	96
rect	90	95	91	96
rect	91	95	92	96
rect	92	95	93	96
rect	93	95	94	96
rect	94	95	95	96
rect	95	95	96	96
rect	96	95	97	96
rect	97	95	98	96
rect	98	95	99	96
rect	99	95	100	96
rect	100	95	101	96
rect	101	95	102	96
rect	102	95	103	96
rect	103	95	104	96
rect	104	95	105	96
rect	105	95	106	96
rect	106	95	107	96
rect	107	95	108	96
rect	108	95	109	96
rect	109	95	110	96
rect	110	95	111	96
rect	111	95	112	96
rect	113	95	114	96
rect	114	95	115	96
rect	115	95	116	96
rect	116	95	117	96
rect	117	95	118	96
rect	118	95	119	96
rect	119	95	120	96
rect	120	95	121	96
rect	122	95	123	96
rect	123	95	124	96
rect	124	95	125	96
rect	125	95	126	96
rect	126	95	127	96
rect	127	95	128	96
rect	128	95	129	96
rect	129	95	130	96
rect	131	95	132	96
rect	132	95	133	96
rect	133	95	134	96
rect	134	95	135	96
rect	135	95	136	96
rect	137	95	138	96
rect	138	95	139	96
rect	140	95	141	96
rect	141	95	142	96
rect	143	95	144	96
rect	144	95	145	96
rect	145	95	146	96
rect	146	95	147	96
rect	147	95	148	96
rect	149	95	150	96
rect	150	95	151	96
rect	152	95	153	96
rect	153	95	154	96
rect	154	95	155	96
rect	155	95	156	96
rect	156	95	157	96
rect	157	95	158	96
rect	158	95	159	96
rect	159	95	160	96
rect	160	95	161	96
rect	161	95	162	96
rect	162	95	163	96
rect	163	95	164	96
rect	165	95	166	96
rect	166	95	167	96
rect	168	95	169	96
rect	169	95	170	96
rect	198	95	199	96
rect	199	95	200	96
rect	201	95	202	96
rect	202	95	203	96
rect	204	95	205	96
rect	205	95	206	96
rect	210	95	211	96
rect	211	95	212	96
rect	212	95	213	96
rect	213	95	214	96
rect	214	95	215	96
rect	215	95	216	96
rect	216	95	217	96
rect	217	95	218	96
rect	218	95	219	96
rect	220	95	221	96
rect	221	95	222	96
rect	223	95	224	96
rect	224	95	225	96
rect	226	95	227	96
rect	227	95	228	96
rect	229	95	230	96
rect	230	95	231	96
rect	232	95	233	96
rect	233	95	234	96
rect	234	95	235	96
rect	235	95	236	96
rect	236	95	237	96
rect	237	95	238	96
rect	238	95	239	96
rect	239	95	240	96
rect	247	95	248	96
rect	248	95	249	96
rect	250	95	251	96
rect	251	95	252	96
rect	253	95	254	96
rect	254	95	255	96
rect	256	95	257	96
rect	257	95	258	96
rect	259	95	260	96
rect	260	95	261	96
rect	262	95	263	96
rect	263	95	264	96
rect	265	95	266	96
rect	266	95	267	96
rect	280	95	281	96
rect	281	95	282	96
rect	282	95	283	96
rect	283	95	284	96
rect	284	95	285	96
rect	301	95	302	96
rect	302	95	303	96
rect	303	95	304	96
rect	304	95	305	96
rect	305	95	306	96
rect	307	95	308	96
rect	308	95	309	96
rect	309	95	310	96
rect	310	95	311	96
rect	311	95	312	96
rect	312	95	313	96
rect	313	95	314	96
rect	314	95	315	96
rect	316	95	317	96
rect	317	95	318	96
rect	319	95	320	96
rect	320	95	321	96
rect	322	95	323	96
rect	323	95	324	96
rect	325	95	326	96
rect	326	95	327	96
rect	327	95	328	96
rect	328	95	329	96
rect	329	95	330	96
rect	331	95	332	96
rect	332	95	333	96
rect	334	95	335	96
rect	335	95	336	96
rect	379	95	380	96
rect	380	95	381	96
rect	385	95	386	96
rect	386	95	387	96
rect	214	104	215	105
rect	215	104	216	105
rect	216	104	217	105
rect	217	104	218	105
rect	218	104	219	105
rect	340	104	341	105
rect	341	104	342	105
rect	379	104	380	105
rect	380	104	381	105
rect	381	104	382	105
rect	382	104	383	105
rect	383	104	384	105
rect	384	104	385	105
rect	385	104	386	105
rect	386	104	387	105
rect	388	104	389	105
rect	389	104	390	105
rect	390	104	391	105
rect	391	104	392	105
rect	392	104	393	105
rect	393	104	394	105
rect	394	104	395	105
rect	395	104	396	105
rect	397	104	398	105
rect	398	104	399	105
rect	399	104	400	105
rect	400	104	401	105
rect	401	104	402	105
rect	403	104	404	105
rect	404	104	405	105
rect	405	104	406	105
rect	406	104	407	105
rect	407	104	408	105
rect	408	104	409	105
rect	409	104	410	105
rect	410	104	411	105
rect	411	104	412	105
rect	412	104	413	105
rect	413	104	414	105
rect	414	104	415	105
rect	415	104	416	105
rect	416	104	417	105
rect	417	104	418	105
rect	418	104	419	105
rect	204	106	205	107
rect	205	106	206	107
rect	206	106	207	107
rect	207	106	208	107
rect	208	106	209	107
rect	209	106	210	107
rect	210	106	211	107
rect	211	106	212	107
rect	212	106	213	107
rect	213	106	214	107
rect	214	106	215	107
rect	215	106	216	107
rect	216	106	217	107
rect	217	106	218	107
rect	218	106	219	107
rect	268	106	269	107
rect	269	106	270	107
rect	271	106	272	107
rect	272	106	273	107
rect	274	106	275	107
rect	275	106	276	107
rect	277	106	278	107
rect	278	106	279	107
rect	298	106	299	107
rect	299	106	300	107
rect	301	106	302	107
rect	302	106	303	107
rect	331	106	332	107
rect	332	106	333	107
rect	334	106	335	107
rect	335	106	336	107
rect	337	106	338	107
rect	338	106	339	107
rect	339	106	340	107
rect	340	106	341	107
rect	341	106	342	107
rect	343	106	344	107
rect	344	106	345	107
rect	346	106	347	107
rect	347	106	348	107
rect	349	106	350	107
rect	350	106	351	107
rect	352	106	353	107
rect	353	106	354	107
rect	354	106	355	107
rect	355	106	356	107
rect	356	106	357	107
rect	358	106	359	107
rect	359	106	360	107
rect	361	106	362	107
rect	362	106	363	107
rect	363	106	364	107
rect	364	106	365	107
rect	365	106	366	107
rect	366	106	367	107
rect	367	106	368	107
rect	368	106	369	107
rect	370	106	371	107
rect	371	106	372	107
rect	372	106	373	107
rect	373	106	374	107
rect	374	106	375	107
rect	375	106	376	107
rect	376	106	377	107
rect	377	106	378	107
rect	378	106	379	107
rect	379	106	380	107
rect	380	106	381	107
rect	381	106	382	107
rect	382	106	383	107
rect	383	106	384	107
rect	384	106	385	107
rect	385	106	386	107
rect	386	106	387	107
rect	388	106	389	107
rect	389	106	390	107
rect	390	106	391	107
rect	391	106	392	107
rect	392	106	393	107
rect	393	106	394	107
rect	394	106	395	107
rect	395	106	396	107
rect	397	106	398	107
rect	398	106	399	107
rect	399	106	400	107
rect	400	106	401	107
rect	401	106	402	107
rect	186	108	187	109
rect	187	108	188	109
rect	189	108	190	109
rect	190	108	191	109
rect	192	108	193	109
rect	193	108	194	109
rect	195	108	196	109
rect	196	108	197	109
rect	198	108	199	109
rect	199	108	200	109
rect	201	108	202	109
rect	202	108	203	109
rect	203	108	204	109
rect	262	108	263	109
rect	263	108	264	109
rect	265	108	266	109
rect	266	108	267	109
rect	267	108	268	109
rect	268	108	269	109
rect	269	108	270	109
rect	271	108	272	109
rect	272	108	273	109
rect	274	108	275	109
rect	275	108	276	109
rect	277	108	278	109
rect	278	108	279	109
rect	280	108	281	109
rect	281	108	282	109
rect	282	108	283	109
rect	283	108	284	109
rect	284	108	285	109
rect	286	108	287	109
rect	287	108	288	109
rect	289	108	290	109
rect	290	108	291	109
rect	292	108	293	109
rect	293	108	294	109
rect	295	108	296	109
rect	296	108	297	109
rect	301	108	302	109
rect	302	108	303	109
rect	304	108	305	109
rect	305	108	306	109
rect	337	108	338	109
rect	338	108	339	109
rect	339	108	340	109
rect	340	108	341	109
rect	341	108	342	109
rect	343	108	344	109
rect	344	108	345	109
rect	346	108	347	109
rect	347	108	348	109
rect	349	108	350	109
rect	350	108	351	109
rect	352	108	353	109
rect	353	108	354	109
rect	354	108	355	109
rect	355	108	356	109
rect	356	108	357	109
rect	358	108	359	109
rect	359	108	360	109
rect	361	108	362	109
rect	362	108	363	109
rect	363	108	364	109
rect	364	108	365	109
rect	365	108	366	109
rect	366	108	367	109
rect	367	108	368	109
rect	368	108	369	109
rect	370	108	371	109
rect	371	108	372	109
rect	372	108	373	109
rect	373	108	374	109
rect	374	108	375	109
rect	375	108	376	109
rect	376	108	377	109
rect	377	108	378	109
rect	388	108	389	109
rect	389	108	390	109
rect	390	108	391	109
rect	391	108	392	109
rect	392	108	393	109
rect	393	108	394	109
rect	394	108	395	109
rect	395	108	396	109
rect	397	108	398	109
rect	398	108	399	109
rect	399	108	400	109
rect	400	108	401	109
rect	401	108	402	109
rect	184	110	185	111
rect	185	110	186	111
rect	186	110	187	111
rect	187	110	188	111
rect	192	110	193	111
rect	193	110	194	111
rect	195	110	196	111
rect	196	110	197	111
rect	198	110	199	111
rect	199	110	200	111
rect	201	110	202	111
rect	202	110	203	111
rect	203	110	204	111
rect	205	110	206	111
rect	206	110	207	111
rect	207	110	208	111
rect	208	110	209	111
rect	209	110	210	111
rect	210	110	211	111
rect	211	110	212	111
rect	212	110	213	111
rect	250	110	251	111
rect	251	110	252	111
rect	253	110	254	111
rect	254	110	255	111
rect	255	110	256	111
rect	256	110	257	111
rect	257	110	258	111
rect	259	110	260	111
rect	260	110	261	111
rect	265	110	266	111
rect	266	110	267	111
rect	267	110	268	111
rect	268	110	269	111
rect	269	110	270	111
rect	271	110	272	111
rect	272	110	273	111
rect	274	110	275	111
rect	275	110	276	111
rect	277	110	278	111
rect	278	110	279	111
rect	280	110	281	111
rect	281	110	282	111
rect	282	110	283	111
rect	283	110	284	111
rect	284	110	285	111
rect	286	110	287	111
rect	287	110	288	111
rect	289	110	290	111
rect	290	110	291	111
rect	292	110	293	111
rect	293	110	294	111
rect	295	110	296	111
rect	296	110	297	111
rect	298	110	299	111
rect	299	110	300	111
rect	300	110	301	111
rect	301	110	302	111
rect	302	110	303	111
rect	304	110	305	111
rect	305	110	306	111
rect	306	110	307	111
rect	307	110	308	111
rect	308	110	309	111
rect	309	110	310	111
rect	310	110	311	111
rect	311	110	312	111
rect	322	110	323	111
rect	323	110	324	111
rect	324	110	325	111
rect	325	110	326	111
rect	326	110	327	111
rect	328	110	329	111
rect	329	110	330	111
rect	330	110	331	111
rect	331	110	332	111
rect	332	110	333	111
rect	334	110	335	111
rect	335	110	336	111
rect	336	110	337	111
rect	337	110	338	111
rect	338	110	339	111
rect	352	110	353	111
rect	353	110	354	111
rect	354	110	355	111
rect	355	110	356	111
rect	356	110	357	111
rect	358	110	359	111
rect	359	110	360	111
rect	361	110	362	111
rect	362	110	363	111
rect	363	110	364	111
rect	364	110	365	111
rect	365	110	366	111
rect	366	110	367	111
rect	367	110	368	111
rect	368	110	369	111
rect	370	110	371	111
rect	371	110	372	111
rect	372	110	373	111
rect	373	110	374	111
rect	374	110	375	111
rect	375	110	376	111
rect	376	110	377	111
rect	377	110	378	111
rect	379	110	380	111
rect	380	110	381	111
rect	381	110	382	111
rect	382	110	383	111
rect	383	110	384	111
rect	384	110	385	111
rect	385	110	386	111
rect	386	110	387	111
rect	174	112	175	113
rect	175	112	176	113
rect	177	112	178	113
rect	178	112	179	113
rect	180	112	181	113
rect	181	112	182	113
rect	182	112	183	113
rect	184	112	185	113
rect	185	112	186	113
rect	186	112	187	113
rect	187	112	188	113
rect	188	112	189	113
rect	195	112	196	113
rect	196	112	197	113
rect	198	112	199	113
rect	199	112	200	113
rect	201	112	202	113
rect	202	112	203	113
rect	203	112	204	113
rect	205	112	206	113
rect	206	112	207	113
rect	207	112	208	113
rect	208	112	209	113
rect	209	112	210	113
rect	210	112	211	113
rect	211	112	212	113
rect	212	112	213	113
rect	214	112	215	113
rect	215	112	216	113
rect	223	112	224	113
rect	224	112	225	113
rect	226	112	227	113
rect	227	112	228	113
rect	229	112	230	113
rect	230	112	231	113
rect	232	112	233	113
rect	233	112	234	113
rect	234	112	235	113
rect	235	112	236	113
rect	236	112	237	113
rect	238	112	239	113
rect	239	112	240	113
rect	241	112	242	113
rect	242	112	243	113
rect	247	112	248	113
rect	248	112	249	113
rect	249	112	250	113
rect	250	112	251	113
rect	251	112	252	113
rect	265	112	266	113
rect	266	112	267	113
rect	267	112	268	113
rect	268	112	269	113
rect	269	112	270	113
rect	271	112	272	113
rect	272	112	273	113
rect	274	112	275	113
rect	275	112	276	113
rect	295	112	296	113
rect	296	112	297	113
rect	298	112	299	113
rect	299	112	300	113
rect	300	112	301	113
rect	301	112	302	113
rect	302	112	303	113
rect	304	112	305	113
rect	305	112	306	113
rect	306	112	307	113
rect	307	112	308	113
rect	308	112	309	113
rect	309	112	310	113
rect	310	112	311	113
rect	311	112	312	113
rect	313	112	314	113
rect	314	112	315	113
rect	316	112	317	113
rect	317	112	318	113
rect	319	112	320	113
rect	320	112	321	113
rect	321	112	322	113
rect	322	112	323	113
rect	323	112	324	113
rect	324	112	325	113
rect	325	112	326	113
rect	326	112	327	113
rect	328	112	329	113
rect	329	112	330	113
rect	330	112	331	113
rect	331	112	332	113
rect	332	112	333	113
rect	334	112	335	113
rect	335	112	336	113
rect	336	112	337	113
rect	337	112	338	113
rect	338	112	339	113
rect	340	112	341	113
rect	341	112	342	113
rect	343	112	344	113
rect	344	112	345	113
rect	346	112	347	113
rect	347	112	348	113
rect	349	112	350	113
rect	350	112	351	113
rect	358	112	359	113
rect	359	112	360	113
rect	361	112	362	113
rect	362	112	363	113
rect	363	112	364	113
rect	364	112	365	113
rect	365	112	366	113
rect	366	112	367	113
rect	367	112	368	113
rect	368	112	369	113
rect	370	112	371	113
rect	371	112	372	113
rect	152	114	153	115
rect	153	114	154	115
rect	154	114	155	115
rect	155	114	156	115
rect	156	114	157	115
rect	157	114	158	115
rect	158	114	159	115
rect	159	114	160	115
rect	160	114	161	115
rect	161	114	162	115
rect	162	114	163	115
rect	163	114	164	115
rect	164	114	165	115
rect	165	114	166	115
rect	166	114	167	115
rect	168	114	169	115
rect	169	114	170	115
rect	171	114	172	115
rect	172	114	173	115
rect	173	114	174	115
rect	180	114	181	115
rect	181	114	182	115
rect	182	114	183	115
rect	184	114	185	115
rect	185	114	186	115
rect	186	114	187	115
rect	187	114	188	115
rect	188	114	189	115
rect	190	114	191	115
rect	191	114	192	115
rect	192	114	193	115
rect	193	114	194	115
rect	194	114	195	115
rect	201	114	202	115
rect	202	114	203	115
rect	203	114	204	115
rect	205	114	206	115
rect	206	114	207	115
rect	207	114	208	115
rect	208	114	209	115
rect	209	114	210	115
rect	210	114	211	115
rect	211	114	212	115
rect	212	114	213	115
rect	214	114	215	115
rect	215	114	216	115
rect	217	114	218	115
rect	218	114	219	115
rect	220	114	221	115
rect	221	114	222	115
rect	229	114	230	115
rect	230	114	231	115
rect	232	114	233	115
rect	233	114	234	115
rect	241	114	242	115
rect	242	114	243	115
rect	244	114	245	115
rect	245	114	246	115
rect	247	114	248	115
rect	248	114	249	115
rect	249	114	250	115
rect	250	114	251	115
rect	251	114	252	115
rect	252	114	253	115
rect	253	114	254	115
rect	254	114	255	115
rect	255	114	256	115
rect	256	114	257	115
rect	257	114	258	115
rect	259	114	260	115
rect	260	114	261	115
rect	262	114	263	115
rect	263	114	264	115
rect	265	114	266	115
rect	266	114	267	115
rect	267	114	268	115
rect	268	114	269	115
rect	269	114	270	115
rect	271	114	272	115
rect	272	114	273	115
rect	274	114	275	115
rect	275	114	276	115
rect	286	114	287	115
rect	287	114	288	115
rect	289	114	290	115
rect	290	114	291	115
rect	292	114	293	115
rect	293	114	294	115
rect	294	114	295	115
rect	295	114	296	115
rect	296	114	297	115
rect	298	114	299	115
rect	299	114	300	115
rect	300	114	301	115
rect	301	114	302	115
rect	302	114	303	115
rect	304	114	305	115
rect	305	114	306	115
rect	306	114	307	115
rect	307	114	308	115
rect	308	114	309	115
rect	309	114	310	115
rect	310	114	311	115
rect	311	114	312	115
rect	313	114	314	115
rect	314	114	315	115
rect	316	114	317	115
rect	317	114	318	115
rect	319	114	320	115
rect	320	114	321	115
rect	321	114	322	115
rect	322	114	323	115
rect	323	114	324	115
rect	324	114	325	115
rect	325	114	326	115
rect	326	114	327	115
rect	328	114	329	115
rect	329	114	330	115
rect	330	114	331	115
rect	331	114	332	115
rect	332	114	333	115
rect	334	114	335	115
rect	335	114	336	115
rect	346	114	347	115
rect	347	114	348	115
rect	349	114	350	115
rect	350	114	351	115
rect	352	114	353	115
rect	353	114	354	115
rect	354	114	355	115
rect	355	114	356	115
rect	356	114	357	115
rect	357	114	358	115
rect	358	114	359	115
rect	359	114	360	115
rect	361	114	362	115
rect	362	114	363	115
rect	363	114	364	115
rect	364	114	365	115
rect	365	114	366	115
rect	366	114	367	115
rect	367	114	368	115
rect	368	114	369	115
rect	90	116	91	117
rect	91	116	92	117
rect	113	116	114	117
rect	114	116	115	117
rect	115	116	116	117
rect	116	116	117	117
rect	117	116	118	117
rect	149	116	150	117
rect	150	116	151	117
rect	151	116	152	117
rect	152	116	153	117
rect	153	116	154	117
rect	154	116	155	117
rect	177	116	178	117
rect	178	116	179	117
rect	179	116	180	117
rect	180	116	181	117
rect	181	116	182	117
rect	182	116	183	117
rect	184	116	185	117
rect	185	116	186	117
rect	186	116	187	117
rect	187	116	188	117
rect	188	116	189	117
rect	190	116	191	117
rect	191	116	192	117
rect	198	116	199	117
rect	199	116	200	117
rect	200	116	201	117
rect	201	116	202	117
rect	202	116	203	117
rect	203	116	204	117
rect	205	116	206	117
rect	206	116	207	117
rect	226	116	227	117
rect	227	116	228	117
rect	228	116	229	117
rect	229	116	230	117
rect	230	116	231	117
rect	232	116	233	117
rect	233	116	234	117
rect	235	116	236	117
rect	236	116	237	117
rect	238	116	239	117
rect	239	116	240	117
rect	240	116	241	117
rect	241	116	242	117
rect	242	116	243	117
rect	244	116	245	117
rect	245	116	246	117
rect	247	116	248	117
rect	248	116	249	117
rect	249	116	250	117
rect	250	116	251	117
rect	251	116	252	117
rect	252	116	253	117
rect	253	116	254	117
rect	254	116	255	117
rect	255	116	256	117
rect	256	116	257	117
rect	257	116	258	117
rect	259	116	260	117
rect	260	116	261	117
rect	262	116	263	117
rect	263	116	264	117
rect	265	116	266	117
rect	266	116	267	117
rect	274	116	275	117
rect	275	116	276	117
rect	277	116	278	117
rect	278	116	279	117
rect	280	116	281	117
rect	281	116	282	117
rect	282	116	283	117
rect	283	116	284	117
rect	284	116	285	117
rect	295	116	296	117
rect	296	116	297	117
rect	298	116	299	117
rect	299	116	300	117
rect	300	116	301	117
rect	301	116	302	117
rect	302	116	303	117
rect	304	116	305	117
rect	305	116	306	117
rect	306	116	307	117
rect	307	116	308	117
rect	308	116	309	117
rect	316	116	317	117
rect	317	116	318	117
rect	319	116	320	117
rect	320	116	321	117
rect	321	116	322	117
rect	322	116	323	117
rect	323	116	324	117
rect	324	116	325	117
rect	325	116	326	117
rect	326	116	327	117
rect	328	116	329	117
rect	329	116	330	117
rect	330	116	331	117
rect	331	116	332	117
rect	332	116	333	117
rect	334	116	335	117
rect	335	116	336	117
rect	337	116	338	117
rect	338	116	339	117
rect	340	116	341	117
rect	341	116	342	117
rect	343	116	344	117
rect	344	116	345	117
rect	345	116	346	117
rect	346	116	347	117
rect	347	116	348	117
rect	349	116	350	117
rect	350	116	351	117
rect	352	116	353	117
rect	353	116	354	117
rect	354	116	355	117
rect	355	116	356	117
rect	356	116	357	117
rect	357	116	358	117
rect	358	116	359	117
rect	359	116	360	117
rect	361	116	362	117
rect	362	116	363	117
rect	41	118	42	119
rect	60	118	61	119
rect	61	118	62	119
rect	62	118	63	119
rect	63	118	64	119
rect	64	118	65	119
rect	65	118	66	119
rect	66	118	67	119
rect	67	118	68	119
rect	69	118	70	119
rect	87	118	88	119
rect	88	118	89	119
rect	110	118	111	119
rect	111	118	112	119
rect	112	118	113	119
rect	113	118	114	119
rect	114	118	115	119
rect	122	118	123	119
rect	123	118	124	119
rect	124	118	125	119
rect	125	118	126	119
rect	126	118	127	119
rect	131	118	132	119
rect	132	118	133	119
rect	133	118	134	119
rect	134	118	135	119
rect	135	118	136	119
rect	140	118	141	119
rect	141	118	142	119
rect	142	118	143	119
rect	143	118	144	119
rect	144	118	145	119
rect	145	118	146	119
rect	146	118	147	119
rect	147	118	148	119
rect	148	118	149	119
rect	149	118	150	119
rect	150	118	151	119
rect	151	118	152	119
rect	171	118	172	119
rect	172	118	173	119
rect	173	118	174	119
rect	175	118	176	119
rect	176	118	177	119
rect	187	118	188	119
rect	188	118	189	119
rect	190	118	191	119
rect	191	118	192	119
rect	193	118	194	119
rect	194	118	195	119
rect	196	118	197	119
rect	197	118	198	119
rect	198	118	199	119
rect	199	118	200	119
rect	200	118	201	119
rect	201	118	202	119
rect	202	118	203	119
rect	203	118	204	119
rect	205	118	206	119
rect	206	118	207	119
rect	208	118	209	119
rect	209	118	210	119
rect	210	118	211	119
rect	211	118	212	119
rect	212	118	213	119
rect	214	118	215	119
rect	215	118	216	119
rect	217	118	218	119
rect	218	118	219	119
rect	220	118	221	119
rect	221	118	222	119
rect	223	118	224	119
rect	224	118	225	119
rect	225	118	226	119
rect	226	118	227	119
rect	227	118	228	119
rect	228	118	229	119
rect	229	118	230	119
rect	230	118	231	119
rect	232	118	233	119
rect	233	118	234	119
rect	235	118	236	119
rect	236	118	237	119
rect	238	118	239	119
rect	239	118	240	119
rect	240	118	241	119
rect	241	118	242	119
rect	242	118	243	119
rect	244	118	245	119
rect	245	118	246	119
rect	247	118	248	119
rect	248	118	249	119
rect	249	118	250	119
rect	250	118	251	119
rect	251	118	252	119
rect	252	118	253	119
rect	253	118	254	119
rect	254	118	255	119
rect	255	118	256	119
rect	256	118	257	119
rect	257	118	258	119
rect	259	118	260	119
rect	260	118	261	119
rect	262	118	263	119
rect	263	118	264	119
rect	265	118	266	119
rect	266	118	267	119
rect	268	118	269	119
rect	269	118	270	119
rect	271	118	272	119
rect	272	118	273	119
rect	273	118	274	119
rect	274	118	275	119
rect	275	118	276	119
rect	277	118	278	119
rect	278	118	279	119
rect	280	118	281	119
rect	281	118	282	119
rect	282	118	283	119
rect	283	118	284	119
rect	284	118	285	119
rect	286	118	287	119
rect	287	118	288	119
rect	289	118	290	119
rect	290	118	291	119
rect	292	118	293	119
rect	293	118	294	119
rect	295	118	296	119
rect	296	118	297	119
rect	298	118	299	119
rect	299	118	300	119
rect	300	118	301	119
rect	301	118	302	119
rect	302	118	303	119
rect	304	118	305	119
rect	305	118	306	119
rect	306	118	307	119
rect	307	118	308	119
rect	308	118	309	119
rect	310	118	311	119
rect	311	118	312	119
rect	313	118	314	119
rect	314	118	315	119
rect	315	118	316	119
rect	316	118	317	119
rect	317	118	318	119
rect	319	118	320	119
rect	320	118	321	119
rect	321	118	322	119
rect	322	118	323	119
rect	323	118	324	119
rect	324	118	325	119
rect	325	118	326	119
rect	326	118	327	119
rect	328	118	329	119
rect	329	118	330	119
rect	330	118	331	119
rect	331	118	332	119
rect	332	118	333	119
rect	334	118	335	119
rect	335	118	336	119
rect	337	118	338	119
rect	338	118	339	119
rect	340	118	341	119
rect	341	118	342	119
rect	343	118	344	119
rect	344	118	345	119
rect	345	118	346	119
rect	346	118	347	119
rect	347	118	348	119
rect	349	118	350	119
rect	350	118	351	119
rect	352	118	353	119
rect	353	118	354	119
rect	354	118	355	119
rect	355	118	356	119
rect	356	118	357	119
rect	38	120	39	121
rect	57	120	58	121
rect	62	120	63	121
rect	63	120	64	121
rect	64	120	65	121
rect	65	120	66	121
rect	66	120	67	121
rect	67	120	68	121
rect	78	120	79	121
rect	79	120	80	121
rect	80	120	81	121
rect	81	120	82	121
rect	82	120	83	121
rect	83	120	84	121
rect	84	120	85	121
rect	85	120	86	121
rect	96	120	97	121
rect	97	120	98	121
rect	98	120	99	121
rect	99	120	100	121
rect	100	120	101	121
rect	101	120	102	121
rect	102	120	103	121
rect	103	120	104	121
rect	104	120	105	121
rect	105	120	106	121
rect	106	120	107	121
rect	107	120	108	121
rect	108	120	109	121
rect	110	120	111	121
rect	111	120	112	121
rect	112	120	113	121
rect	113	120	114	121
rect	114	120	115	121
rect	116	120	117	121
rect	117	120	118	121
rect	119	120	120	121
rect	120	120	121	121
rect	121	120	122	121
rect	122	120	123	121
rect	123	120	124	121
rect	124	120	125	121
rect	125	120	126	121
rect	126	120	127	121
rect	128	120	129	121
rect	129	120	130	121
rect	130	120	131	121
rect	131	120	132	121
rect	132	120	133	121
rect	133	120	134	121
rect	134	120	135	121
rect	135	120	136	121
rect	137	120	138	121
rect	138	120	139	121
rect	139	120	140	121
rect	140	120	141	121
rect	141	120	142	121
rect	142	120	143	121
rect	143	120	144	121
rect	144	120	145	121
rect	145	120	146	121
rect	146	120	147	121
rect	147	120	148	121
rect	148	120	149	121
rect	149	120	150	121
rect	150	120	151	121
rect	151	120	152	121
rect	153	120	154	121
rect	154	120	155	121
rect	156	120	157	121
rect	157	120	158	121
rect	158	120	159	121
rect	159	120	160	121
rect	160	120	161	121
rect	161	120	162	121
rect	162	120	163	121
rect	163	120	164	121
rect	164	120	165	121
rect	165	120	166	121
rect	166	120	167	121
rect	168	120	169	121
rect	169	120	170	121
rect	170	120	171	121
rect	171	120	172	121
rect	172	120	173	121
rect	173	120	174	121
rect	175	120	176	121
rect	176	120	177	121
rect	178	120	179	121
rect	179	120	180	121
rect	180	120	181	121
rect	181	120	182	121
rect	182	120	183	121
rect	184	120	185	121
rect	185	120	186	121
rect	187	120	188	121
rect	188	120	189	121
rect	190	120	191	121
rect	191	120	192	121
rect	193	120	194	121
rect	194	120	195	121
rect	196	120	197	121
rect	197	120	198	121
rect	198	120	199	121
rect	199	120	200	121
rect	200	120	201	121
rect	201	120	202	121
rect	202	120	203	121
rect	203	120	204	121
rect	205	120	206	121
rect	206	120	207	121
rect	208	120	209	121
rect	209	120	210	121
rect	210	120	211	121
rect	211	120	212	121
rect	212	120	213	121
rect	214	120	215	121
rect	215	120	216	121
rect	217	120	218	121
rect	218	120	219	121
rect	220	120	221	121
rect	221	120	222	121
rect	223	120	224	121
rect	224	120	225	121
rect	225	120	226	121
rect	226	120	227	121
rect	227	120	228	121
rect	228	120	229	121
rect	229	120	230	121
rect	230	120	231	121
rect	232	120	233	121
rect	233	120	234	121
rect	235	120	236	121
rect	236	120	237	121
rect	238	120	239	121
rect	239	120	240	121
rect	240	120	241	121
rect	241	120	242	121
rect	242	120	243	121
rect	244	120	245	121
rect	245	120	246	121
rect	247	120	248	121
rect	248	120	249	121
rect	249	120	250	121
rect	250	120	251	121
rect	251	120	252	121
rect	252	120	253	121
rect	253	120	254	121
rect	254	120	255	121
rect	255	120	256	121
rect	256	120	257	121
rect	257	120	258	121
rect	259	120	260	121
rect	260	120	261	121
rect	262	120	263	121
rect	263	120	264	121
rect	265	120	266	121
rect	266	120	267	121
rect	268	120	269	121
rect	269	120	270	121
rect	271	120	272	121
rect	272	120	273	121
rect	273	120	274	121
rect	274	120	275	121
rect	275	120	276	121
rect	277	120	278	121
rect	278	120	279	121
rect	280	120	281	121
rect	281	120	282	121
rect	282	120	283	121
rect	283	120	284	121
rect	284	120	285	121
rect	286	120	287	121
rect	287	120	288	121
rect	289	120	290	121
rect	290	120	291	121
rect	292	120	293	121
rect	293	120	294	121
rect	295	120	296	121
rect	296	120	297	121
rect	298	120	299	121
rect	299	120	300	121
rect	300	120	301	121
rect	301	120	302	121
rect	302	120	303	121
rect	304	120	305	121
rect	305	120	306	121
rect	306	120	307	121
rect	307	120	308	121
rect	308	120	309	121
rect	310	120	311	121
rect	311	120	312	121
rect	313	120	314	121
rect	314	120	315	121
rect	315	120	316	121
rect	316	120	317	121
rect	317	120	318	121
rect	319	120	320	121
rect	320	120	321	121
rect	334	120	335	121
rect	335	120	336	121
rect	337	120	338	121
rect	338	120	339	121
rect	340	120	341	121
rect	341	120	342	121
rect	343	120	344	121
rect	344	120	345	121
rect	345	120	346	121
rect	346	120	347	121
rect	347	120	348	121
rect	349	120	350	121
rect	350	120	351	121
rect	352	120	353	121
rect	353	120	354	121
rect	354	120	355	121
rect	355	120	356	121
rect	356	120	357	121
rect	358	120	359	121
rect	359	120	360	121
rect	361	120	362	121
rect	362	120	363	121
rect	364	120	365	121
rect	365	120	366	121
rect	32	122	33	123
rect	33	122	34	123
rect	35	122	36	123
rect	36	122	37	123
rect	37	122	38	123
rect	38	122	39	123
rect	40	122	41	123
rect	41	122	42	123
rect	43	122	44	123
rect	44	122	45	123
rect	45	122	46	123
rect	46	122	47	123
rect	47	122	48	123
rect	48	122	49	123
rect	49	122	50	123
rect	50	122	51	123
rect	51	122	52	123
rect	52	122	53	123
rect	53	122	54	123
rect	54	122	55	123
rect	55	122	56	123
rect	56	122	57	123
rect	57	122	58	123
rect	59	122	60	123
rect	60	122	61	123
rect	62	122	63	123
rect	63	122	64	123
rect	64	122	65	123
rect	65	122	66	123
rect	66	122	67	123
rect	67	122	68	123
rect	68	122	69	123
rect	69	122	70	123
rect	71	122	72	123
rect	72	122	73	123
rect	73	122	74	123
rect	74	122	75	123
rect	75	122	76	123
rect	76	122	77	123
rect	77	122	78	123
rect	78	122	79	123
rect	79	122	80	123
rect	80	122	81	123
rect	81	122	82	123
rect	82	122	83	123
rect	83	122	84	123
rect	84	122	85	123
rect	85	122	86	123
rect	87	122	88	123
rect	88	122	89	123
rect	90	122	91	123
rect	91	122	92	123
rect	93	122	94	123
rect	94	122	95	123
rect	96	122	97	123
rect	97	122	98	123
rect	98	122	99	123
rect	99	122	100	123
rect	100	122	101	123
rect	101	122	102	123
rect	102	122	103	123
rect	103	122	104	123
rect	104	122	105	123
rect	105	122	106	123
rect	106	122	107	123
rect	107	122	108	123
rect	108	122	109	123
rect	110	122	111	123
rect	111	122	112	123
rect	112	122	113	123
rect	113	122	114	123
rect	114	122	115	123
rect	116	122	117	123
rect	117	122	118	123
rect	119	122	120	123
rect	120	122	121	123
rect	121	122	122	123
rect	122	122	123	123
rect	123	122	124	123
rect	124	122	125	123
rect	125	122	126	123
rect	126	122	127	123
rect	128	122	129	123
rect	129	122	130	123
rect	130	122	131	123
rect	131	122	132	123
rect	132	122	133	123
rect	133	122	134	123
rect	134	122	135	123
rect	135	122	136	123
rect	137	122	138	123
rect	138	122	139	123
rect	139	122	140	123
rect	140	122	141	123
rect	141	122	142	123
rect	142	122	143	123
rect	143	122	144	123
rect	144	122	145	123
rect	145	122	146	123
rect	146	122	147	123
rect	147	122	148	123
rect	148	122	149	123
rect	149	122	150	123
rect	150	122	151	123
rect	151	122	152	123
rect	153	122	154	123
rect	154	122	155	123
rect	156	122	157	123
rect	157	122	158	123
rect	168	122	169	123
rect	169	122	170	123
rect	170	122	171	123
rect	171	122	172	123
rect	172	122	173	123
rect	173	122	174	123
rect	175	122	176	123
rect	176	122	177	123
rect	178	122	179	123
rect	179	122	180	123
rect	180	122	181	123
rect	181	122	182	123
rect	182	122	183	123
rect	184	122	185	123
rect	185	122	186	123
rect	187	122	188	123
rect	188	122	189	123
rect	190	122	191	123
rect	191	122	192	123
rect	193	122	194	123
rect	194	122	195	123
rect	196	122	197	123
rect	197	122	198	123
rect	198	122	199	123
rect	199	122	200	123
rect	200	122	201	123
rect	201	122	202	123
rect	202	122	203	123
rect	203	122	204	123
rect	205	122	206	123
rect	206	122	207	123
rect	208	122	209	123
rect	209	122	210	123
rect	226	122	227	123
rect	227	122	228	123
rect	228	122	229	123
rect	229	122	230	123
rect	230	122	231	123
rect	238	122	239	123
rect	239	122	240	123
rect	240	122	241	123
rect	241	122	242	123
rect	242	122	243	123
rect	244	122	245	123
rect	245	122	246	123
rect	247	122	248	123
rect	248	122	249	123
rect	249	122	250	123
rect	250	122	251	123
rect	251	122	252	123
rect	252	122	253	123
rect	253	122	254	123
rect	254	122	255	123
rect	255	122	256	123
rect	256	122	257	123
rect	257	122	258	123
rect	259	122	260	123
rect	260	122	261	123
rect	262	122	263	123
rect	263	122	264	123
rect	265	122	266	123
rect	266	122	267	123
rect	268	122	269	123
rect	269	122	270	123
rect	271	122	272	123
rect	272	122	273	123
rect	273	122	274	123
rect	274	122	275	123
rect	275	122	276	123
rect	277	122	278	123
rect	278	122	279	123
rect	280	122	281	123
rect	281	122	282	123
rect	282	122	283	123
rect	283	122	284	123
rect	284	122	285	123
rect	286	122	287	123
rect	287	122	288	123
rect	289	122	290	123
rect	290	122	291	123
rect	292	122	293	123
rect	293	122	294	123
rect	295	122	296	123
rect	296	122	297	123
rect	298	122	299	123
rect	299	122	300	123
rect	300	122	301	123
rect	301	122	302	123
rect	302	122	303	123
rect	304	122	305	123
rect	305	122	306	123
rect	306	122	307	123
rect	307	122	308	123
rect	308	122	309	123
rect	310	122	311	123
rect	311	122	312	123
rect	313	122	314	123
rect	314	122	315	123
rect	319	122	320	123
rect	320	122	321	123
rect	322	122	323	123
rect	323	122	324	123
rect	324	122	325	123
rect	325	122	326	123
rect	326	122	327	123
rect	328	122	329	123
rect	329	122	330	123
rect	330	122	331	123
rect	331	122	332	123
rect	332	122	333	123
rect	361	122	362	123
rect	362	122	363	123
rect	364	122	365	123
rect	365	122	366	123
rect	367	122	368	123
rect	368	122	369	123
rect	19	124	20	125
rect	20	124	21	125
rect	29	124	30	125
rect	35	124	36	125
rect	36	124	37	125
rect	37	124	38	125
rect	38	124	39	125
rect	40	124	41	125
rect	41	124	42	125
rect	43	124	44	125
rect	44	124	45	125
rect	45	124	46	125
rect	46	124	47	125
rect	47	124	48	125
rect	48	124	49	125
rect	49	124	50	125
rect	50	124	51	125
rect	51	124	52	125
rect	52	124	53	125
rect	53	124	54	125
rect	54	124	55	125
rect	55	124	56	125
rect	56	124	57	125
rect	57	124	58	125
rect	59	124	60	125
rect	60	124	61	125
rect	62	124	63	125
rect	63	124	64	125
rect	64	124	65	125
rect	65	124	66	125
rect	66	124	67	125
rect	67	124	68	125
rect	68	124	69	125
rect	69	124	70	125
rect	71	124	72	125
rect	72	124	73	125
rect	73	124	74	125
rect	74	124	75	125
rect	75	124	76	125
rect	76	124	77	125
rect	77	124	78	125
rect	78	124	79	125
rect	79	124	80	125
rect	80	124	81	125
rect	81	124	82	125
rect	82	124	83	125
rect	83	124	84	125
rect	84	124	85	125
rect	85	124	86	125
rect	87	124	88	125
rect	88	124	89	125
rect	90	124	91	125
rect	91	124	92	125
rect	93	124	94	125
rect	94	124	95	125
rect	96	124	97	125
rect	97	124	98	125
rect	98	124	99	125
rect	99	124	100	125
rect	100	124	101	125
rect	101	124	102	125
rect	102	124	103	125
rect	103	124	104	125
rect	104	124	105	125
rect	105	124	106	125
rect	106	124	107	125
rect	107	124	108	125
rect	108	124	109	125
rect	110	124	111	125
rect	111	124	112	125
rect	112	124	113	125
rect	113	124	114	125
rect	114	124	115	125
rect	116	124	117	125
rect	117	124	118	125
rect	119	124	120	125
rect	120	124	121	125
rect	121	124	122	125
rect	122	124	123	125
rect	123	124	124	125
rect	124	124	125	125
rect	125	124	126	125
rect	126	124	127	125
rect	128	124	129	125
rect	129	124	130	125
rect	130	124	131	125
rect	131	124	132	125
rect	132	124	133	125
rect	133	124	134	125
rect	134	124	135	125
rect	135	124	136	125
rect	137	124	138	125
rect	138	124	139	125
rect	139	124	140	125
rect	140	124	141	125
rect	141	124	142	125
rect	142	124	143	125
rect	143	124	144	125
rect	144	124	145	125
rect	145	124	146	125
rect	146	124	147	125
rect	147	124	148	125
rect	148	124	149	125
rect	149	124	150	125
rect	150	124	151	125
rect	151	124	152	125
rect	153	124	154	125
rect	154	124	155	125
rect	156	124	157	125
rect	157	124	158	125
rect	159	124	160	125
rect	160	124	161	125
rect	161	124	162	125
rect	162	124	163	125
rect	163	124	164	125
rect	164	124	165	125
rect	165	124	166	125
rect	166	124	167	125
rect	167	124	168	125
rect	168	124	169	125
rect	169	124	170	125
rect	170	124	171	125
rect	171	124	172	125
rect	172	124	173	125
rect	173	124	174	125
rect	175	124	176	125
rect	176	124	177	125
rect	178	124	179	125
rect	179	124	180	125
rect	180	124	181	125
rect	181	124	182	125
rect	182	124	183	125
rect	184	124	185	125
rect	185	124	186	125
rect	187	124	188	125
rect	188	124	189	125
rect	190	124	191	125
rect	191	124	192	125
rect	193	124	194	125
rect	194	124	195	125
rect	196	124	197	125
rect	197	124	198	125
rect	198	124	199	125
rect	199	124	200	125
rect	200	124	201	125
rect	201	124	202	125
rect	202	124	203	125
rect	203	124	204	125
rect	205	124	206	125
rect	206	124	207	125
rect	208	124	209	125
rect	209	124	210	125
rect	211	124	212	125
rect	212	124	213	125
rect	214	124	215	125
rect	215	124	216	125
rect	217	124	218	125
rect	218	124	219	125
rect	220	124	221	125
rect	221	124	222	125
rect	223	124	224	125
rect	224	124	225	125
rect	226	124	227	125
rect	227	124	228	125
rect	228	124	229	125
rect	229	124	230	125
rect	230	124	231	125
rect	231	124	232	125
rect	232	124	233	125
rect	233	124	234	125
rect	235	124	236	125
rect	236	124	237	125
rect	237	124	238	125
rect	238	124	239	125
rect	239	124	240	125
rect	240	124	241	125
rect	241	124	242	125
rect	242	124	243	125
rect	244	124	245	125
rect	245	124	246	125
rect	247	124	248	125
rect	248	124	249	125
rect	271	124	272	125
rect	272	124	273	125
rect	273	124	274	125
rect	274	124	275	125
rect	275	124	276	125
rect	277	124	278	125
rect	278	124	279	125
rect	280	124	281	125
rect	281	124	282	125
rect	292	124	293	125
rect	293	124	294	125
rect	295	124	296	125
rect	296	124	297	125
rect	298	124	299	125
rect	299	124	300	125
rect	300	124	301	125
rect	301	124	302	125
rect	302	124	303	125
rect	304	124	305	125
rect	305	124	306	125
rect	306	124	307	125
rect	307	124	308	125
rect	308	124	309	125
rect	310	124	311	125
rect	311	124	312	125
rect	313	124	314	125
rect	314	124	315	125
rect	316	124	317	125
rect	317	124	318	125
rect	355	124	356	125
rect	356	124	357	125
rect	358	124	359	125
rect	359	124	360	125
rect	397	124	398	125
rect	398	124	399	125
rect	399	124	400	125
rect	400	124	401	125
rect	401	124	402	125
rect	403	124	404	125
rect	404	124	405	125
rect	405	124	406	125
rect	406	124	407	125
rect	407	124	408	125
rect	408	124	409	125
rect	409	124	410	125
rect	410	124	411	125
rect	411	124	412	125
rect	412	124	413	125
rect	413	124	414	125
rect	414	124	415	125
rect	415	124	416	125
rect	12	126	13	127
rect	13	126	14	127
rect	14	126	15	127
rect	15	126	16	127
rect	16	126	17	127
rect	17	126	18	127
rect	19	126	20	127
rect	20	126	21	127
rect	22	126	23	127
rect	23	126	24	127
rect	24	126	25	127
rect	25	126	26	127
rect	26	126	27	127
rect	27	126	28	127
rect	28	126	29	127
rect	29	126	30	127
rect	31	126	32	127
rect	32	126	33	127
rect	33	126	34	127
rect	34	126	35	127
rect	35	126	36	127
rect	36	126	37	127
rect	37	126	38	127
rect	38	126	39	127
rect	40	126	41	127
rect	41	126	42	127
rect	43	126	44	127
rect	44	126	45	127
rect	45	126	46	127
rect	46	126	47	127
rect	47	126	48	127
rect	48	126	49	127
rect	49	126	50	127
rect	50	126	51	127
rect	51	126	52	127
rect	52	126	53	127
rect	53	126	54	127
rect	54	126	55	127
rect	55	126	56	127
rect	56	126	57	127
rect	57	126	58	127
rect	59	126	60	127
rect	60	126	61	127
rect	62	126	63	127
rect	63	126	64	127
rect	64	126	65	127
rect	65	126	66	127
rect	66	126	67	127
rect	67	126	68	127
rect	68	126	69	127
rect	69	126	70	127
rect	71	126	72	127
rect	72	126	73	127
rect	73	126	74	127
rect	74	126	75	127
rect	75	126	76	127
rect	76	126	77	127
rect	77	126	78	127
rect	78	126	79	127
rect	79	126	80	127
rect	80	126	81	127
rect	81	126	82	127
rect	82	126	83	127
rect	83	126	84	127
rect	84	126	85	127
rect	85	126	86	127
rect	87	126	88	127
rect	88	126	89	127
rect	90	126	91	127
rect	91	126	92	127
rect	93	126	94	127
rect	94	126	95	127
rect	96	126	97	127
rect	97	126	98	127
rect	98	126	99	127
rect	99	126	100	127
rect	100	126	101	127
rect	101	126	102	127
rect	102	126	103	127
rect	103	126	104	127
rect	104	126	105	127
rect	105	126	106	127
rect	106	126	107	127
rect	107	126	108	127
rect	108	126	109	127
rect	110	126	111	127
rect	111	126	112	127
rect	112	126	113	127
rect	113	126	114	127
rect	114	126	115	127
rect	116	126	117	127
rect	117	126	118	127
rect	119	126	120	127
rect	120	126	121	127
rect	121	126	122	127
rect	122	126	123	127
rect	123	126	124	127
rect	124	126	125	127
rect	125	126	126	127
rect	126	126	127	127
rect	128	126	129	127
rect	129	126	130	127
rect	130	126	131	127
rect	131	126	132	127
rect	132	126	133	127
rect	133	126	134	127
rect	134	126	135	127
rect	135	126	136	127
rect	137	126	138	127
rect	138	126	139	127
rect	139	126	140	127
rect	140	126	141	127
rect	141	126	142	127
rect	142	126	143	127
rect	143	126	144	127
rect	144	126	145	127
rect	145	126	146	127
rect	146	126	147	127
rect	147	126	148	127
rect	148	126	149	127
rect	149	126	150	127
rect	150	126	151	127
rect	151	126	152	127
rect	153	126	154	127
rect	154	126	155	127
rect	156	126	157	127
rect	157	126	158	127
rect	159	126	160	127
rect	160	126	161	127
rect	161	126	162	127
rect	162	126	163	127
rect	163	126	164	127
rect	164	126	165	127
rect	165	126	166	127
rect	166	126	167	127
rect	167	126	168	127
rect	168	126	169	127
rect	169	126	170	127
rect	170	126	171	127
rect	171	126	172	127
rect	172	126	173	127
rect	173	126	174	127
rect	175	126	176	127
rect	176	126	177	127
rect	178	126	179	127
rect	179	126	180	127
rect	180	126	181	127
rect	181	126	182	127
rect	182	126	183	127
rect	184	126	185	127
rect	185	126	186	127
rect	187	126	188	127
rect	188	126	189	127
rect	190	126	191	127
rect	191	126	192	127
rect	193	126	194	127
rect	194	126	195	127
rect	196	126	197	127
rect	197	126	198	127
rect	198	126	199	127
rect	199	126	200	127
rect	200	126	201	127
rect	201	126	202	127
rect	202	126	203	127
rect	203	126	204	127
rect	205	126	206	127
rect	206	126	207	127
rect	208	126	209	127
rect	209	126	210	127
rect	211	126	212	127
rect	212	126	213	127
rect	214	126	215	127
rect	215	126	216	127
rect	217	126	218	127
rect	218	126	219	127
rect	220	126	221	127
rect	221	126	222	127
rect	223	126	224	127
rect	224	126	225	127
rect	226	126	227	127
rect	227	126	228	127
rect	228	126	229	127
rect	229	126	230	127
rect	230	126	231	127
rect	231	126	232	127
rect	232	126	233	127
rect	233	126	234	127
rect	235	126	236	127
rect	236	126	237	127
rect	237	126	238	127
rect	238	126	239	127
rect	239	126	240	127
rect	240	126	241	127
rect	241	126	242	127
rect	242	126	243	127
rect	244	126	245	127
rect	245	126	246	127
rect	247	126	248	127
rect	248	126	249	127
rect	250	126	251	127
rect	251	126	252	127
rect	259	126	260	127
rect	260	126	261	127
rect	262	126	263	127
rect	263	126	264	127
rect	265	126	266	127
rect	266	126	267	127
rect	268	126	269	127
rect	269	126	270	127
rect	270	126	271	127
rect	271	126	272	127
rect	272	126	273	127
rect	289	126	290	127
rect	290	126	291	127
rect	291	126	292	127
rect	292	126	293	127
rect	293	126	294	127
rect	295	126	296	127
rect	296	126	297	127
rect	298	126	299	127
rect	299	126	300	127
rect	328	126	329	127
rect	329	126	330	127
rect	349	126	350	127
rect	350	126	351	127
rect	352	126	353	127
rect	353	126	354	127
rect	355	126	356	127
rect	356	126	357	127
rect	358	126	359	127
rect	359	126	360	127
rect	361	126	362	127
rect	362	126	363	127
rect	364	126	365	127
rect	365	126	366	127
rect	367	126	368	127
rect	368	126	369	127
rect	370	126	371	127
rect	371	126	372	127
rect	373	126	374	127
rect	374	126	375	127
rect	375	126	376	127
rect	376	126	377	127
rect	377	126	378	127
rect	379	126	380	127
rect	380	126	381	127
rect	381	126	382	127
rect	382	126	383	127
rect	383	126	384	127
rect	384	126	385	127
rect	385	126	386	127
rect	386	126	387	127
rect	388	126	389	127
rect	389	126	390	127
rect	390	126	391	127
rect	391	126	392	127
rect	392	126	393	127
rect	393	126	394	127
rect	394	126	395	127
rect	395	126	396	127
rect	217	135	218	136
rect	218	135	219	136
rect	220	135	221	136
rect	221	135	222	136
rect	223	135	224	136
rect	224	135	225	136
rect	226	135	227	136
rect	227	135	228	136
rect	229	135	230	136
rect	230	135	231	136
rect	202	137	203	138
rect	203	137	204	138
rect	205	137	206	138
rect	206	137	207	138
rect	208	137	209	138
rect	209	137	210	138
rect	217	137	218	138
rect	218	137	219	138
rect	220	137	221	138
rect	221	137	222	138
rect	223	137	224	138
rect	224	137	225	138
rect	238	137	239	138
rect	239	137	240	138
rect	240	137	241	138
rect	241	137	242	138
rect	242	137	243	138
rect	244	137	245	138
rect	245	137	246	138
rect	247	137	248	138
rect	248	137	249	138
rect	250	137	251	138
rect	251	137	252	138
rect	253	137	254	138
rect	254	137	255	138
rect	255	137	256	138
rect	256	137	257	138
rect	257	137	258	138
rect	258	137	259	138
rect	259	137	260	138
rect	260	137	261	138
rect	307	137	308	138
rect	308	137	309	138
rect	309	137	310	138
rect	310	137	311	138
rect	311	137	312	138
rect	313	137	314	138
rect	314	137	315	138
rect	150	139	151	140
rect	151	139	152	140
rect	153	139	154	140
rect	154	139	155	140
rect	156	139	157	140
rect	157	139	158	140
rect	159	139	160	140
rect	160	139	161	140
rect	161	139	162	140
rect	162	139	163	140
rect	163	139	164	140
rect	164	139	165	140
rect	165	139	166	140
rect	166	139	167	140
rect	167	139	168	140
rect	168	139	169	140
rect	169	139	170	140
rect	170	139	171	140
rect	171	139	172	140
rect	172	139	173	140
rect	173	139	174	140
rect	175	139	176	140
rect	176	139	177	140
rect	178	139	179	140
rect	179	139	180	140
rect	180	139	181	140
rect	181	139	182	140
rect	182	139	183	140
rect	183	139	184	140
rect	184	139	185	140
rect	185	139	186	140
rect	187	139	188	140
rect	188	139	189	140
rect	190	139	191	140
rect	191	139	192	140
rect	193	139	194	140
rect	194	139	195	140
rect	196	139	197	140
rect	197	139	198	140
rect	198	139	199	140
rect	199	139	200	140
rect	200	139	201	140
rect	202	139	203	140
rect	203	139	204	140
rect	205	139	206	140
rect	206	139	207	140
rect	208	139	209	140
rect	209	139	210	140
rect	210	139	211	140
rect	211	139	212	140
rect	212	139	213	140
rect	214	139	215	140
rect	215	139	216	140
rect	217	139	218	140
rect	218	139	219	140
rect	220	139	221	140
rect	221	139	222	140
rect	223	139	224	140
rect	224	139	225	140
rect	225	139	226	140
rect	226	139	227	140
rect	227	139	228	140
rect	229	139	230	140
rect	230	139	231	140
rect	232	139	233	140
rect	233	139	234	140
rect	235	139	236	140
rect	236	139	237	140
rect	237	139	238	140
rect	238	139	239	140
rect	239	139	240	140
rect	240	139	241	140
rect	241	139	242	140
rect	242	139	243	140
rect	244	139	245	140
rect	245	139	246	140
rect	247	139	248	140
rect	248	139	249	140
rect	250	139	251	140
rect	251	139	252	140
rect	253	139	254	140
rect	254	139	255	140
rect	255	139	256	140
rect	256	139	257	140
rect	257	139	258	140
rect	258	139	259	140
rect	259	139	260	140
rect	260	139	261	140
rect	261	139	262	140
rect	262	139	263	140
rect	263	139	264	140
rect	265	139	266	140
rect	266	139	267	140
rect	277	139	278	140
rect	278	139	279	140
rect	280	139	281	140
rect	281	139	282	140
rect	283	139	284	140
rect	284	139	285	140
rect	286	139	287	140
rect	287	139	288	140
rect	298	139	299	140
rect	299	139	300	140
rect	301	139	302	140
rect	302	139	303	140
rect	304	139	305	140
rect	305	139	306	140
rect	307	139	308	140
rect	308	139	309	140
rect	309	139	310	140
rect	310	139	311	140
rect	311	139	312	140
rect	313	139	314	140
rect	314	139	315	140
rect	184	141	185	142
rect	185	141	186	142
rect	187	141	188	142
rect	188	141	189	142
rect	190	141	191	142
rect	191	141	192	142
rect	193	141	194	142
rect	194	141	195	142
rect	196	141	197	142
rect	197	141	198	142
rect	198	141	199	142
rect	199	141	200	142
rect	200	141	201	142
rect	202	141	203	142
rect	203	141	204	142
rect	205	141	206	142
rect	206	141	207	142
rect	226	141	227	142
rect	227	141	228	142
rect	235	141	236	142
rect	236	141	237	142
rect	237	141	238	142
rect	238	141	239	142
rect	239	141	240	142
rect	240	141	241	142
rect	241	141	242	142
rect	242	141	243	142
rect	244	141	245	142
rect	245	141	246	142
rect	247	141	248	142
rect	248	141	249	142
rect	250	141	251	142
rect	251	141	252	142
rect	253	141	254	142
rect	254	141	255	142
rect	268	141	269	142
rect	269	141	270	142
rect	270	141	271	142
rect	271	141	272	142
rect	272	141	273	142
rect	277	141	278	142
rect	278	141	279	142
rect	292	141	293	142
rect	293	141	294	142
rect	295	141	296	142
rect	296	141	297	142
rect	297	141	298	142
rect	298	141	299	142
rect	299	141	300	142
rect	319	141	320	142
rect	320	141	321	142
rect	322	141	323	142
rect	323	141	324	142
rect	325	141	326	142
rect	326	141	327	142
rect	190	143	191	144
rect	191	143	192	144
rect	193	143	194	144
rect	194	143	195	144
rect	196	143	197	144
rect	197	143	198	144
rect	198	143	199	144
rect	199	143	200	144
rect	200	143	201	144
rect	202	143	203	144
rect	203	143	204	144
rect	205	143	206	144
rect	206	143	207	144
rect	223	143	224	144
rect	224	143	225	144
rect	226	143	227	144
rect	227	143	228	144
rect	228	143	229	144
rect	229	143	230	144
rect	230	143	231	144
rect	232	143	233	144
rect	233	143	234	144
rect	244	143	245	144
rect	245	143	246	144
rect	247	143	248	144
rect	248	143	249	144
rect	250	143	251	144
rect	251	143	252	144
rect	253	143	254	144
rect	254	143	255	144
rect	256	143	257	144
rect	257	143	258	144
rect	258	143	259	144
rect	259	143	260	144
rect	260	143	261	144
rect	265	143	266	144
rect	266	143	267	144
rect	268	143	269	144
rect	269	143	270	144
rect	270	143	271	144
rect	271	143	272	144
rect	272	143	273	144
rect	273	143	274	144
rect	274	143	275	144
rect	275	143	276	144
rect	277	143	278	144
rect	278	143	279	144
rect	286	143	287	144
rect	287	143	288	144
rect	289	143	290	144
rect	290	143	291	144
rect	292	143	293	144
rect	293	143	294	144
rect	295	143	296	144
rect	296	143	297	144
rect	313	143	314	144
rect	314	143	315	144
rect	316	143	317	144
rect	317	143	318	144
rect	318	143	319	144
rect	319	143	320	144
rect	320	143	321	144
rect	322	143	323	144
rect	323	143	324	144
rect	370	143	371	144
rect	371	143	372	144
rect	372	143	373	144
rect	373	143	374	144
rect	374	143	375	144
rect	376	143	377	144
rect	377	143	378	144
rect	379	143	380	144
rect	380	143	381	144
rect	381	143	382	144
rect	93	145	94	146
rect	94	145	95	146
rect	95	145	96	146
rect	96	145	97	146
rect	97	145	98	146
rect	159	145	160	146
rect	160	145	161	146
rect	161	145	162	146
rect	162	145	163	146
rect	163	145	164	146
rect	164	145	165	146
rect	165	145	166	146
rect	166	145	167	146
rect	181	145	182	146
rect	182	145	183	146
rect	184	145	185	146
rect	185	145	186	146
rect	187	145	188	146
rect	188	145	189	146
rect	189	145	190	146
rect	190	145	191	146
rect	191	145	192	146
rect	193	145	194	146
rect	194	145	195	146
rect	196	145	197	146
rect	197	145	198	146
rect	198	145	199	146
rect	199	145	200	146
rect	200	145	201	146
rect	202	145	203	146
rect	203	145	204	146
rect	205	145	206	146
rect	206	145	207	146
rect	208	145	209	146
rect	209	145	210	146
rect	210	145	211	146
rect	211	145	212	146
rect	212	145	213	146
rect	214	145	215	146
rect	215	145	216	146
rect	217	145	218	146
rect	218	145	219	146
rect	220	145	221	146
rect	221	145	222	146
rect	222	145	223	146
rect	223	145	224	146
rect	224	145	225	146
rect	226	145	227	146
rect	227	145	228	146
rect	228	145	229	146
rect	229	145	230	146
rect	230	145	231	146
rect	232	145	233	146
rect	233	145	234	146
rect	235	145	236	146
rect	236	145	237	146
rect	237	145	238	146
rect	238	145	239	146
rect	239	145	240	146
rect	240	145	241	146
rect	241	145	242	146
rect	242	145	243	146
rect	243	145	244	146
rect	244	145	245	146
rect	245	145	246	146
rect	247	145	248	146
rect	248	145	249	146
rect	250	145	251	146
rect	251	145	252	146
rect	253	145	254	146
rect	254	145	255	146
rect	256	145	257	146
rect	257	145	258	146
rect	258	145	259	146
rect	259	145	260	146
rect	260	145	261	146
rect	262	145	263	146
rect	263	145	264	146
rect	264	145	265	146
rect	265	145	266	146
rect	266	145	267	146
rect	268	145	269	146
rect	269	145	270	146
rect	270	145	271	146
rect	271	145	272	146
rect	272	145	273	146
rect	273	145	274	146
rect	274	145	275	146
rect	275	145	276	146
rect	277	145	278	146
rect	278	145	279	146
rect	280	145	281	146
rect	281	145	282	146
rect	283	145	284	146
rect	284	145	285	146
rect	285	145	286	146
rect	286	145	287	146
rect	287	145	288	146
rect	289	145	290	146
rect	290	145	291	146
rect	292	145	293	146
rect	293	145	294	146
rect	295	145	296	146
rect	296	145	297	146
rect	298	145	299	146
rect	299	145	300	146
rect	300	145	301	146
rect	301	145	302	146
rect	302	145	303	146
rect	304	145	305	146
rect	305	145	306	146
rect	307	145	308	146
rect	308	145	309	146
rect	309	145	310	146
rect	310	145	311	146
rect	311	145	312	146
rect	312	145	313	146
rect	313	145	314	146
rect	314	145	315	146
rect	316	145	317	146
rect	317	145	318	146
rect	318	145	319	146
rect	319	145	320	146
rect	320	145	321	146
rect	322	145	323	146
rect	323	145	324	146
rect	324	145	325	146
rect	325	145	326	146
rect	326	145	327	146
rect	328	145	329	146
rect	329	145	330	146
rect	331	145	332	146
rect	332	145	333	146
rect	334	145	335	146
rect	335	145	336	146
rect	337	145	338	146
rect	338	145	339	146
rect	340	145	341	146
rect	341	145	342	146
rect	343	145	344	146
rect	344	145	345	146
rect	345	145	346	146
rect	346	145	347	146
rect	347	145	348	146
rect	348	145	349	146
rect	349	145	350	146
rect	350	145	351	146
rect	351	145	352	146
rect	353	145	354	146
rect	355	145	356	146
rect	356	145	357	146
rect	358	145	359	146
rect	359	145	360	146
rect	360	145	361	146
rect	361	145	362	146
rect	362	145	363	146
rect	364	145	365	146
rect	365	145	366	146
rect	367	145	368	146
rect	368	145	369	146
rect	369	145	370	146
rect	370	145	371	146
rect	371	145	372	146
rect	372	145	373	146
rect	373	145	374	146
rect	374	145	375	146
rect	376	145	377	146
rect	377	145	378	146
rect	379	145	380	146
rect	380	145	381	146
rect	381	145	382	146
rect	383	145	384	146
rect	384	145	385	146
rect	385	145	386	146
rect	386	145	387	146
rect	388	145	389	146
rect	389	145	390	146
rect	390	145	391	146
rect	391	145	392	146
rect	392	145	393	146
rect	393	145	394	146
rect	394	145	395	146
rect	395	145	396	146
rect	397	145	398	146
rect	398	145	399	146
rect	399	145	400	146
rect	400	145	401	146
rect	401	145	402	146
rect	403	145	404	146
rect	404	145	405	146
rect	405	145	406	146
rect	406	145	407	146
rect	407	145	408	146
rect	408	145	409	146
rect	409	145	410	146
rect	90	147	91	148
rect	91	147	92	148
rect	92	147	93	148
rect	93	147	94	148
rect	94	147	95	148
rect	137	147	138	148
rect	138	147	139	148
rect	139	147	140	148
rect	159	147	160	148
rect	160	147	161	148
rect	161	147	162	148
rect	162	147	163	148
rect	163	147	164	148
rect	164	147	165	148
rect	165	147	166	148
rect	166	147	167	148
rect	168	147	169	148
rect	169	147	170	148
rect	170	147	171	148
rect	171	147	172	148
rect	172	147	173	148
rect	173	147	174	148
rect	175	147	176	148
rect	176	147	177	148
rect	178	147	179	148
rect	179	147	180	148
rect	181	147	182	148
rect	182	147	183	148
rect	184	147	185	148
rect	185	147	186	148
rect	187	147	188	148
rect	188	147	189	148
rect	189	147	190	148
rect	190	147	191	148
rect	191	147	192	148
rect	193	147	194	148
rect	194	147	195	148
rect	196	147	197	148
rect	197	147	198	148
rect	198	147	199	148
rect	199	147	200	148
rect	200	147	201	148
rect	202	147	203	148
rect	203	147	204	148
rect	205	147	206	148
rect	206	147	207	148
rect	208	147	209	148
rect	209	147	210	148
rect	210	147	211	148
rect	211	147	212	148
rect	212	147	213	148
rect	214	147	215	148
rect	215	147	216	148
rect	217	147	218	148
rect	218	147	219	148
rect	220	147	221	148
rect	221	147	222	148
rect	222	147	223	148
rect	223	147	224	148
rect	224	147	225	148
rect	226	147	227	148
rect	227	147	228	148
rect	228	147	229	148
rect	229	147	230	148
rect	230	147	231	148
rect	232	147	233	148
rect	233	147	234	148
rect	235	147	236	148
rect	236	147	237	148
rect	237	147	238	148
rect	238	147	239	148
rect	239	147	240	148
rect	240	147	241	148
rect	241	147	242	148
rect	242	147	243	148
rect	243	147	244	148
rect	244	147	245	148
rect	245	147	246	148
rect	247	147	248	148
rect	248	147	249	148
rect	250	147	251	148
rect	251	147	252	148
rect	253	147	254	148
rect	254	147	255	148
rect	256	147	257	148
rect	257	147	258	148
rect	258	147	259	148
rect	259	147	260	148
rect	260	147	261	148
rect	262	147	263	148
rect	263	147	264	148
rect	264	147	265	148
rect	265	147	266	148
rect	266	147	267	148
rect	268	147	269	148
rect	269	147	270	148
rect	270	147	271	148
rect	271	147	272	148
rect	272	147	273	148
rect	273	147	274	148
rect	274	147	275	148
rect	275	147	276	148
rect	277	147	278	148
rect	278	147	279	148
rect	280	147	281	148
rect	281	147	282	148
rect	283	147	284	148
rect	284	147	285	148
rect	285	147	286	148
rect	286	147	287	148
rect	287	147	288	148
rect	289	147	290	148
rect	290	147	291	148
rect	292	147	293	148
rect	293	147	294	148
rect	295	147	296	148
rect	296	147	297	148
rect	298	147	299	148
rect	299	147	300	148
rect	313	147	314	148
rect	314	147	315	148
rect	316	147	317	148
rect	317	147	318	148
rect	318	147	319	148
rect	319	147	320	148
rect	320	147	321	148
rect	322	147	323	148
rect	323	147	324	148
rect	324	147	325	148
rect	325	147	326	148
rect	326	147	327	148
rect	328	147	329	148
rect	329	147	330	148
rect	347	147	348	148
rect	348	147	349	148
rect	349	147	350	148
rect	350	147	351	148
rect	351	147	352	148
rect	353	147	354	148
rect	355	147	356	148
rect	356	147	357	148
rect	367	147	368	148
rect	368	147	369	148
rect	369	147	370	148
rect	370	147	371	148
rect	371	147	372	148
rect	372	147	373	148
rect	43	149	44	150
rect	44	149	45	150
rect	45	149	46	150
rect	46	149	47	150
rect	87	149	88	150
rect	88	149	89	150
rect	89	149	90	150
rect	90	149	91	150
rect	91	149	92	150
rect	92	149	93	150
rect	93	149	94	150
rect	94	149	95	150
rect	96	149	97	150
rect	97	149	98	150
rect	99	149	100	150
rect	100	149	101	150
rect	101	149	102	150
rect	102	149	103	150
rect	103	149	104	150
rect	104	149	105	150
rect	105	149	106	150
rect	106	149	107	150
rect	128	149	129	150
rect	129	149	130	150
rect	131	149	132	150
rect	132	149	133	150
rect	133	149	134	150
rect	134	149	135	150
rect	135	149	136	150
rect	136	149	137	150
rect	156	149	157	150
rect	157	149	158	150
rect	159	149	160	150
rect	160	149	161	150
rect	161	149	162	150
rect	162	149	163	150
rect	163	149	164	150
rect	178	149	179	150
rect	179	149	180	150
rect	181	149	182	150
rect	182	149	183	150
rect	184	149	185	150
rect	185	149	186	150
rect	187	149	188	150
rect	188	149	189	150
rect	193	149	194	150
rect	194	149	195	150
rect	196	149	197	150
rect	197	149	198	150
rect	198	149	199	150
rect	199	149	200	150
rect	200	149	201	150
rect	202	149	203	150
rect	203	149	204	150
rect	205	149	206	150
rect	206	149	207	150
rect	208	149	209	150
rect	209	149	210	150
rect	214	149	215	150
rect	215	149	216	150
rect	217	149	218	150
rect	218	149	219	150
rect	220	149	221	150
rect	221	149	222	150
rect	222	149	223	150
rect	223	149	224	150
rect	224	149	225	150
rect	226	149	227	150
rect	227	149	228	150
rect	238	149	239	150
rect	239	149	240	150
rect	240	149	241	150
rect	241	149	242	150
rect	242	149	243	150
rect	243	149	244	150
rect	244	149	245	150
rect	245	149	246	150
rect	253	149	254	150
rect	254	149	255	150
rect	256	149	257	150
rect	257	149	258	150
rect	258	149	259	150
rect	259	149	260	150
rect	260	149	261	150
rect	262	149	263	150
rect	263	149	264	150
rect	274	149	275	150
rect	275	149	276	150
rect	277	149	278	150
rect	278	149	279	150
rect	280	149	281	150
rect	281	149	282	150
rect	283	149	284	150
rect	284	149	285	150
rect	285	149	286	150
rect	286	149	287	150
rect	287	149	288	150
rect	289	149	290	150
rect	290	149	291	150
rect	292	149	293	150
rect	293	149	294	150
rect	310	149	311	150
rect	311	149	312	150
rect	313	149	314	150
rect	314	149	315	150
rect	316	149	317	150
rect	317	149	318	150
rect	318	149	319	150
rect	319	149	320	150
rect	320	149	321	150
rect	322	149	323	150
rect	323	149	324	150
rect	324	149	325	150
rect	325	149	326	150
rect	326	149	327	150
rect	328	149	329	150
rect	329	149	330	150
rect	330	149	331	150
rect	331	149	332	150
rect	332	149	333	150
rect	343	149	344	150
rect	344	149	345	150
rect	345	149	346	150
rect	347	149	348	150
rect	348	149	349	150
rect	355	149	356	150
rect	356	149	357	150
rect	357	149	358	150
rect	358	149	359	150
rect	359	149	360	150
rect	360	149	361	150
rect	361	149	362	150
rect	362	149	363	150
rect	364	149	365	150
rect	365	149	366	150
rect	366	149	367	150
rect	367	149	368	150
rect	368	149	369	150
rect	369	149	370	150
rect	37	151	38	152
rect	38	151	39	152
rect	40	151	41	152
rect	41	151	42	152
rect	42	151	43	152
rect	43	151	44	152
rect	44	151	45	152
rect	45	151	46	152
rect	46	151	47	152
rect	48	151	49	152
rect	49	151	50	152
rect	50	151	51	152
rect	51	151	52	152
rect	52	151	53	152
rect	53	151	54	152
rect	54	151	55	152
rect	56	151	57	152
rect	57	151	58	152
rect	59	151	60	152
rect	60	151	61	152
rect	62	151	63	152
rect	63	151	64	152
rect	64	151	65	152
rect	65	151	66	152
rect	66	151	67	152
rect	67	151	68	152
rect	68	151	69	152
rect	69	151	70	152
rect	71	151	72	152
rect	72	151	73	152
rect	73	151	74	152
rect	74	151	75	152
rect	75	151	76	152
rect	76	151	77	152
rect	77	151	78	152
rect	78	151	79	152
rect	79	151	80	152
rect	80	151	81	152
rect	81	151	82	152
rect	82	151	83	152
rect	83	151	84	152
rect	84	151	85	152
rect	85	151	86	152
rect	86	151	87	152
rect	87	151	88	152
rect	88	151	89	152
rect	89	151	90	152
rect	90	151	91	152
rect	91	151	92	152
rect	92	151	93	152
rect	93	151	94	152
rect	94	151	95	152
rect	96	151	97	152
rect	97	151	98	152
rect	99	151	100	152
rect	100	151	101	152
rect	101	151	102	152
rect	102	151	103	152
rect	103	151	104	152
rect	104	151	105	152
rect	105	151	106	152
rect	106	151	107	152
rect	108	151	109	152
rect	109	151	110	152
rect	110	151	111	152
rect	111	151	112	152
rect	129	151	130	152
rect	153	151	154	152
rect	154	151	155	152
rect	155	151	156	152
rect	156	151	157	152
rect	157	151	158	152
rect	159	151	160	152
rect	160	151	161	152
rect	175	151	176	152
rect	176	151	177	152
rect	177	151	178	152
rect	178	151	179	152
rect	179	151	180	152
rect	181	151	182	152
rect	182	151	183	152
rect	184	151	185	152
rect	185	151	186	152
rect	187	151	188	152
rect	188	151	189	152
rect	190	151	191	152
rect	191	151	192	152
rect	196	151	197	152
rect	197	151	198	152
rect	198	151	199	152
rect	199	151	200	152
rect	200	151	201	152
rect	202	151	203	152
rect	203	151	204	152
rect	205	151	206	152
rect	206	151	207	152
rect	208	151	209	152
rect	209	151	210	152
rect	211	151	212	152
rect	212	151	213	152
rect	220	151	221	152
rect	221	151	222	152
rect	222	151	223	152
rect	223	151	224	152
rect	224	151	225	152
rect	226	151	227	152
rect	227	151	228	152
rect	229	151	230	152
rect	230	151	231	152
rect	232	151	233	152
rect	233	151	234	152
rect	235	151	236	152
rect	236	151	237	152
rect	238	151	239	152
rect	239	151	240	152
rect	240	151	241	152
rect	241	151	242	152
rect	242	151	243	152
rect	243	151	244	152
rect	244	151	245	152
rect	245	151	246	152
rect	250	151	251	152
rect	251	151	252	152
rect	252	151	253	152
rect	253	151	254	152
rect	254	151	255	152
rect	256	151	257	152
rect	257	151	258	152
rect	283	151	284	152
rect	284	151	285	152
rect	285	151	286	152
rect	286	151	287	152
rect	287	151	288	152
rect	289	151	290	152
rect	290	151	291	152
rect	292	151	293	152
rect	293	151	294	152
rect	304	151	305	152
rect	305	151	306	152
rect	307	151	308	152
rect	308	151	309	152
rect	310	151	311	152
rect	311	151	312	152
rect	313	151	314	152
rect	314	151	315	152
rect	316	151	317	152
rect	317	151	318	152
rect	322	151	323	152
rect	323	151	324	152
rect	324	151	325	152
rect	325	151	326	152
rect	326	151	327	152
rect	328	151	329	152
rect	329	151	330	152
rect	340	151	341	152
rect	341	151	342	152
rect	342	151	343	152
rect	343	151	344	152
rect	344	151	345	152
rect	345	151	346	152
rect	347	151	348	152
rect	348	151	349	152
rect	350	151	351	152
rect	351	151	352	152
rect	353	151	354	152
rect	354	151	355	152
rect	355	151	356	152
rect	356	151	357	152
rect	357	151	358	152
rect	358	151	359	152
rect	359	151	360	152
rect	360	151	361	152
rect	361	151	362	152
rect	362	151	363	152
rect	364	151	365	152
rect	365	151	366	152
rect	366	151	367	152
rect	22	153	23	154
rect	23	153	24	154
rect	24	153	25	154
rect	25	153	26	154
rect	26	153	27	154
rect	27	153	28	154
rect	28	153	29	154
rect	29	153	30	154
rect	31	153	32	154
rect	32	153	33	154
rect	33	153	34	154
rect	34	153	35	154
rect	35	153	36	154
rect	36	153	37	154
rect	37	153	38	154
rect	38	153	39	154
rect	40	153	41	154
rect	41	153	42	154
rect	42	153	43	154
rect	43	153	44	154
rect	44	153	45	154
rect	45	153	46	154
rect	46	153	47	154
rect	48	153	49	154
rect	49	153	50	154
rect	50	153	51	154
rect	51	153	52	154
rect	52	153	53	154
rect	53	153	54	154
rect	54	153	55	154
rect	59	153	60	154
rect	60	153	61	154
rect	62	153	63	154
rect	63	153	64	154
rect	64	153	65	154
rect	76	153	77	154
rect	77	153	78	154
rect	78	153	79	154
rect	79	153	80	154
rect	80	153	81	154
rect	81	153	82	154
rect	82	153	83	154
rect	83	153	84	154
rect	84	153	85	154
rect	85	153	86	154
rect	86	153	87	154
rect	87	153	88	154
rect	88	153	89	154
rect	89	153	90	154
rect	90	153	91	154
rect	91	153	92	154
rect	92	153	93	154
rect	93	153	94	154
rect	94	153	95	154
rect	96	153	97	154
rect	97	153	98	154
rect	99	153	100	154
rect	100	153	101	154
rect	101	153	102	154
rect	102	153	103	154
rect	103	153	104	154
rect	104	153	105	154
rect	105	153	106	154
rect	106	153	107	154
rect	108	153	109	154
rect	109	153	110	154
rect	110	153	111	154
rect	111	153	112	154
rect	112	153	113	154
rect	113	153	114	154
rect	114	153	115	154
rect	115	153	116	154
rect	117	153	118	154
rect	118	153	119	154
rect	120	153	121	154
rect	121	153	122	154
rect	122	153	123	154
rect	123	153	124	154
rect	124	153	125	154
rect	125	153	126	154
rect	126	153	127	154
rect	127	153	128	154
rect	129	153	130	154
rect	130	153	131	154
rect	131	153	132	154
rect	132	153	133	154
rect	133	153	134	154
rect	134	153	135	154
rect	135	153	136	154
rect	136	153	137	154
rect	138	153	139	154
rect	139	153	140	154
rect	141	153	142	154
rect	142	153	143	154
rect	143	153	144	154
rect	144	153	145	154
rect	145	153	146	154
rect	146	153	147	154
rect	147	153	148	154
rect	148	153	149	154
rect	150	153	151	154
rect	151	153	152	154
rect	152	153	153	154
rect	153	153	154	154
rect	154	153	155	154
rect	155	153	156	154
rect	156	153	157	154
rect	157	153	158	154
rect	159	153	160	154
rect	160	153	161	154
rect	162	153	163	154
rect	163	153	164	154
rect	165	153	166	154
rect	166	153	167	154
rect	168	153	169	154
rect	169	153	170	154
rect	170	153	171	154
rect	171	153	172	154
rect	172	153	173	154
rect	173	153	174	154
rect	174	153	175	154
rect	175	153	176	154
rect	176	153	177	154
rect	177	153	178	154
rect	178	153	179	154
rect	179	153	180	154
rect	181	153	182	154
rect	182	153	183	154
rect	184	153	185	154
rect	185	153	186	154
rect	187	153	188	154
rect	188	153	189	154
rect	190	153	191	154
rect	191	153	192	154
rect	193	153	194	154
rect	194	153	195	154
rect	195	153	196	154
rect	196	153	197	154
rect	197	153	198	154
rect	198	153	199	154
rect	199	153	200	154
rect	200	153	201	154
rect	202	153	203	154
rect	203	153	204	154
rect	205	153	206	154
rect	206	153	207	154
rect	208	153	209	154
rect	209	153	210	154
rect	211	153	212	154
rect	212	153	213	154
rect	214	153	215	154
rect	215	153	216	154
rect	217	153	218	154
rect	218	153	219	154
rect	219	153	220	154
rect	220	153	221	154
rect	221	153	222	154
rect	222	153	223	154
rect	223	153	224	154
rect	224	153	225	154
rect	226	153	227	154
rect	227	153	228	154
rect	229	153	230	154
rect	230	153	231	154
rect	232	153	233	154
rect	233	153	234	154
rect	235	153	236	154
rect	236	153	237	154
rect	238	153	239	154
rect	239	153	240	154
rect	240	153	241	154
rect	241	153	242	154
rect	242	153	243	154
rect	243	153	244	154
rect	244	153	245	154
rect	245	153	246	154
rect	247	153	248	154
rect	248	153	249	154
rect	249	153	250	154
rect	250	153	251	154
rect	251	153	252	154
rect	252	153	253	154
rect	253	153	254	154
rect	254	153	255	154
rect	256	153	257	154
rect	257	153	258	154
rect	259	153	260	154
rect	260	153	261	154
rect	262	153	263	154
rect	263	153	264	154
rect	265	153	266	154
rect	266	153	267	154
rect	268	153	269	154
rect	269	153	270	154
rect	270	153	271	154
rect	271	153	272	154
rect	272	153	273	154
rect	274	153	275	154
rect	275	153	276	154
rect	277	153	278	154
rect	278	153	279	154
rect	280	153	281	154
rect	281	153	282	154
rect	282	153	283	154
rect	283	153	284	154
rect	284	153	285	154
rect	285	153	286	154
rect	286	153	287	154
rect	287	153	288	154
rect	289	153	290	154
rect	290	153	291	154
rect	292	153	293	154
rect	293	153	294	154
rect	295	153	296	154
rect	296	153	297	154
rect	298	153	299	154
rect	299	153	300	154
rect	301	153	302	154
rect	302	153	303	154
rect	303	153	304	154
rect	304	153	305	154
rect	305	153	306	154
rect	307	153	308	154
rect	308	153	309	154
rect	310	153	311	154
rect	311	153	312	154
rect	313	153	314	154
rect	314	153	315	154
rect	316	153	317	154
rect	317	153	318	154
rect	319	153	320	154
rect	320	153	321	154
rect	321	153	322	154
rect	322	153	323	154
rect	323	153	324	154
rect	324	153	325	154
rect	325	153	326	154
rect	326	153	327	154
rect	328	153	329	154
rect	329	153	330	154
rect	331	153	332	154
rect	332	153	333	154
rect	333	153	334	154
rect	334	153	335	154
rect	335	153	336	154
rect	337	153	338	154
rect	338	153	339	154
rect	339	153	340	154
rect	340	153	341	154
rect	341	153	342	154
rect	342	153	343	154
rect	343	153	344	154
rect	344	153	345	154
rect	345	153	346	154
rect	347	153	348	154
rect	348	153	349	154
rect	350	153	351	154
rect	351	153	352	154
rect	353	153	354	154
rect	354	153	355	154
rect	355	153	356	154
rect	356	153	357	154
rect	357	153	358	154
rect	388	153	389	154
rect	389	153	390	154
rect	390	153	391	154
rect	397	153	398	154
rect	398	153	399	154
rect	399	153	400	154
rect	400	153	401	154
rect	401	153	402	154
rect	31	155	32	156
rect	32	155	33	156
rect	33	155	34	156
rect	34	155	35	156
rect	40	155	41	156
rect	41	155	42	156
rect	42	155	43	156
rect	43	155	44	156
rect	57	155	58	156
rect	58	155	59	156
rect	59	155	60	156
rect	60	155	61	156
rect	71	155	72	156
rect	72	155	73	156
rect	73	155	74	156
rect	74	155	75	156
rect	76	155	77	156
rect	77	155	78	156
rect	78	155	79	156
rect	79	155	80	156
rect	80	155	81	156
rect	81	155	82	156
rect	82	155	83	156
rect	83	155	84	156
rect	84	155	85	156
rect	85	155	86	156
rect	86	155	87	156
rect	87	155	88	156
rect	88	155	89	156
rect	89	155	90	156
rect	90	155	91	156
rect	91	155	92	156
rect	92	155	93	156
rect	93	155	94	156
rect	94	155	95	156
rect	96	155	97	156
rect	97	155	98	156
rect	99	155	100	156
rect	100	155	101	156
rect	101	155	102	156
rect	102	155	103	156
rect	103	155	104	156
rect	104	155	105	156
rect	105	155	106	156
rect	106	155	107	156
rect	108	155	109	156
rect	109	155	110	156
rect	110	155	111	156
rect	111	155	112	156
rect	112	155	113	156
rect	113	155	114	156
rect	114	155	115	156
rect	115	155	116	156
rect	117	155	118	156
rect	118	155	119	156
rect	120	155	121	156
rect	121	155	122	156
rect	122	155	123	156
rect	123	155	124	156
rect	124	155	125	156
rect	125	155	126	156
rect	126	155	127	156
rect	127	155	128	156
rect	129	155	130	156
rect	130	155	131	156
rect	131	155	132	156
rect	132	155	133	156
rect	133	155	134	156
rect	134	155	135	156
rect	135	155	136	156
rect	136	155	137	156
rect	138	155	139	156
rect	139	155	140	156
rect	141	155	142	156
rect	142	155	143	156
rect	143	155	144	156
rect	144	155	145	156
rect	145	155	146	156
rect	146	155	147	156
rect	147	155	148	156
rect	148	155	149	156
rect	150	155	151	156
rect	151	155	152	156
rect	152	155	153	156
rect	153	155	154	156
rect	154	155	155	156
rect	155	155	156	156
rect	156	155	157	156
rect	157	155	158	156
rect	159	155	160	156
rect	160	155	161	156
rect	162	155	163	156
rect	163	155	164	156
rect	165	155	166	156
rect	166	155	167	156
rect	168	155	169	156
rect	169	155	170	156
rect	170	155	171	156
rect	171	155	172	156
rect	172	155	173	156
rect	173	155	174	156
rect	174	155	175	156
rect	175	155	176	156
rect	176	155	177	156
rect	177	155	178	156
rect	178	155	179	156
rect	179	155	180	156
rect	181	155	182	156
rect	182	155	183	156
rect	184	155	185	156
rect	185	155	186	156
rect	187	155	188	156
rect	188	155	189	156
rect	190	155	191	156
rect	191	155	192	156
rect	193	155	194	156
rect	194	155	195	156
rect	195	155	196	156
rect	196	155	197	156
rect	197	155	198	156
rect	198	155	199	156
rect	199	155	200	156
rect	200	155	201	156
rect	202	155	203	156
rect	203	155	204	156
rect	205	155	206	156
rect	206	155	207	156
rect	208	155	209	156
rect	209	155	210	156
rect	211	155	212	156
rect	212	155	213	156
rect	214	155	215	156
rect	215	155	216	156
rect	217	155	218	156
rect	218	155	219	156
rect	219	155	220	156
rect	220	155	221	156
rect	221	155	222	156
rect	222	155	223	156
rect	223	155	224	156
rect	224	155	225	156
rect	226	155	227	156
rect	227	155	228	156
rect	229	155	230	156
rect	230	155	231	156
rect	232	155	233	156
rect	233	155	234	156
rect	235	155	236	156
rect	236	155	237	156
rect	238	155	239	156
rect	239	155	240	156
rect	240	155	241	156
rect	241	155	242	156
rect	242	155	243	156
rect	243	155	244	156
rect	244	155	245	156
rect	245	155	246	156
rect	247	155	248	156
rect	248	155	249	156
rect	249	155	250	156
rect	250	155	251	156
rect	251	155	252	156
rect	252	155	253	156
rect	253	155	254	156
rect	254	155	255	156
rect	256	155	257	156
rect	257	155	258	156
rect	259	155	260	156
rect	260	155	261	156
rect	262	155	263	156
rect	263	155	264	156
rect	265	155	266	156
rect	266	155	267	156
rect	268	155	269	156
rect	269	155	270	156
rect	270	155	271	156
rect	271	155	272	156
rect	272	155	273	156
rect	274	155	275	156
rect	275	155	276	156
rect	277	155	278	156
rect	278	155	279	156
rect	280	155	281	156
rect	281	155	282	156
rect	282	155	283	156
rect	283	155	284	156
rect	284	155	285	156
rect	285	155	286	156
rect	286	155	287	156
rect	287	155	288	156
rect	289	155	290	156
rect	290	155	291	156
rect	292	155	293	156
rect	293	155	294	156
rect	295	155	296	156
rect	296	155	297	156
rect	298	155	299	156
rect	299	155	300	156
rect	301	155	302	156
rect	302	155	303	156
rect	303	155	304	156
rect	304	155	305	156
rect	305	155	306	156
rect	307	155	308	156
rect	308	155	309	156
rect	310	155	311	156
rect	311	155	312	156
rect	313	155	314	156
rect	314	155	315	156
rect	316	155	317	156
rect	317	155	318	156
rect	319	155	320	156
rect	320	155	321	156
rect	321	155	322	156
rect	322	155	323	156
rect	323	155	324	156
rect	337	155	338	156
rect	338	155	339	156
rect	339	155	340	156
rect	340	155	341	156
rect	341	155	342	156
rect	342	155	343	156
rect	343	155	344	156
rect	344	155	345	156
rect	345	155	346	156
rect	347	155	348	156
rect	348	155	349	156
rect	350	155	351	156
rect	351	155	352	156
rect	353	155	354	156
rect	354	155	355	156
rect	364	155	365	156
rect	365	155	366	156
rect	366	155	367	156
rect	368	155	369	156
rect	369	155	370	156
rect	371	155	372	156
rect	372	155	373	156
rect	374	155	375	156
rect	379	155	380	156
rect	380	155	381	156
rect	381	155	382	156
rect	383	155	384	156
rect	384	155	385	156
rect	385	155	386	156
rect	386	155	387	156
rect	387	155	388	156
rect	388	155	389	156
rect	389	155	390	156
rect	390	155	391	156
rect	392	155	393	156
rect	393	155	394	156
rect	414	155	415	156
rect	415	155	416	156
rect	416	155	417	156
rect	417	155	418	156
rect	418	155	419	156
rect	249	164	250	165
rect	250	164	251	165
rect	251	164	252	165
rect	252	164	253	165
rect	253	164	254	165
rect	254	164	255	165
rect	256	164	257	165
rect	257	164	258	165
rect	259	164	260	165
rect	260	164	261	165
rect	262	164	263	165
rect	263	164	264	165
rect	265	164	266	165
rect	266	164	267	165
rect	267	164	268	165
rect	268	164	269	165
rect	269	164	270	165
rect	270	164	271	165
rect	271	164	272	165
rect	272	164	273	165
rect	277	164	278	165
rect	278	164	279	165
rect	280	164	281	165
rect	331	164	332	165
rect	243	166	244	167
rect	244	166	245	167
rect	245	166	246	167
rect	276	166	277	167
rect	277	166	278	167
rect	278	166	279	167
rect	280	166	281	167
rect	282	166	283	167
rect	283	166	284	167
rect	284	166	285	167
rect	285	166	286	167
rect	286	166	287	167
rect	287	166	288	167
rect	289	166	290	167
rect	290	166	291	167
rect	292	166	293	167
rect	293	166	294	167
rect	295	166	296	167
rect	296	166	297	167
rect	298	166	299	167
rect	299	166	300	167
rect	300	166	301	167
rect	301	166	302	167
rect	302	166	303	167
rect	304	166	305	167
rect	305	166	306	167
rect	307	166	308	167
rect	308	166	309	167
rect	319	166	320	167
rect	320	166	321	167
rect	322	166	323	167
rect	323	166	324	167
rect	324	166	325	167
rect	325	166	326	167
rect	326	166	327	167
rect	328	166	329	167
rect	246	168	247	169
rect	247	168	248	169
rect	249	168	250	169
rect	250	168	251	169
rect	251	168	252	169
rect	252	168	253	169
rect	253	168	254	169
rect	254	168	255	169
rect	270	168	271	169
rect	271	168	272	169
rect	272	168	273	169
rect	273	168	274	169
rect	274	168	275	169
rect	276	168	277	169
rect	277	168	278	169
rect	278	168	279	169
rect	307	168	308	169
rect	308	168	309	169
rect	309	168	310	169
rect	310	168	311	169
rect	311	168	312	169
rect	313	168	314	169
rect	314	168	315	169
rect	316	168	317	169
rect	317	168	318	169
rect	318	168	319	169
rect	319	168	320	169
rect	320	168	321	169
rect	232	170	233	171
rect	233	170	234	171
rect	235	170	236	171
rect	236	170	237	171
rect	238	170	239	171
rect	239	170	240	171
rect	241	170	242	171
rect	243	170	244	171
rect	244	170	245	171
rect	246	170	247	171
rect	247	170	248	171
rect	249	170	250	171
rect	250	170	251	171
rect	265	170	266	171
rect	266	170	267	171
rect	267	170	268	171
rect	268	170	269	171
rect	270	170	271	171
rect	271	170	272	171
rect	272	170	273	171
rect	273	170	274	171
rect	274	170	275	171
rect	276	170	277	171
rect	277	170	278	171
rect	298	170	299	171
rect	299	170	300	171
rect	300	170	301	171
rect	301	170	302	171
rect	302	170	303	171
rect	304	170	305	171
rect	316	170	317	171
rect	208	172	209	173
rect	209	172	210	173
rect	211	172	212	173
rect	212	172	213	173
rect	214	172	215	173
rect	215	172	216	173
rect	217	172	218	173
rect	218	172	219	173
rect	220	172	221	173
rect	221	172	222	173
rect	222	172	223	173
rect	223	172	224	173
rect	224	172	225	173
rect	226	172	227	173
rect	227	172	228	173
rect	229	172	230	173
rect	235	172	236	173
rect	236	172	237	173
rect	238	172	239	173
rect	239	172	240	173
rect	241	172	242	173
rect	243	172	244	173
rect	244	172	245	173
rect	246	172	247	173
rect	247	172	248	173
rect	249	172	250	173
rect	250	172	251	173
rect	252	172	253	173
rect	253	172	254	173
rect	259	172	260	173
rect	260	172	261	173
rect	262	172	263	173
rect	263	172	264	173
rect	264	172	265	173
rect	265	172	266	173
rect	273	172	274	173
rect	274	172	275	173
rect	276	172	277	173
rect	277	172	278	173
rect	279	172	280	173
rect	280	172	281	173
rect	282	172	283	173
rect	283	172	284	173
rect	284	172	285	173
rect	285	172	286	173
rect	286	172	287	173
rect	287	172	288	173
rect	289	172	290	173
rect	290	172	291	173
rect	292	172	293	173
rect	293	172	294	173
rect	295	172	296	173
rect	296	172	297	173
rect	297	172	298	173
rect	298	172	299	173
rect	299	172	300	173
rect	300	172	301	173
rect	301	172	302	173
rect	302	172	303	173
rect	304	172	305	173
rect	306	172	307	173
rect	307	172	308	173
rect	308	172	309	173
rect	309	172	310	173
rect	310	172	311	173
rect	311	172	312	173
rect	313	172	314	173
rect	314	172	315	173
rect	315	172	316	173
rect	316	172	317	173
rect	318	172	319	173
rect	319	172	320	173
rect	320	172	321	173
rect	321	172	322	173
rect	322	172	323	173
rect	323	172	324	173
rect	324	172	325	173
rect	325	172	326	173
rect	326	172	327	173
rect	328	172	329	173
rect	330	172	331	173
rect	331	172	332	173
rect	333	172	334	173
rect	334	172	335	173
rect	335	172	336	173
rect	336	172	337	173
rect	337	172	338	173
rect	338	172	339	173
rect	339	172	340	173
rect	340	172	341	173
rect	341	172	342	173
rect	342	172	343	173
rect	343	172	344	173
rect	344	172	345	173
rect	345	172	346	173
rect	347	172	348	173
rect	348	172	349	173
rect	350	172	351	173
rect	351	172	352	173
rect	352	172	353	173
rect	353	172	354	173
rect	354	172	355	173
rect	355	172	356	173
rect	356	172	357	173
rect	357	172	358	173
rect	359	172	360	173
rect	360	172	361	173
rect	361	172	362	173
rect	362	172	363	173
rect	363	172	364	173
rect	364	172	365	173
rect	365	172	366	173
rect	366	172	367	173
rect	368	172	369	173
rect	369	172	370	173
rect	371	172	372	173
rect	372	172	373	173
rect	51	174	52	175
rect	52	174	53	175
rect	53	174	54	175
rect	54	174	55	175
rect	55	174	56	175
rect	57	174	58	175
rect	58	174	59	175
rect	59	174	60	175
rect	60	174	61	175
rect	61	174	62	175
rect	62	174	63	175
rect	63	174	64	175
rect	64	174	65	175
rect	66	174	67	175
rect	67	174	68	175
rect	68	174	69	175
rect	69	174	70	175
rect	70	174	71	175
rect	71	174	72	175
rect	72	174	73	175
rect	73	174	74	175
rect	74	174	75	175
rect	75	174	76	175
rect	76	174	77	175
rect	77	174	78	175
rect	78	174	79	175
rect	79	174	80	175
rect	80	174	81	175
rect	81	174	82	175
rect	82	174	83	175
rect	83	174	84	175
rect	84	174	85	175
rect	85	174	86	175
rect	86	174	87	175
rect	87	174	88	175
rect	88	174	89	175
rect	89	174	90	175
rect	90	174	91	175
rect	91	174	92	175
rect	92	174	93	175
rect	93	174	94	175
rect	94	174	95	175
rect	96	174	97	175
rect	97	174	98	175
rect	99	174	100	175
rect	100	174	101	175
rect	101	174	102	175
rect	102	174	103	175
rect	103	174	104	175
rect	104	174	105	175
rect	105	174	106	175
rect	106	174	107	175
rect	108	174	109	175
rect	109	174	110	175
rect	110	174	111	175
rect	111	174	112	175
rect	112	174	113	175
rect	113	174	114	175
rect	114	174	115	175
rect	115	174	116	175
rect	117	174	118	175
rect	118	174	119	175
rect	120	174	121	175
rect	121	174	122	175
rect	122	174	123	175
rect	123	174	124	175
rect	124	174	125	175
rect	125	174	126	175
rect	126	174	127	175
rect	127	174	128	175
rect	129	174	130	175
rect	130	174	131	175
rect	131	174	132	175
rect	132	174	133	175
rect	133	174	134	175
rect	134	174	135	175
rect	135	174	136	175
rect	136	174	137	175
rect	138	174	139	175
rect	139	174	140	175
rect	141	174	142	175
rect	142	174	143	175
rect	143	174	144	175
rect	144	174	145	175
rect	145	174	146	175
rect	146	174	147	175
rect	147	174	148	175
rect	148	174	149	175
rect	150	174	151	175
rect	151	174	152	175
rect	152	174	153	175
rect	153	174	154	175
rect	154	174	155	175
rect	155	174	156	175
rect	156	174	157	175
rect	157	174	158	175
rect	159	174	160	175
rect	160	174	161	175
rect	162	174	163	175
rect	163	174	164	175
rect	165	174	166	175
rect	166	174	167	175
rect	168	174	169	175
rect	169	174	170	175
rect	170	174	171	175
rect	171	174	172	175
rect	172	174	173	175
rect	174	174	175	175
rect	175	174	176	175
rect	176	174	177	175
rect	178	174	179	175
rect	179	174	180	175
rect	180	174	181	175
rect	181	174	182	175
rect	182	174	183	175
rect	184	174	185	175
rect	185	174	186	175
rect	187	174	188	175
rect	188	174	189	175
rect	190	174	191	175
rect	191	174	192	175
rect	193	174	194	175
rect	194	174	195	175
rect	195	174	196	175
rect	196	174	197	175
rect	197	174	198	175
rect	198	174	199	175
rect	199	174	200	175
rect	200	174	201	175
rect	202	174	203	175
rect	203	174	204	175
rect	205	174	206	175
rect	206	174	207	175
rect	207	174	208	175
rect	208	174	209	175
rect	209	174	210	175
rect	211	174	212	175
rect	212	174	213	175
rect	214	174	215	175
rect	215	174	216	175
rect	217	174	218	175
rect	218	174	219	175
rect	220	174	221	175
rect	221	174	222	175
rect	222	174	223	175
rect	223	174	224	175
rect	224	174	225	175
rect	226	174	227	175
rect	227	174	228	175
rect	229	174	230	175
rect	231	174	232	175
rect	232	174	233	175
rect	233	174	234	175
rect	234	174	235	175
rect	235	174	236	175
rect	236	174	237	175
rect	238	174	239	175
rect	239	174	240	175
rect	241	174	242	175
rect	243	174	244	175
rect	244	174	245	175
rect	246	174	247	175
rect	247	174	248	175
rect	249	174	250	175
rect	250	174	251	175
rect	252	174	253	175
rect	253	174	254	175
rect	255	174	256	175
rect	256	174	257	175
rect	257	174	258	175
rect	258	174	259	175
rect	259	174	260	175
rect	260	174	261	175
rect	262	174	263	175
rect	263	174	264	175
rect	264	174	265	175
rect	265	174	266	175
rect	267	174	268	175
rect	268	174	269	175
rect	270	174	271	175
rect	271	174	272	175
rect	273	174	274	175
rect	274	174	275	175
rect	276	174	277	175
rect	277	174	278	175
rect	279	174	280	175
rect	280	174	281	175
rect	282	174	283	175
rect	283	174	284	175
rect	284	174	285	175
rect	285	174	286	175
rect	286	174	287	175
rect	287	174	288	175
rect	289	174	290	175
rect	290	174	291	175
rect	295	174	296	175
rect	296	174	297	175
rect	297	174	298	175
rect	298	174	299	175
rect	299	174	300	175
rect	300	174	301	175
rect	301	174	302	175
rect	302	174	303	175
rect	304	174	305	175
rect	306	174	307	175
rect	307	174	308	175
rect	308	174	309	175
rect	309	174	310	175
rect	310	174	311	175
rect	311	174	312	175
rect	313	174	314	175
rect	150	176	151	177
rect	151	176	152	177
rect	193	176	194	177
rect	194	176	195	177
rect	195	176	196	177
rect	196	176	197	177
rect	197	176	198	177
rect	198	176	199	177
rect	199	176	200	177
rect	200	176	201	177
rect	202	176	203	177
rect	203	176	204	177
rect	205	176	206	177
rect	206	176	207	177
rect	207	176	208	177
rect	220	176	221	177
rect	221	176	222	177
rect	222	176	223	177
rect	223	176	224	177
rect	224	176	225	177
rect	226	176	227	177
rect	227	176	228	177
rect	229	176	230	177
rect	231	176	232	177
rect	232	176	233	177
rect	233	176	234	177
rect	234	176	235	177
rect	235	176	236	177
rect	236	176	237	177
rect	238	176	239	177
rect	239	176	240	177
rect	241	176	242	177
rect	243	176	244	177
rect	244	176	245	177
rect	246	176	247	177
rect	247	176	248	177
rect	249	176	250	177
rect	250	176	251	177
rect	252	176	253	177
rect	253	176	254	177
rect	255	176	256	177
rect	256	176	257	177
rect	257	176	258	177
rect	258	176	259	177
rect	259	176	260	177
rect	260	176	261	177
rect	262	176	263	177
rect	263	176	264	177
rect	264	176	265	177
rect	265	176	266	177
rect	267	176	268	177
rect	268	176	269	177
rect	270	176	271	177
rect	271	176	272	177
rect	273	176	274	177
rect	274	176	275	177
rect	276	176	277	177
rect	277	176	278	177
rect	279	176	280	177
rect	280	176	281	177
rect	282	176	283	177
rect	283	176	284	177
rect	284	176	285	177
rect	285	176	286	177
rect	286	176	287	177
rect	287	176	288	177
rect	289	176	290	177
rect	294	176	295	177
rect	295	176	296	177
rect	296	176	297	177
rect	297	176	298	177
rect	298	176	299	177
rect	299	176	300	177
rect	300	176	301	177
rect	301	176	302	177
rect	302	176	303	177
rect	304	176	305	177
rect	306	176	307	177
rect	307	176	308	177
rect	308	176	309	177
rect	309	176	310	177
rect	310	176	311	177
rect	311	176	312	177
rect	354	176	355	177
rect	355	176	356	177
rect	356	176	357	177
rect	357	176	358	177
rect	359	176	360	177
rect	360	176	361	177
rect	361	176	362	177
rect	362	176	363	177
rect	363	176	364	177
rect	364	176	365	177
rect	365	176	366	177
rect	366	176	367	177
rect	138	178	139	179
rect	139	178	140	179
rect	141	178	142	179
rect	142	178	143	179
rect	143	178	144	179
rect	144	178	145	179
rect	145	178	146	179
rect	146	178	147	179
rect	147	178	148	179
rect	148	178	149	179
rect	178	178	179	179
rect	179	178	180	179
rect	180	178	181	179
rect	181	178	182	179
rect	182	178	183	179
rect	193	178	194	179
rect	194	178	195	179
rect	195	178	196	179
rect	196	178	197	179
rect	197	178	198	179
rect	198	178	199	179
rect	199	178	200	179
rect	200	178	201	179
rect	214	178	215	179
rect	215	178	216	179
rect	217	178	218	179
rect	218	178	219	179
rect	219	178	220	179
rect	220	178	221	179
rect	221	178	222	179
rect	222	178	223	179
rect	223	178	224	179
rect	224	178	225	179
rect	226	178	227	179
rect	227	178	228	179
rect	229	178	230	179
rect	231	178	232	179
rect	232	178	233	179
rect	238	178	239	179
rect	239	178	240	179
rect	241	178	242	179
rect	243	178	244	179
rect	244	178	245	179
rect	246	178	247	179
rect	247	178	248	179
rect	249	178	250	179
rect	250	178	251	179
rect	252	178	253	179
rect	253	178	254	179
rect	255	178	256	179
rect	256	178	257	179
rect	264	178	265	179
rect	265	178	266	179
rect	267	178	268	179
rect	268	178	269	179
rect	270	178	271	179
rect	271	178	272	179
rect	273	178	274	179
rect	274	178	275	179
rect	276	178	277	179
rect	277	178	278	179
rect	279	178	280	179
rect	280	178	281	179
rect	282	178	283	179
rect	283	178	284	179
rect	284	178	285	179
rect	285	178	286	179
rect	286	178	287	179
rect	287	178	288	179
rect	289	178	290	179
rect	291	178	292	179
rect	292	178	293	179
rect	294	178	295	179
rect	295	178	296	179
rect	296	178	297	179
rect	297	178	298	179
rect	298	178	299	179
rect	299	178	300	179
rect	300	178	301	179
rect	301	178	302	179
rect	302	178	303	179
rect	304	178	305	179
rect	306	178	307	179
rect	307	178	308	179
rect	308	178	309	179
rect	309	178	310	179
rect	310	178	311	179
rect	311	178	312	179
rect	312	178	313	179
rect	313	178	314	179
rect	315	178	316	179
rect	316	178	317	179
rect	318	178	319	179
rect	319	178	320	179
rect	320	178	321	179
rect	321	178	322	179
rect	322	178	323	179
rect	323	178	324	179
rect	324	178	325	179
rect	325	178	326	179
rect	326	178	327	179
rect	345	178	346	179
rect	347	178	348	179
rect	348	178	349	179
rect	369	178	370	179
rect	371	178	372	179
rect	372	178	373	179
rect	373	178	374	179
rect	374	178	375	179
rect	375	178	376	179
rect	376	178	377	179
rect	377	178	378	179
rect	378	178	379	179
rect	379	178	380	179
rect	380	178	381	179
rect	381	178	382	179
rect	43	180	44	181
rect	129	180	130	181
rect	130	180	131	181
rect	131	180	132	181
rect	132	180	133	181
rect	133	180	134	181
rect	134	180	135	181
rect	135	180	136	181
rect	136	180	137	181
rect	174	180	175	181
rect	175	180	176	181
rect	176	180	177	181
rect	177	180	178	181
rect	178	180	179	181
rect	179	180	180	181
rect	180	180	181	181
rect	181	180	182	181
rect	182	180	183	181
rect	183	180	184	181
rect	184	180	185	181
rect	185	180	186	181
rect	187	180	188	181
rect	188	180	189	181
rect	190	180	191	181
rect	191	180	192	181
rect	193	180	194	181
rect	194	180	195	181
rect	195	180	196	181
rect	196	180	197	181
rect	197	180	198	181
rect	198	180	199	181
rect	199	180	200	181
rect	200	180	201	181
rect	201	180	202	181
rect	202	180	203	181
rect	203	180	204	181
rect	204	180	205	181
rect	206	180	207	181
rect	207	180	208	181
rect	209	180	210	181
rect	211	180	212	181
rect	212	180	213	181
rect	213	180	214	181
rect	214	180	215	181
rect	215	180	216	181
rect	217	180	218	181
rect	218	180	219	181
rect	219	180	220	181
rect	220	180	221	181
rect	221	180	222	181
rect	222	180	223	181
rect	223	180	224	181
rect	224	180	225	181
rect	226	180	227	181
rect	227	180	228	181
rect	229	180	230	181
rect	231	180	232	181
rect	232	180	233	181
rect	234	180	235	181
rect	235	180	236	181
rect	236	180	237	181
rect	237	180	238	181
rect	238	180	239	181
rect	239	180	240	181
rect	241	180	242	181
rect	243	180	244	181
rect	244	180	245	181
rect	246	180	247	181
rect	247	180	248	181
rect	249	180	250	181
rect	250	180	251	181
rect	252	180	253	181
rect	253	180	254	181
rect	255	180	256	181
rect	256	180	257	181
rect	258	180	259	181
rect	259	180	260	181
rect	260	180	261	181
rect	262	180	263	181
rect	264	180	265	181
rect	265	180	266	181
rect	267	180	268	181
rect	268	180	269	181
rect	270	180	271	181
rect	271	180	272	181
rect	273	180	274	181
rect	274	180	275	181
rect	276	180	277	181
rect	277	180	278	181
rect	279	180	280	181
rect	280	180	281	181
rect	282	180	283	181
rect	283	180	284	181
rect	289	180	290	181
rect	291	180	292	181
rect	292	180	293	181
rect	294	180	295	181
rect	295	180	296	181
rect	342	180	343	181
rect	343	180	344	181
rect	345	180	346	181
rect	357	180	358	181
rect	358	180	359	181
rect	360	180	361	181
rect	361	180	362	181
rect	362	180	363	181
rect	363	180	364	181
rect	364	180	365	181
rect	365	180	366	181
rect	366	180	367	181
rect	367	180	368	181
rect	369	180	370	181
rect	395	180	396	181
rect	396	180	397	181
rect	36	182	37	183
rect	37	182	38	183
rect	38	182	39	183
rect	39	182	40	183
rect	40	182	41	183
rect	41	182	42	183
rect	43	182	44	183
rect	44	182	45	183
rect	99	182	100	183
rect	120	182	121	183
rect	121	182	122	183
rect	122	182	123	183
rect	123	182	124	183
rect	124	182	125	183
rect	125	182	126	183
rect	126	182	127	183
rect	127	182	128	183
rect	165	182	166	183
rect	166	182	167	183
rect	167	182	168	183
rect	169	182	170	183
rect	170	182	171	183
rect	171	182	172	183
rect	172	182	173	183
rect	173	182	174	183
rect	184	182	185	183
rect	185	182	186	183
rect	190	182	191	183
rect	191	182	192	183
rect	193	182	194	183
rect	194	182	195	183
rect	195	182	196	183
rect	196	182	197	183
rect	197	182	198	183
rect	198	182	199	183
rect	199	182	200	183
rect	200	182	201	183
rect	201	182	202	183
rect	215	182	216	183
rect	221	182	222	183
rect	222	182	223	183
rect	223	182	224	183
rect	224	182	225	183
rect	229	182	230	183
rect	231	182	232	183
rect	232	182	233	183
rect	234	182	235	183
rect	235	182	236	183
rect	236	182	237	183
rect	237	182	238	183
rect	238	182	239	183
rect	239	182	240	183
rect	262	182	263	183
rect	264	182	265	183
rect	265	182	266	183
rect	267	182	268	183
rect	268	182	269	183
rect	270	182	271	183
rect	271	182	272	183
rect	273	182	274	183
rect	274	182	275	183
rect	276	182	277	183
rect	277	182	278	183
rect	279	182	280	183
rect	280	182	281	183
rect	282	182	283	183
rect	283	182	284	183
rect	285	182	286	183
rect	286	182	287	183
rect	287	182	288	183
rect	288	182	289	183
rect	289	182	290	183
rect	291	182	292	183
rect	292	182	293	183
rect	294	182	295	183
rect	295	182	296	183
rect	297	182	298	183
rect	298	182	299	183
rect	299	182	300	183
rect	300	182	301	183
rect	301	182	302	183
rect	302	182	303	183
rect	304	182	305	183
rect	306	182	307	183
rect	307	182	308	183
rect	308	182	309	183
rect	309	182	310	183
rect	310	182	311	183
rect	311	182	312	183
rect	312	182	313	183
rect	313	182	314	183
rect	315	182	316	183
rect	316	182	317	183
rect	318	182	319	183
rect	319	182	320	183
rect	320	182	321	183
rect	321	182	322	183
rect	322	182	323	183
rect	323	182	324	183
rect	324	182	325	183
rect	325	182	326	183
rect	326	182	327	183
rect	327	182	328	183
rect	328	182	329	183
rect	330	182	331	183
rect	331	182	332	183
rect	333	182	334	183
rect	334	182	335	183
rect	335	182	336	183
rect	336	182	337	183
rect	337	182	338	183
rect	338	182	339	183
rect	339	182	340	183
rect	340	182	341	183
rect	342	182	343	183
rect	343	182	344	183
rect	345	182	346	183
rect	346	182	347	183
rect	347	182	348	183
rect	348	182	349	183
rect	349	182	350	183
rect	350	182	351	183
rect	351	182	352	183
rect	352	182	353	183
rect	354	182	355	183
rect	355	182	356	183
rect	357	182	358	183
rect	358	182	359	183
rect	360	182	361	183
rect	361	182	362	183
rect	362	182	363	183
rect	363	182	364	183
rect	364	182	365	183
rect	365	182	366	183
rect	366	182	367	183
rect	367	182	368	183
rect	369	182	370	183
rect	370	182	371	183
rect	389	182	390	183
rect	390	182	391	183
rect	395	182	396	183
rect	396	182	397	183
rect	398	182	399	183
rect	399	182	400	183
rect	400	182	401	183
rect	401	182	402	183
rect	402	182	403	183
rect	403	182	404	183
rect	404	182	405	183
rect	405	182	406	183
rect	406	182	407	183
rect	407	182	408	183
rect	408	182	409	183
rect	409	182	410	183
rect	411	182	412	183
rect	412	182	413	183
rect	9	184	10	185
rect	10	184	11	185
rect	11	184	12	185
rect	12	184	13	185
rect	13	184	14	185
rect	37	184	38	185
rect	38	184	39	185
rect	52	184	53	185
rect	53	184	54	185
rect	54	184	55	185
rect	55	184	56	185
rect	66	184	67	185
rect	96	184	97	185
rect	108	184	109	185
rect	109	184	110	185
rect	110	184	111	185
rect	111	184	112	185
rect	112	184	113	185
rect	113	184	114	185
rect	114	184	115	185
rect	115	184	116	185
rect	117	184	118	185
rect	118	184	119	185
rect	162	184	163	185
rect	163	184	164	185
rect	164	184	165	185
rect	165	184	166	185
rect	166	184	167	185
rect	167	184	168	185
rect	169	184	170	185
rect	170	184	171	185
rect	187	184	188	185
rect	188	184	189	185
rect	189	184	190	185
rect	190	184	191	185
rect	191	184	192	185
rect	193	184	194	185
rect	194	184	195	185
rect	195	184	196	185
rect	196	184	197	185
rect	197	184	198	185
rect	198	184	199	185
rect	199	184	200	185
rect	200	184	201	185
rect	201	184	202	185
rect	203	184	204	185
rect	204	184	205	185
rect	206	184	207	185
rect	207	184	208	185
rect	209	184	210	185
rect	210	184	211	185
rect	212	184	213	185
rect	213	184	214	185
rect	215	184	216	185
rect	216	184	217	185
rect	217	184	218	185
rect	218	184	219	185
rect	219	184	220	185
rect	221	184	222	185
rect	222	184	223	185
rect	223	184	224	185
rect	224	184	225	185
rect	225	184	226	185
rect	226	184	227	185
rect	227	184	228	185
rect	228	184	229	185
rect	229	184	230	185
rect	231	184	232	185
rect	232	184	233	185
rect	234	184	235	185
rect	235	184	236	185
rect	236	184	237	185
rect	237	184	238	185
rect	238	184	239	185
rect	239	184	240	185
rect	240	184	241	185
rect	241	184	242	185
rect	243	184	244	185
rect	244	184	245	185
rect	246	184	247	185
rect	247	184	248	185
rect	249	184	250	185
rect	250	184	251	185
rect	252	184	253	185
rect	253	184	254	185
rect	255	184	256	185
rect	256	184	257	185
rect	258	184	259	185
rect	259	184	260	185
rect	260	184	261	185
rect	261	184	262	185
rect	262	184	263	185
rect	264	184	265	185
rect	265	184	266	185
rect	267	184	268	185
rect	268	184	269	185
rect	270	184	271	185
rect	271	184	272	185
rect	273	184	274	185
rect	274	184	275	185
rect	276	184	277	185
rect	277	184	278	185
rect	279	184	280	185
rect	280	184	281	185
rect	282	184	283	185
rect	283	184	284	185
rect	285	184	286	185
rect	286	184	287	185
rect	287	184	288	185
rect	288	184	289	185
rect	289	184	290	185
rect	291	184	292	185
rect	292	184	293	185
rect	294	184	295	185
rect	295	184	296	185
rect	297	184	298	185
rect	298	184	299	185
rect	299	184	300	185
rect	300	184	301	185
rect	301	184	302	185
rect	302	184	303	185
rect	327	184	328	185
rect	328	184	329	185
rect	330	184	331	185
rect	331	184	332	185
rect	333	184	334	185
rect	334	184	335	185
rect	335	184	336	185
rect	336	184	337	185
rect	337	184	338	185
rect	338	184	339	185
rect	339	184	340	185
rect	340	184	341	185
rect	342	184	343	185
rect	343	184	344	185
rect	345	184	346	185
rect	346	184	347	185
rect	347	184	348	185
rect	348	184	349	185
rect	349	184	350	185
rect	350	184	351	185
rect	351	184	352	185
rect	352	184	353	185
rect	354	184	355	185
rect	355	184	356	185
rect	357	184	358	185
rect	358	184	359	185
rect	360	184	361	185
rect	361	184	362	185
rect	362	184	363	185
rect	363	184	364	185
rect	364	184	365	185
rect	365	184	366	185
rect	366	184	367	185
rect	367	184	368	185
rect	369	184	370	185
rect	370	184	371	185
rect	372	184	373	185
rect	373	184	374	185
rect	374	184	375	185
rect	375	184	376	185
rect	376	184	377	185
rect	377	184	378	185
rect	378	184	379	185
rect	379	184	380	185
rect	380	184	381	185
rect	381	184	382	185
rect	382	184	383	185
rect	383	184	384	185
rect	384	184	385	185
rect	385	184	386	185
rect	386	184	387	185
rect	387	184	388	185
rect	392	184	393	185
rect	393	184	394	185
rect	395	184	396	185
rect	396	184	397	185
rect	398	184	399	185
rect	399	184	400	185
rect	400	184	401	185
rect	401	184	402	185
rect	402	184	403	185
rect	403	184	404	185
rect	404	184	405	185
rect	405	184	406	185
rect	406	184	407	185
rect	407	184	408	185
rect	408	184	409	185
rect	409	184	410	185
rect	313	193	314	194
rect	315	193	316	194
rect	316	193	317	194
rect	318	193	319	194
rect	319	193	320	194
rect	321	193	322	194
rect	322	193	323	194
rect	323	193	324	194
rect	324	193	325	194
rect	325	193	326	194
rect	327	193	328	194
rect	328	193	329	194
rect	330	193	331	194
rect	331	193	332	194
rect	311	195	312	196
rect	313	195	314	196
rect	315	195	316	196
rect	316	195	317	196
rect	318	195	319	196
rect	319	195	320	196
rect	321	195	322	196
rect	322	195	323	196
rect	323	195	324	196
rect	324	195	325	196
rect	325	195	326	196
rect	206	197	207	198
rect	207	197	208	198
rect	209	197	210	198
rect	210	197	211	198
rect	212	197	213	198
rect	213	197	214	198
rect	215	197	216	198
rect	216	197	217	198
rect	217	197	218	198
rect	218	197	219	198
rect	219	197	220	198
rect	220	197	221	198
rect	221	197	222	198
rect	222	197	223	198
rect	223	197	224	198
rect	224	197	225	198
rect	225	197	226	198
rect	226	197	227	198
rect	318	197	319	198
rect	319	197	320	198
rect	321	197	322	198
rect	322	197	323	198
rect	323	197	324	198
rect	324	197	325	198
rect	207	199	208	200
rect	209	199	210	200
rect	210	199	211	200
rect	212	199	213	200
rect	213	199	214	200
rect	317	199	318	200
rect	318	199	319	200
rect	319	199	320	200
rect	212	201	213	202
rect	213	201	214	202
rect	214	201	215	202
rect	243	201	244	202
rect	244	201	245	202
rect	246	201	247	202
rect	247	201	248	202
rect	249	201	250	202
rect	250	201	251	202
rect	252	201	253	202
rect	253	201	254	202
rect	255	201	256	202
rect	256	201	257	202
rect	258	201	259	202
rect	259	201	260	202
rect	320	201	321	202
rect	321	201	322	202
rect	322	201	323	202
rect	323	201	324	202
rect	324	201	325	202
rect	326	201	327	202
rect	327	201	328	202
rect	328	201	329	202
rect	330	201	331	202
rect	331	201	332	202
rect	332	201	333	202
rect	333	201	334	202
rect	334	201	335	202
rect	335	201	336	202
rect	336	201	337	202
rect	337	201	338	202
rect	339	201	340	202
rect	340	201	341	202
rect	342	201	343	202
rect	343	201	344	202
rect	49	203	50	204
rect	50	203	51	204
rect	52	203	53	204
rect	53	203	54	204
rect	54	203	55	204
rect	55	203	56	204
rect	213	203	214	204
rect	214	203	215	204
rect	216	203	217	204
rect	217	203	218	204
rect	218	203	219	204
rect	219	203	220	204
rect	220	203	221	204
rect	221	203	222	204
rect	222	203	223	204
rect	223	203	224	204
rect	224	203	225	204
rect	225	203	226	204
rect	226	203	227	204
rect	227	203	228	204
rect	228	203	229	204
rect	229	203	230	204
rect	231	203	232	204
rect	232	203	233	204
rect	234	203	235	204
rect	235	203	236	204
rect	236	203	237	204
rect	237	203	238	204
rect	238	203	239	204
rect	239	203	240	204
rect	240	203	241	204
rect	241	203	242	204
rect	242	203	243	204
rect	243	203	244	204
rect	244	203	245	204
rect	246	203	247	204
rect	247	203	248	204
rect	330	203	331	204
rect	344	203	345	204
rect	345	203	346	204
rect	346	203	347	204
rect	347	203	348	204
rect	348	203	349	204
rect	349	203	350	204
rect	350	203	351	204
rect	351	203	352	204
rect	352	203	353	204
rect	354	203	355	204
rect	355	203	356	204
rect	357	203	358	204
rect	358	203	359	204
rect	360	203	361	204
rect	361	203	362	204
rect	362	203	363	204
rect	363	203	364	204
rect	364	203	365	204
rect	365	203	366	204
rect	366	203	367	204
rect	367	203	368	204
rect	46	205	47	206
rect	47	205	48	206
rect	48	205	49	206
rect	49	205	50	206
rect	50	205	51	206
rect	52	205	53	206
rect	150	205	151	206
rect	151	205	152	206
rect	153	205	154	206
rect	154	205	155	206
rect	155	205	156	206
rect	156	205	157	206
rect	157	205	158	206
rect	158	205	159	206
rect	250	205	251	206
rect	252	205	253	206
rect	253	205	254	206
rect	255	205	256	206
rect	256	205	257	206
rect	262	205	263	206
rect	263	205	264	206
rect	264	205	265	206
rect	265	205	266	206
rect	270	205	271	206
rect	271	205	272	206
rect	272	205	273	206
rect	282	205	283	206
rect	283	205	284	206
rect	284	205	285	206
rect	308	205	309	206
rect	309	205	310	206
rect	311	205	312	206
rect	313	205	314	206
rect	315	205	316	206
rect	317	205	318	206
rect	318	205	319	206
rect	320	205	321	206
rect	321	205	322	206
rect	322	205	323	206
rect	323	205	324	206
rect	324	205	325	206
rect	326	205	327	206
rect	327	205	328	206
rect	328	205	329	206
rect	329	205	330	206
rect	330	205	331	206
rect	332	205	333	206
rect	333	205	334	206
rect	334	205	335	206
rect	335	205	336	206
rect	336	205	337	206
rect	337	205	338	206
rect	339	205	340	206
rect	340	205	341	206
rect	40	207	41	208
rect	41	207	42	208
rect	43	207	44	208
rect	44	207	45	208
rect	45	207	46	208
rect	46	207	47	208
rect	120	207	121	208
rect	121	207	122	208
rect	122	207	123	208
rect	123	207	124	208
rect	124	207	125	208
rect	125	207	126	208
rect	138	207	139	208
rect	139	207	140	208
rect	141	207	142	208
rect	142	207	143	208
rect	143	207	144	208
rect	144	207	145	208
rect	145	207	146	208
rect	146	207	147	208
rect	147	207	148	208
rect	148	207	149	208
rect	149	207	150	208
rect	181	207	182	208
rect	182	207	183	208
rect	225	207	226	208
rect	226	207	227	208
rect	227	207	228	208
rect	228	207	229	208
rect	229	207	230	208
rect	231	207	232	208
rect	232	207	233	208
rect	234	207	235	208
rect	235	207	236	208
rect	236	207	237	208
rect	237	207	238	208
rect	238	207	239	208
rect	239	207	240	208
rect	240	207	241	208
rect	241	207	242	208
rect	242	207	243	208
rect	243	207	244	208
rect	244	207	245	208
rect	259	207	260	208
rect	260	207	261	208
rect	262	207	263	208
rect	263	207	264	208
rect	264	207	265	208
rect	265	207	266	208
rect	266	207	267	208
rect	267	207	268	208
rect	268	207	269	208
rect	269	207	270	208
rect	270	207	271	208
rect	271	207	272	208
rect	272	207	273	208
rect	274	207	275	208
rect	275	207	276	208
rect	276	207	277	208
rect	277	207	278	208
rect	279	207	280	208
rect	280	207	281	208
rect	281	207	282	208
rect	282	207	283	208
rect	283	207	284	208
rect	284	207	285	208
rect	286	207	287	208
rect	287	207	288	208
rect	288	207	289	208
rect	289	207	290	208
rect	313	207	314	208
rect	315	207	316	208
rect	317	207	318	208
rect	318	207	319	208
rect	320	207	321	208
rect	321	207	322	208
rect	322	207	323	208
rect	323	207	324	208
rect	324	207	325	208
rect	326	207	327	208
rect	327	207	328	208
rect	341	207	342	208
rect	342	207	343	208
rect	344	207	345	208
rect	345	207	346	208
rect	346	207	347	208
rect	347	207	348	208
rect	348	207	349	208
rect	349	207	350	208
rect	350	207	351	208
rect	351	207	352	208
rect	352	207	353	208
rect	28	209	29	210
rect	29	209	30	210
rect	31	209	32	210
rect	32	209	33	210
rect	33	209	34	210
rect	34	209	35	210
rect	35	209	36	210
rect	36	209	37	210
rect	37	209	38	210
rect	38	209	39	210
rect	39	209	40	210
rect	40	209	41	210
rect	41	209	42	210
rect	43	209	44	210
rect	44	209	45	210
rect	45	209	46	210
rect	46	209	47	210
rect	48	209	49	210
rect	49	209	50	210
rect	50	209	51	210
rect	52	209	53	210
rect	54	209	55	210
rect	55	209	56	210
rect	57	209	58	210
rect	58	209	59	210
rect	59	209	60	210
rect	60	209	61	210
rect	62	209	63	210
rect	63	209	64	210
rect	64	209	65	210
rect	65	209	66	210
rect	66	209	67	210
rect	68	209	69	210
rect	69	209	70	210
rect	70	209	71	210
rect	71	209	72	210
rect	72	209	73	210
rect	73	209	74	210
rect	74	209	75	210
rect	75	209	76	210
rect	76	209	77	210
rect	77	209	78	210
rect	78	209	79	210
rect	79	209	80	210
rect	80	209	81	210
rect	81	209	82	210
rect	82	209	83	210
rect	83	209	84	210
rect	84	209	85	210
rect	85	209	86	210
rect	86	209	87	210
rect	87	209	88	210
rect	88	209	89	210
rect	89	209	90	210
rect	90	209	91	210
rect	91	209	92	210
rect	92	209	93	210
rect	93	209	94	210
rect	94	209	95	210
rect	95	209	96	210
rect	96	209	97	210
rect	98	209	99	210
rect	99	209	100	210
rect	100	209	101	210
rect	102	209	103	210
rect	103	209	104	210
rect	104	209	105	210
rect	105	209	106	210
rect	106	209	107	210
rect	107	209	108	210
rect	108	209	109	210
rect	109	209	110	210
rect	110	209	111	210
rect	111	209	112	210
rect	112	209	113	210
rect	113	209	114	210
rect	114	209	115	210
rect	115	209	116	210
rect	117	209	118	210
rect	118	209	119	210
rect	119	209	120	210
rect	120	209	121	210
rect	121	209	122	210
rect	122	209	123	210
rect	123	209	124	210
rect	124	209	125	210
rect	125	209	126	210
rect	127	209	128	210
rect	129	209	130	210
rect	130	209	131	210
rect	131	209	132	210
rect	132	209	133	210
rect	133	209	134	210
rect	134	209	135	210
rect	135	209	136	210
rect	136	209	137	210
rect	137	209	138	210
rect	138	209	139	210
rect	139	209	140	210
rect	141	209	142	210
rect	142	209	143	210
rect	143	209	144	210
rect	144	209	145	210
rect	145	209	146	210
rect	146	209	147	210
rect	147	209	148	210
rect	148	209	149	210
rect	149	209	150	210
rect	151	209	152	210
rect	153	209	154	210
rect	154	209	155	210
rect	155	209	156	210
rect	156	209	157	210
rect	157	209	158	210
rect	158	209	159	210
rect	160	209	161	210
rect	161	209	162	210
rect	162	209	163	210
rect	163	209	164	210
rect	164	209	165	210
rect	165	209	166	210
rect	166	209	167	210
rect	167	209	168	210
rect	169	209	170	210
rect	170	209	171	210
rect	172	209	173	210
rect	173	209	174	210
rect	175	209	176	210
rect	176	209	177	210
rect	177	209	178	210
rect	178	209	179	210
rect	179	209	180	210
rect	180	209	181	210
rect	181	209	182	210
rect	182	209	183	210
rect	183	209	184	210
rect	184	209	185	210
rect	185	209	186	210
rect	187	209	188	210
rect	188	209	189	210
rect	189	209	190	210
rect	190	209	191	210
rect	191	209	192	210
rect	192	209	193	210
rect	193	209	194	210
rect	194	209	195	210
rect	195	209	196	210
rect	196	209	197	210
rect	197	209	198	210
rect	198	209	199	210
rect	199	209	200	210
rect	200	209	201	210
rect	201	209	202	210
rect	203	209	204	210
rect	204	209	205	210
rect	205	209	206	210
rect	207	209	208	210
rect	209	209	210	210
rect	210	209	211	210
rect	211	209	212	210
rect	213	209	214	210
rect	214	209	215	210
rect	216	209	217	210
rect	217	209	218	210
rect	218	209	219	210
rect	219	209	220	210
rect	220	209	221	210
rect	221	209	222	210
rect	222	209	223	210
rect	223	209	224	210
rect	225	209	226	210
rect	226	209	227	210
rect	227	209	228	210
rect	228	209	229	210
rect	229	209	230	210
rect	231	209	232	210
rect	232	209	233	210
rect	234	209	235	210
rect	235	209	236	210
rect	236	209	237	210
rect	237	209	238	210
rect	238	209	239	210
rect	239	209	240	210
rect	240	209	241	210
rect	241	209	242	210
rect	242	209	243	210
rect	243	209	244	210
rect	244	209	245	210
rect	245	209	246	210
rect	246	209	247	210
rect	247	209	248	210
rect	248	209	249	210
rect	250	209	251	210
rect	252	209	253	210
rect	253	209	254	210
rect	255	209	256	210
rect	256	209	257	210
rect	257	209	258	210
rect	259	209	260	210
rect	260	209	261	210
rect	262	209	263	210
rect	263	209	264	210
rect	268	209	269	210
rect	269	209	270	210
rect	270	209	271	210
rect	271	209	272	210
rect	272	209	273	210
rect	274	209	275	210
rect	275	209	276	210
rect	276	209	277	210
rect	277	209	278	210
rect	279	209	280	210
rect	280	209	281	210
rect	281	209	282	210
rect	282	209	283	210
rect	283	209	284	210
rect	284	209	285	210
rect	286	209	287	210
rect	287	209	288	210
rect	288	209	289	210
rect	289	209	290	210
rect	290	209	291	210
rect	291	209	292	210
rect	292	209	293	210
rect	302	209	303	210
rect	303	209	304	210
rect	305	209	306	210
rect	306	209	307	210
rect	308	209	309	210
rect	309	209	310	210
rect	311	209	312	210
rect	312	209	313	210
rect	313	209	314	210
rect	323	209	324	210
rect	324	209	325	210
rect	326	209	327	210
rect	327	209	328	210
rect	329	209	330	210
rect	330	209	331	210
rect	332	209	333	210
rect	333	209	334	210
rect	334	209	335	210
rect	335	209	336	210
rect	336	209	337	210
rect	337	209	338	210
rect	339	209	340	210
rect	341	209	342	210
rect	342	209	343	210
rect	344	209	345	210
rect	345	209	346	210
rect	346	209	347	210
rect	347	209	348	210
rect	348	209	349	210
rect	349	209	350	210
rect	350	209	351	210
rect	351	209	352	210
rect	352	209	353	210
rect	353	209	354	210
rect	354	209	355	210
rect	355	209	356	210
rect	389	209	390	210
rect	390	209	391	210
rect	392	209	393	210
rect	393	209	394	210
rect	395	209	396	210
rect	396	209	397	210
rect	15	211	16	212
rect	16	211	17	212
rect	27	211	28	212
rect	28	211	29	212
rect	29	211	30	212
rect	39	211	40	212
rect	40	211	41	212
rect	41	211	42	212
rect	43	211	44	212
rect	44	211	45	212
rect	45	211	46	212
rect	46	211	47	212
rect	48	211	49	212
rect	49	211	50	212
rect	50	211	51	212
rect	68	211	69	212
rect	69	211	70	212
rect	70	211	71	212
rect	71	211	72	212
rect	72	211	73	212
rect	73	211	74	212
rect	74	211	75	212
rect	129	211	130	212
rect	130	211	131	212
rect	131	211	132	212
rect	132	211	133	212
rect	133	211	134	212
rect	134	211	135	212
rect	139	211	140	212
rect	148	211	149	212
rect	149	211	150	212
rect	151	211	152	212
rect	175	211	176	212
rect	176	211	177	212
rect	177	211	178	212
rect	178	211	179	212
rect	179	211	180	212
rect	234	211	235	212
rect	235	211	236	212
rect	236	211	237	212
rect	237	211	238	212
rect	238	211	239	212
rect	239	211	240	212
rect	240	211	241	212
rect	241	211	242	212
rect	242	211	243	212
rect	243	211	244	212
rect	244	211	245	212
rect	245	211	246	212
rect	255	211	256	212
rect	256	211	257	212
rect	257	211	258	212
rect	259	211	260	212
rect	260	211	261	212
rect	262	211	263	212
rect	263	211	264	212
rect	265	211	266	212
rect	266	211	267	212
rect	268	211	269	212
rect	269	211	270	212
rect	270	211	271	212
rect	271	211	272	212
rect	272	211	273	212
rect	274	211	275	212
rect	275	211	276	212
rect	276	211	277	212
rect	277	211	278	212
rect	279	211	280	212
rect	280	211	281	212
rect	281	211	282	212
rect	282	211	283	212
rect	283	211	284	212
rect	284	211	285	212
rect	286	211	287	212
rect	287	211	288	212
rect	288	211	289	212
rect	289	211	290	212
rect	290	211	291	212
rect	291	211	292	212
rect	292	211	293	212
rect	293	211	294	212
rect	294	211	295	212
rect	295	211	296	212
rect	297	211	298	212
rect	298	211	299	212
rect	299	211	300	212
rect	300	211	301	212
rect	302	211	303	212
rect	303	211	304	212
rect	305	211	306	212
rect	306	211	307	212
rect	308	211	309	212
rect	309	211	310	212
rect	311	211	312	212
rect	312	211	313	212
rect	313	211	314	212
rect	314	211	315	212
rect	315	211	316	212
rect	317	211	318	212
rect	318	211	319	212
rect	320	211	321	212
rect	321	211	322	212
rect	323	211	324	212
rect	324	211	325	212
rect	326	211	327	212
rect	327	211	328	212
rect	329	211	330	212
rect	330	211	331	212
rect	332	211	333	212
rect	333	211	334	212
rect	334	211	335	212
rect	335	211	336	212
rect	336	211	337	212
rect	337	211	338	212
rect	369	211	370	212
rect	370	211	371	212
rect	371	211	372	212
rect	372	211	373	212
rect	373	211	374	212
rect	374	211	375	212
rect	375	211	376	212
rect	376	211	377	212
rect	377	211	378	212
rect	378	211	379	212
rect	379	211	380	212
rect	380	211	381	212
rect	381	211	382	212
rect	382	211	383	212
rect	383	211	384	212
rect	384	211	385	212
rect	386	211	387	212
rect	387	211	388	212
rect	388	211	389	212
rect	389	211	390	212
rect	390	211	391	212
rect	9	213	10	214
rect	10	213	11	214
rect	11	213	12	214
rect	12	213	13	214
rect	13	213	14	214
rect	14	213	15	214
rect	15	213	16	214
rect	16	213	17	214
rect	18	213	19	214
rect	19	213	20	214
rect	20	213	21	214
rect	21	213	22	214
rect	22	213	23	214
rect	23	213	24	214
rect	25	213	26	214
rect	27	213	28	214
rect	28	213	29	214
rect	29	213	30	214
rect	30	213	31	214
rect	31	213	32	214
rect	32	213	33	214
rect	33	213	34	214
rect	34	213	35	214
rect	35	213	36	214
rect	36	213	37	214
rect	37	213	38	214
rect	39	213	40	214
rect	40	213	41	214
rect	41	213	42	214
rect	43	213	44	214
rect	44	213	45	214
rect	45	213	46	214
rect	46	213	47	214
rect	48	213	49	214
rect	49	213	50	214
rect	50	213	51	214
rect	51	213	52	214
rect	52	213	53	214
rect	54	213	55	214
rect	55	213	56	214
rect	57	213	58	214
rect	58	213	59	214
rect	59	213	60	214
rect	60	213	61	214
rect	62	213	63	214
rect	63	213	64	214
rect	64	213	65	214
rect	65	213	66	214
rect	66	213	67	214
rect	67	213	68	214
rect	68	213	69	214
rect	69	213	70	214
rect	70	213	71	214
rect	71	213	72	214
rect	72	213	73	214
rect	73	213	74	214
rect	74	213	75	214
rect	76	213	77	214
rect	77	213	78	214
rect	78	213	79	214
rect	79	213	80	214
rect	80	213	81	214
rect	81	213	82	214
rect	82	213	83	214
rect	83	213	84	214
rect	84	213	85	214
rect	85	213	86	214
rect	86	213	87	214
rect	87	213	88	214
rect	88	213	89	214
rect	89	213	90	214
rect	90	213	91	214
rect	91	213	92	214
rect	92	213	93	214
rect	93	213	94	214
rect	94	213	95	214
rect	95	213	96	214
rect	96	213	97	214
rect	97	213	98	214
rect	99	213	100	214
rect	100	213	101	214
rect	102	213	103	214
rect	103	213	104	214
rect	104	213	105	214
rect	105	213	106	214
rect	106	213	107	214
rect	107	213	108	214
rect	108	213	109	214
rect	109	213	110	214
rect	110	213	111	214
rect	111	213	112	214
rect	112	213	113	214
rect	113	213	114	214
rect	114	213	115	214
rect	115	213	116	214
rect	116	213	117	214
rect	118	213	119	214
rect	119	213	120	214
rect	120	213	121	214
rect	121	213	122	214
rect	122	213	123	214
rect	123	213	124	214
rect	124	213	125	214
rect	125	213	126	214
rect	127	213	128	214
rect	128	213	129	214
rect	129	213	130	214
rect	130	213	131	214
rect	131	213	132	214
rect	132	213	133	214
rect	133	213	134	214
rect	134	213	135	214
rect	136	213	137	214
rect	137	213	138	214
rect	139	213	140	214
rect	140	213	141	214
rect	141	213	142	214
rect	142	213	143	214
rect	143	213	144	214
rect	144	213	145	214
rect	145	213	146	214
rect	146	213	147	214
rect	148	213	149	214
rect	149	213	150	214
rect	151	213	152	214
rect	152	213	153	214
rect	153	213	154	214
rect	154	213	155	214
rect	155	213	156	214
rect	156	213	157	214
rect	157	213	158	214
rect	158	213	159	214
rect	160	213	161	214
rect	161	213	162	214
rect	162	213	163	214
rect	163	213	164	214
rect	164	213	165	214
rect	165	213	166	214
rect	166	213	167	214
rect	167	213	168	214
rect	169	213	170	214
rect	170	213	171	214
rect	172	213	173	214
rect	173	213	174	214
rect	174	213	175	214
rect	175	213	176	214
rect	176	213	177	214
rect	177	213	178	214
rect	178	213	179	214
rect	179	213	180	214
rect	181	213	182	214
rect	182	213	183	214
rect	183	213	184	214
rect	184	213	185	214
rect	185	213	186	214
rect	187	213	188	214
rect	188	213	189	214
rect	189	213	190	214
rect	190	213	191	214
rect	191	213	192	214
rect	192	213	193	214
rect	193	213	194	214
rect	194	213	195	214
rect	195	213	196	214
rect	196	213	197	214
rect	197	213	198	214
rect	198	213	199	214
rect	199	213	200	214
rect	200	213	201	214
rect	201	213	202	214
rect	203	213	204	214
rect	204	213	205	214
rect	205	213	206	214
rect	207	213	208	214
rect	209	213	210	214
rect	210	213	211	214
rect	211	213	212	214
rect	213	213	214	214
rect	214	213	215	214
rect	216	213	217	214
rect	217	213	218	214
rect	218	213	219	214
rect	219	213	220	214
rect	220	213	221	214
rect	221	213	222	214
rect	222	213	223	214
rect	223	213	224	214
rect	225	213	226	214
rect	226	213	227	214
rect	227	213	228	214
rect	228	213	229	214
rect	229	213	230	214
rect	231	213	232	214
rect	232	213	233	214
rect	233	213	234	214
rect	234	213	235	214
rect	235	213	236	214
rect	236	213	237	214
rect	237	213	238	214
rect	238	213	239	214
rect	239	213	240	214
rect	240	213	241	214
rect	241	213	242	214
rect	242	213	243	214
rect	243	213	244	214
rect	244	213	245	214
rect	245	213	246	214
rect	247	213	248	214
rect	248	213	249	214
rect	250	213	251	214
rect	252	213	253	214
rect	253	213	254	214
rect	254	213	255	214
rect	255	213	256	214
rect	256	213	257	214
rect	257	213	258	214
rect	259	213	260	214
rect	260	213	261	214
rect	262	213	263	214
rect	263	213	264	214
rect	265	213	266	214
rect	266	213	267	214
rect	268	213	269	214
rect	269	213	270	214
rect	270	213	271	214
rect	271	213	272	214
rect	272	213	273	214
rect	274	213	275	214
rect	275	213	276	214
rect	276	213	277	214
rect	277	213	278	214
rect	279	213	280	214
rect	280	213	281	214
rect	281	213	282	214
rect	282	213	283	214
rect	283	213	284	214
rect	284	213	285	214
rect	286	213	287	214
rect	287	213	288	214
rect	288	213	289	214
rect	289	213	290	214
rect	290	213	291	214
rect	291	213	292	214
rect	292	213	293	214
rect	293	213	294	214
rect	294	213	295	214
rect	295	213	296	214
rect	297	213	298	214
rect	298	213	299	214
rect	299	213	300	214
rect	300	213	301	214
rect	302	213	303	214
rect	303	213	304	214
rect	305	213	306	214
rect	306	213	307	214
rect	308	213	309	214
rect	309	213	310	214
rect	311	213	312	214
rect	312	213	313	214
rect	313	213	314	214
rect	314	213	315	214
rect	315	213	316	214
rect	317	213	318	214
rect	318	213	319	214
rect	320	213	321	214
rect	321	213	322	214
rect	323	213	324	214
rect	324	213	325	214
rect	326	213	327	214
rect	327	213	328	214
rect	329	213	330	214
rect	330	213	331	214
rect	332	213	333	214
rect	333	213	334	214
rect	334	213	335	214
rect	335	213	336	214
rect	336	213	337	214
rect	337	213	338	214
rect	338	213	339	214
rect	339	213	340	214
rect	341	213	342	214
rect	342	213	343	214
rect	344	213	345	214
rect	345	213	346	214
rect	346	213	347	214
rect	347	213	348	214
rect	348	213	349	214
rect	349	213	350	214
rect	350	213	351	214
rect	351	213	352	214
rect	360	213	361	214
rect	361	213	362	214
rect	362	213	363	214
rect	363	213	364	214
rect	364	213	365	214
rect	365	213	366	214
rect	366	213	367	214
rect	367	213	368	214
rect	369	213	370	214
rect	370	213	371	214
rect	388	213	389	214
rect	389	213	390	214
rect	390	213	391	214
rect	391	213	392	214
rect	392	213	393	214
rect	393	213	394	214
rect	9	215	10	216
rect	10	215	11	216
rect	11	215	12	216
rect	12	215	13	216
rect	13	215	14	216
rect	25	215	26	216
rect	27	215	28	216
rect	28	215	29	216
rect	29	215	30	216
rect	30	215	31	216
rect	31	215	32	216
rect	32	215	33	216
rect	33	215	34	216
rect	34	215	35	216
rect	43	215	44	216
rect	44	215	45	216
rect	45	215	46	216
rect	46	215	47	216
rect	48	215	49	216
rect	49	215	50	216
rect	62	215	63	216
rect	63	215	64	216
rect	64	215	65	216
rect	65	215	66	216
rect	66	215	67	216
rect	67	215	68	216
rect	68	215	69	216
rect	69	215	70	216
rect	70	215	71	216
rect	71	215	72	216
rect	82	215	83	216
rect	83	215	84	216
rect	84	215	85	216
rect	85	215	86	216
rect	86	215	87	216
rect	87	215	88	216
rect	88	215	89	216
rect	89	215	90	216
rect	90	215	91	216
rect	91	215	92	216
rect	92	215	93	216
rect	93	215	94	216
rect	94	215	95	216
rect	95	215	96	216
rect	96	215	97	216
rect	97	215	98	216
rect	99	215	100	216
rect	100	215	101	216
rect	102	215	103	216
rect	103	215	104	216
rect	104	215	105	216
rect	105	215	106	216
rect	106	215	107	216
rect	107	215	108	216
rect	108	215	109	216
rect	109	215	110	216
rect	110	215	111	216
rect	111	215	112	216
rect	112	215	113	216
rect	113	215	114	216
rect	114	215	115	216
rect	115	215	116	216
rect	116	215	117	216
rect	118	215	119	216
rect	119	215	120	216
rect	120	215	121	216
rect	121	215	122	216
rect	122	215	123	216
rect	123	215	124	216
rect	124	215	125	216
rect	125	215	126	216
rect	127	215	128	216
rect	128	215	129	216
rect	129	215	130	216
rect	130	215	131	216
rect	131	215	132	216
rect	132	215	133	216
rect	133	215	134	216
rect	134	215	135	216
rect	136	215	137	216
rect	137	215	138	216
rect	139	215	140	216
rect	140	215	141	216
rect	141	215	142	216
rect	142	215	143	216
rect	143	215	144	216
rect	144	215	145	216
rect	145	215	146	216
rect	146	215	147	216
rect	148	215	149	216
rect	149	215	150	216
rect	151	215	152	216
rect	152	215	153	216
rect	153	215	154	216
rect	154	215	155	216
rect	155	215	156	216
rect	156	215	157	216
rect	157	215	158	216
rect	158	215	159	216
rect	160	215	161	216
rect	161	215	162	216
rect	172	215	173	216
rect	173	215	174	216
rect	174	215	175	216
rect	175	215	176	216
rect	176	215	177	216
rect	209	215	210	216
rect	210	215	211	216
rect	211	215	212	216
rect	213	215	214	216
rect	214	215	215	216
rect	216	215	217	216
rect	217	215	218	216
rect	218	215	219	216
rect	219	215	220	216
rect	220	215	221	216
rect	221	215	222	216
rect	222	215	223	216
rect	223	215	224	216
rect	225	215	226	216
rect	226	215	227	216
rect	231	215	232	216
rect	232	215	233	216
rect	233	215	234	216
rect	234	215	235	216
rect	235	215	236	216
rect	236	215	237	216
rect	237	215	238	216
rect	238	215	239	216
rect	239	215	240	216
rect	240	215	241	216
rect	241	215	242	216
rect	242	215	243	216
rect	252	215	253	216
rect	253	215	254	216
rect	254	215	255	216
rect	255	215	256	216
rect	256	215	257	216
rect	257	215	258	216
rect	259	215	260	216
rect	260	215	261	216
rect	262	215	263	216
rect	263	215	264	216
rect	265	215	266	216
rect	266	215	267	216
rect	268	215	269	216
rect	269	215	270	216
rect	279	215	280	216
rect	280	215	281	216
rect	281	215	282	216
rect	297	215	298	216
rect	298	215	299	216
rect	299	215	300	216
rect	300	215	301	216
rect	302	215	303	216
rect	303	215	304	216
rect	305	215	306	216
rect	306	215	307	216
rect	308	215	309	216
rect	309	215	310	216
rect	311	215	312	216
rect	312	215	313	216
rect	313	215	314	216
rect	314	215	315	216
rect	315	215	316	216
rect	317	215	318	216
rect	318	215	319	216
rect	320	215	321	216
rect	321	215	322	216
rect	323	215	324	216
rect	324	215	325	216
rect	326	215	327	216
rect	327	215	328	216
rect	329	215	330	216
rect	330	215	331	216
rect	332	215	333	216
rect	333	215	334	216
rect	334	215	335	216
rect	335	215	336	216
rect	336	215	337	216
rect	337	215	338	216
rect	338	215	339	216
rect	339	215	340	216
rect	341	215	342	216
rect	342	215	343	216
rect	344	215	345	216
rect	345	215	346	216
rect	346	215	347	216
rect	347	215	348	216
rect	348	215	349	216
rect	349	215	350	216
rect	350	215	351	216
rect	351	215	352	216
rect	353	215	354	216
rect	354	215	355	216
rect	355	215	356	216
rect	356	215	357	216
rect	357	215	358	216
rect	358	215	359	216
rect	359	215	360	216
rect	360	215	361	216
rect	361	215	362	216
rect	362	215	363	216
rect	363	215	364	216
rect	364	215	365	216
rect	365	215	366	216
rect	366	215	367	216
rect	367	215	368	216
rect	369	215	370	216
rect	370	215	371	216
rect	372	215	373	216
rect	373	215	374	216
rect	374	215	375	216
rect	375	215	376	216
rect	376	215	377	216
rect	377	215	378	216
rect	378	215	379	216
rect	379	215	380	216
rect	380	215	381	216
rect	381	215	382	216
rect	382	215	383	216
rect	383	215	384	216
rect	384	215	385	216
rect	241	224	242	225
rect	242	224	243	225
rect	244	224	245	225
rect	245	224	246	225
rect	247	224	248	225
rect	248	224	249	225
rect	250	224	251	225
rect	251	224	252	225
rect	253	224	254	225
rect	254	224	255	225
rect	255	224	256	225
rect	256	224	257	225
rect	257	224	258	225
rect	259	224	260	225
rect	260	224	261	225
rect	262	224	263	225
rect	263	224	264	225
rect	265	224	266	225
rect	266	224	267	225
rect	262	226	263	227
rect	263	226	264	227
rect	265	226	266	227
rect	181	228	182	229
rect	182	228	183	229
rect	183	228	184	229
rect	184	228	185	229
rect	185	228	186	229
rect	186	228	187	229
rect	187	228	188	229
rect	250	228	251	229
rect	251	228	252	229
rect	259	228	260	229
rect	260	228	261	229
rect	261	228	262	229
rect	262	228	263	229
rect	263	228	264	229
rect	265	228	266	229
rect	267	228	268	229
rect	268	228	269	229
rect	269	228	270	229
rect	271	228	272	229
rect	272	228	273	229
rect	274	228	275	229
rect	275	228	276	229
rect	151	230	152	231
rect	152	230	153	231
rect	153	230	154	231
rect	154	230	155	231
rect	155	230	156	231
rect	156	230	157	231
rect	157	230	158	231
rect	158	230	159	231
rect	160	230	161	231
rect	178	230	179	231
rect	179	230	180	231
rect	180	230	181	231
rect	181	230	182	231
rect	182	230	183	231
rect	183	230	184	231
rect	184	230	185	231
rect	222	230	223	231
rect	223	230	224	231
rect	249	230	250	231
rect	250	230	251	231
rect	251	230	252	231
rect	252	230	253	231
rect	253	230	254	231
rect	254	230	255	231
rect	255	230	256	231
rect	256	230	257	231
rect	257	230	258	231
rect	258	230	259	231
rect	259	230	260	231
rect	274	230	275	231
rect	57	232	58	233
rect	58	232	59	233
rect	59	232	60	233
rect	136	232	137	233
rect	138	232	139	233
rect	139	232	140	233
rect	140	232	141	233
rect	141	232	142	233
rect	142	232	143	233
rect	143	232	144	233
rect	144	232	145	233
rect	145	232	146	233
rect	146	232	147	233
rect	148	232	149	233
rect	171	232	172	233
rect	172	232	173	233
rect	173	232	174	233
rect	174	232	175	233
rect	175	232	176	233
rect	176	232	177	233
rect	177	232	178	233
rect	178	232	179	233
rect	204	232	205	233
rect	205	232	206	233
rect	207	232	208	233
rect	208	232	209	233
rect	209	232	210	233
rect	216	232	217	233
rect	217	232	218	233
rect	218	232	219	233
rect	219	232	220	233
rect	220	232	221	233
rect	221	232	222	233
rect	222	232	223	233
rect	223	232	224	233
rect	224	232	225	233
rect	225	232	226	233
rect	226	232	227	233
rect	228	232	229	233
rect	229	232	230	233
rect	230	232	231	233
rect	231	232	232	233
rect	247	232	248	233
rect	249	232	250	233
rect	250	232	251	233
rect	251	232	252	233
rect	252	232	253	233
rect	253	232	254	233
rect	254	232	255	233
rect	255	232	256	233
rect	256	232	257	233
rect	257	232	258	233
rect	258	232	259	233
rect	259	232	260	233
rect	261	232	262	233
rect	262	232	263	233
rect	263	232	264	233
rect	265	232	266	233
rect	267	232	268	233
rect	268	232	269	233
rect	269	232	270	233
rect	271	232	272	233
rect	54	234	55	235
rect	55	234	56	235
rect	56	234	57	235
rect	102	234	103	235
rect	103	234	104	235
rect	104	234	105	235
rect	105	234	106	235
rect	135	234	136	235
rect	136	234	137	235
rect	138	234	139	235
rect	139	234	140	235
rect	140	234	141	235
rect	141	234	142	235
rect	142	234	143	235
rect	143	234	144	235
rect	144	234	145	235
rect	145	234	146	235
rect	146	234	147	235
rect	169	234	170	235
rect	171	234	172	235
rect	172	234	173	235
rect	173	234	174	235
rect	174	234	175	235
rect	175	234	176	235
rect	198	234	199	235
rect	199	234	200	235
rect	200	234	201	235
rect	201	234	202	235
rect	202	234	203	235
rect	203	234	204	235
rect	204	234	205	235
rect	205	234	206	235
rect	215	234	216	235
rect	216	234	217	235
rect	217	234	218	235
rect	218	234	219	235
rect	219	234	220	235
rect	244	234	245	235
rect	245	234	246	235
rect	246	234	247	235
rect	247	234	248	235
rect	249	234	250	235
rect	250	234	251	235
rect	326	234	327	235
rect	327	234	328	235
rect	329	234	330	235
rect	330	234	331	235
rect	332	234	333	235
rect	333	234	334	235
rect	335	234	336	235
rect	51	236	52	237
rect	52	236	53	237
rect	53	236	54	237
rect	99	236	100	237
rect	100	236	101	237
rect	101	236	102	237
rect	102	236	103	237
rect	103	236	104	237
rect	104	236	105	237
rect	105	236	106	237
rect	107	236	108	237
rect	108	236	109	237
rect	127	236	128	237
rect	128	236	129	237
rect	129	236	130	237
rect	130	236	131	237
rect	131	236	132	237
rect	132	236	133	237
rect	133	236	134	237
rect	135	236	136	237
rect	136	236	137	237
rect	138	236	139	237
rect	139	236	140	237
rect	160	236	161	237
rect	162	236	163	237
rect	163	236	164	237
rect	164	236	165	237
rect	166	236	167	237
rect	167	236	168	237
rect	168	236	169	237
rect	169	236	170	237
rect	171	236	172	237
rect	172	236	173	237
rect	194	236	195	237
rect	195	236	196	237
rect	196	236	197	237
rect	198	236	199	237
rect	199	236	200	237
rect	200	236	201	237
rect	201	236	202	237
rect	202	236	203	237
rect	203	236	204	237
rect	204	236	205	237
rect	205	236	206	237
rect	206	236	207	237
rect	207	236	208	237
rect	208	236	209	237
rect	209	236	210	237
rect	211	236	212	237
rect	212	236	213	237
rect	213	236	214	237
rect	215	236	216	237
rect	216	236	217	237
rect	217	236	218	237
rect	218	236	219	237
rect	219	236	220	237
rect	221	236	222	237
rect	222	236	223	237
rect	223	236	224	237
rect	224	236	225	237
rect	225	236	226	237
rect	226	236	227	237
rect	228	236	229	237
rect	229	236	230	237
rect	230	236	231	237
rect	231	236	232	237
rect	233	236	234	237
rect	234	236	235	237
rect	235	236	236	237
rect	236	236	237	237
rect	237	236	238	237
rect	238	236	239	237
rect	239	236	240	237
rect	240	236	241	237
rect	241	236	242	237
rect	242	236	243	237
rect	243	236	244	237
rect	244	236	245	237
rect	245	236	246	237
rect	246	236	247	237
rect	247	236	248	237
rect	249	236	250	237
rect	250	236	251	237
rect	252	236	253	237
rect	253	236	254	237
rect	254	236	255	237
rect	255	236	256	237
rect	256	236	257	237
rect	257	236	258	237
rect	258	236	259	237
rect	259	236	260	237
rect	261	236	262	237
rect	262	236	263	237
rect	263	236	264	237
rect	265	236	266	237
rect	267	236	268	237
rect	268	236	269	237
rect	269	236	270	237
rect	271	236	272	237
rect	273	236	274	237
rect	274	236	275	237
rect	276	236	277	237
rect	277	236	278	237
rect	278	236	279	237
rect	279	236	280	237
rect	280	236	281	237
rect	281	236	282	237
rect	283	236	284	237
rect	284	236	285	237
rect	320	236	321	237
rect	321	236	322	237
rect	323	236	324	237
rect	324	236	325	237
rect	325	236	326	237
rect	326	236	327	237
rect	327	236	328	237
rect	329	236	330	237
rect	330	236	331	237
rect	332	236	333	237
rect	333	236	334	237
rect	341	236	342	237
rect	342	236	343	237
rect	344	236	345	237
rect	345	236	346	237
rect	48	238	49	239
rect	49	238	50	239
rect	50	238	51	239
rect	81	238	82	239
rect	82	238	83	239
rect	83	238	84	239
rect	84	238	85	239
rect	85	238	86	239
rect	86	238	87	239
rect	87	238	88	239
rect	88	238	89	239
rect	89	238	90	239
rect	90	238	91	239
rect	91	238	92	239
rect	93	238	94	239
rect	94	238	95	239
rect	95	238	96	239
rect	96	238	97	239
rect	97	238	98	239
rect	98	238	99	239
rect	99	238	100	239
rect	100	238	101	239
rect	101	238	102	239
rect	102	238	103	239
rect	103	238	104	239
rect	104	238	105	239
rect	105	238	106	239
rect	107	238	108	239
rect	108	238	109	239
rect	110	238	111	239
rect	111	238	112	239
rect	112	238	113	239
rect	113	238	114	239
rect	114	238	115	239
rect	115	238	116	239
rect	116	238	117	239
rect	117	238	118	239
rect	119	238	120	239
rect	120	238	121	239
rect	121	238	122	239
rect	122	238	123	239
rect	123	238	124	239
rect	124	238	125	239
rect	125	238	126	239
rect	126	238	127	239
rect	127	238	128	239
rect	128	238	129	239
rect	129	238	130	239
rect	130	238	131	239
rect	131	238	132	239
rect	132	238	133	239
rect	133	238	134	239
rect	135	238	136	239
rect	136	238	137	239
rect	138	238	139	239
rect	139	238	140	239
rect	141	238	142	239
rect	142	238	143	239
rect	143	238	144	239
rect	144	238	145	239
rect	145	238	146	239
rect	146	238	147	239
rect	147	238	148	239
rect	148	238	149	239
rect	150	238	151	239
rect	151	238	152	239
rect	152	238	153	239
rect	153	238	154	239
rect	154	238	155	239
rect	155	238	156	239
rect	156	238	157	239
rect	157	238	158	239
rect	166	238	167	239
rect	167	238	168	239
rect	168	238	169	239
rect	169	238	170	239
rect	171	238	172	239
rect	172	238	173	239
rect	174	238	175	239
rect	175	238	176	239
rect	177	238	178	239
rect	178	238	179	239
rect	180	238	181	239
rect	181	238	182	239
rect	182	238	183	239
rect	183	238	184	239
rect	184	238	185	239
rect	186	238	187	239
rect	187	238	188	239
rect	189	238	190	239
rect	190	238	191	239
rect	191	238	192	239
rect	192	238	193	239
rect	193	238	194	239
rect	194	238	195	239
rect	195	238	196	239
rect	196	238	197	239
rect	198	238	199	239
rect	199	238	200	239
rect	200	238	201	239
rect	201	238	202	239
rect	202	238	203	239
rect	203	238	204	239
rect	204	238	205	239
rect	205	238	206	239
rect	206	238	207	239
rect	207	238	208	239
rect	208	238	209	239
rect	209	238	210	239
rect	211	238	212	239
rect	212	238	213	239
rect	213	238	214	239
rect	215	238	216	239
rect	216	238	217	239
rect	217	238	218	239
rect	218	238	219	239
rect	219	238	220	239
rect	221	238	222	239
rect	222	238	223	239
rect	223	238	224	239
rect	224	238	225	239
rect	225	238	226	239
rect	226	238	227	239
rect	228	238	229	239
rect	229	238	230	239
rect	230	238	231	239
rect	231	238	232	239
rect	233	238	234	239
rect	234	238	235	239
rect	235	238	236	239
rect	236	238	237	239
rect	237	238	238	239
rect	238	238	239	239
rect	239	238	240	239
rect	240	238	241	239
rect	241	238	242	239
rect	242	238	243	239
rect	243	238	244	239
rect	244	238	245	239
rect	245	238	246	239
rect	246	238	247	239
rect	247	238	248	239
rect	249	238	250	239
rect	250	238	251	239
rect	252	238	253	239
rect	253	238	254	239
rect	254	238	255	239
rect	255	238	256	239
rect	256	238	257	239
rect	257	238	258	239
rect	258	238	259	239
rect	259	238	260	239
rect	261	238	262	239
rect	262	238	263	239
rect	263	238	264	239
rect	265	238	266	239
rect	267	238	268	239
rect	268	238	269	239
rect	269	238	270	239
rect	271	238	272	239
rect	273	238	274	239
rect	274	238	275	239
rect	276	238	277	239
rect	277	238	278	239
rect	278	238	279	239
rect	279	238	280	239
rect	280	238	281	239
rect	281	238	282	239
rect	283	238	284	239
rect	284	238	285	239
rect	285	238	286	239
rect	286	238	287	239
rect	287	238	288	239
rect	288	238	289	239
rect	289	238	290	239
rect	290	238	291	239
rect	291	238	292	239
rect	292	238	293	239
rect	293	238	294	239
rect	294	238	295	239
rect	295	238	296	239
rect	296	238	297	239
rect	297	238	298	239
rect	298	238	299	239
rect	299	238	300	239
rect	300	238	301	239
rect	302	238	303	239
rect	303	238	304	239
rect	305	238	306	239
rect	306	238	307	239
rect	308	238	309	239
rect	309	238	310	239
rect	311	238	312	239
rect	312	238	313	239
rect	313	238	314	239
rect	314	238	315	239
rect	315	238	316	239
rect	317	238	318	239
rect	318	238	319	239
rect	319	238	320	239
rect	320	238	321	239
rect	321	238	322	239
rect	323	238	324	239
rect	329	238	330	239
rect	330	238	331	239
rect	332	238	333	239
rect	333	238	334	239
rect	334	238	335	239
rect	335	238	336	239
rect	337	238	338	239
rect	338	238	339	239
rect	25	240	26	241
rect	36	240	37	241
rect	37	240	38	241
rect	39	240	40	241
rect	40	240	41	241
rect	41	240	42	241
rect	42	240	43	241
rect	43	240	44	241
rect	44	240	45	241
rect	45	240	46	241
rect	46	240	47	241
rect	47	240	48	241
rect	76	240	77	241
rect	77	240	78	241
rect	78	240	79	241
rect	79	240	80	241
rect	81	240	82	241
rect	82	240	83	241
rect	83	240	84	241
rect	84	240	85	241
rect	85	240	86	241
rect	86	240	87	241
rect	87	240	88	241
rect	88	240	89	241
rect	89	240	90	241
rect	90	240	91	241
rect	91	240	92	241
rect	93	240	94	241
rect	94	240	95	241
rect	95	240	96	241
rect	96	240	97	241
rect	97	240	98	241
rect	98	240	99	241
rect	99	240	100	241
rect	100	240	101	241
rect	101	240	102	241
rect	102	240	103	241
rect	103	240	104	241
rect	104	240	105	241
rect	105	240	106	241
rect	107	240	108	241
rect	108	240	109	241
rect	110	240	111	241
rect	111	240	112	241
rect	112	240	113	241
rect	113	240	114	241
rect	114	240	115	241
rect	115	240	116	241
rect	116	240	117	241
rect	117	240	118	241
rect	119	240	120	241
rect	120	240	121	241
rect	121	240	122	241
rect	122	240	123	241
rect	123	240	124	241
rect	124	240	125	241
rect	125	240	126	241
rect	126	240	127	241
rect	127	240	128	241
rect	128	240	129	241
rect	129	240	130	241
rect	130	240	131	241
rect	131	240	132	241
rect	132	240	133	241
rect	133	240	134	241
rect	135	240	136	241
rect	136	240	137	241
rect	138	240	139	241
rect	139	240	140	241
rect	141	240	142	241
rect	142	240	143	241
rect	143	240	144	241
rect	144	240	145	241
rect	145	240	146	241
rect	146	240	147	241
rect	147	240	148	241
rect	148	240	149	241
rect	150	240	151	241
rect	151	240	152	241
rect	152	240	153	241
rect	153	240	154	241
rect	154	240	155	241
rect	155	240	156	241
rect	156	240	157	241
rect	157	240	158	241
rect	159	240	160	241
rect	160	240	161	241
rect	162	240	163	241
rect	163	240	164	241
rect	164	240	165	241
rect	165	240	166	241
rect	166	240	167	241
rect	167	240	168	241
rect	168	240	169	241
rect	169	240	170	241
rect	171	240	172	241
rect	172	240	173	241
rect	174	240	175	241
rect	175	240	176	241
rect	177	240	178	241
rect	178	240	179	241
rect	180	240	181	241
rect	181	240	182	241
rect	182	240	183	241
rect	183	240	184	241
rect	184	240	185	241
rect	186	240	187	241
rect	187	240	188	241
rect	189	240	190	241
rect	190	240	191	241
rect	191	240	192	241
rect	192	240	193	241
rect	193	240	194	241
rect	194	240	195	241
rect	195	240	196	241
rect	196	240	197	241
rect	198	240	199	241
rect	199	240	200	241
rect	200	240	201	241
rect	201	240	202	241
rect	202	240	203	241
rect	203	240	204	241
rect	204	240	205	241
rect	205	240	206	241
rect	206	240	207	241
rect	207	240	208	241
rect	208	240	209	241
rect	209	240	210	241
rect	211	240	212	241
rect	212	240	213	241
rect	213	240	214	241
rect	215	240	216	241
rect	216	240	217	241
rect	217	240	218	241
rect	218	240	219	241
rect	219	240	220	241
rect	221	240	222	241
rect	222	240	223	241
rect	223	240	224	241
rect	224	240	225	241
rect	225	240	226	241
rect	226	240	227	241
rect	228	240	229	241
rect	229	240	230	241
rect	230	240	231	241
rect	231	240	232	241
rect	233	240	234	241
rect	234	240	235	241
rect	235	240	236	241
rect	236	240	237	241
rect	237	240	238	241
rect	238	240	239	241
rect	239	240	240	241
rect	240	240	241	241
rect	241	240	242	241
rect	242	240	243	241
rect	243	240	244	241
rect	244	240	245	241
rect	245	240	246	241
rect	246	240	247	241
rect	247	240	248	241
rect	249	240	250	241
rect	250	240	251	241
rect	252	240	253	241
rect	253	240	254	241
rect	254	240	255	241
rect	255	240	256	241
rect	256	240	257	241
rect	257	240	258	241
rect	258	240	259	241
rect	259	240	260	241
rect	261	240	262	241
rect	262	240	263	241
rect	263	240	264	241
rect	265	240	266	241
rect	267	240	268	241
rect	268	240	269	241
rect	269	240	270	241
rect	271	240	272	241
rect	273	240	274	241
rect	274	240	275	241
rect	276	240	277	241
rect	277	240	278	241
rect	278	240	279	241
rect	279	240	280	241
rect	280	240	281	241
rect	281	240	282	241
rect	283	240	284	241
rect	284	240	285	241
rect	285	240	286	241
rect	286	240	287	241
rect	287	240	288	241
rect	288	240	289	241
rect	289	240	290	241
rect	290	240	291	241
rect	291	240	292	241
rect	292	240	293	241
rect	293	240	294	241
rect	294	240	295	241
rect	295	240	296	241
rect	296	240	297	241
rect	297	240	298	241
rect	298	240	299	241
rect	299	240	300	241
rect	300	240	301	241
rect	302	240	303	241
rect	303	240	304	241
rect	305	240	306	241
rect	306	240	307	241
rect	308	240	309	241
rect	309	240	310	241
rect	311	240	312	241
rect	312	240	313	241
rect	313	240	314	241
rect	314	240	315	241
rect	315	240	316	241
rect	317	240	318	241
rect	318	240	319	241
rect	319	240	320	241
rect	320	240	321	241
rect	321	240	322	241
rect	323	240	324	241
rect	325	240	326	241
rect	326	240	327	241
rect	332	240	333	241
rect	333	240	334	241
rect	334	240	335	241
rect	335	240	336	241
rect	337	240	338	241
rect	338	240	339	241
rect	340	240	341	241
rect	341	240	342	241
rect	342	240	343	241
rect	344	240	345	241
rect	345	240	346	241
rect	346	240	347	241
rect	347	240	348	241
rect	348	240	349	241
rect	350	240	351	241
rect	351	240	352	241
rect	353	240	354	241
rect	354	240	355	241
rect	355	240	356	241
rect	356	240	357	241
rect	357	240	358	241
rect	358	240	359	241
rect	359	240	360	241
rect	360	240	361	241
rect	361	240	362	241
rect	18	242	19	243
rect	19	242	20	243
rect	20	242	21	243
rect	21	242	22	243
rect	22	242	23	243
rect	23	242	24	243
rect	25	242	26	243
rect	26	242	27	243
rect	31	242	32	243
rect	32	242	33	243
rect	33	242	34	243
rect	34	242	35	243
rect	35	242	36	243
rect	36	242	37	243
rect	37	242	38	243
rect	73	242	74	243
rect	74	242	75	243
rect	75	242	76	243
rect	76	242	77	243
rect	77	242	78	243
rect	78	242	79	243
rect	79	242	80	243
rect	81	242	82	243
rect	82	242	83	243
rect	93	242	94	243
rect	94	242	95	243
rect	95	242	96	243
rect	96	242	97	243
rect	97	242	98	243
rect	98	242	99	243
rect	99	242	100	243
rect	100	242	101	243
rect	101	242	102	243
rect	102	242	103	243
rect	103	242	104	243
rect	104	242	105	243
rect	105	242	106	243
rect	107	242	108	243
rect	108	242	109	243
rect	110	242	111	243
rect	111	242	112	243
rect	112	242	113	243
rect	113	242	114	243
rect	114	242	115	243
rect	115	242	116	243
rect	116	242	117	243
rect	117	242	118	243
rect	119	242	120	243
rect	120	242	121	243
rect	121	242	122	243
rect	122	242	123	243
rect	123	242	124	243
rect	124	242	125	243
rect	125	242	126	243
rect	126	242	127	243
rect	127	242	128	243
rect	128	242	129	243
rect	129	242	130	243
rect	130	242	131	243
rect	131	242	132	243
rect	132	242	133	243
rect	133	242	134	243
rect	135	242	136	243
rect	136	242	137	243
rect	138	242	139	243
rect	139	242	140	243
rect	141	242	142	243
rect	142	242	143	243
rect	143	242	144	243
rect	144	242	145	243
rect	145	242	146	243
rect	146	242	147	243
rect	147	242	148	243
rect	148	242	149	243
rect	150	242	151	243
rect	151	242	152	243
rect	152	242	153	243
rect	153	242	154	243
rect	154	242	155	243
rect	155	242	156	243
rect	156	242	157	243
rect	157	242	158	243
rect	159	242	160	243
rect	160	242	161	243
rect	162	242	163	243
rect	163	242	164	243
rect	164	242	165	243
rect	165	242	166	243
rect	166	242	167	243
rect	167	242	168	243
rect	168	242	169	243
rect	169	242	170	243
rect	171	242	172	243
rect	172	242	173	243
rect	174	242	175	243
rect	175	242	176	243
rect	177	242	178	243
rect	178	242	179	243
rect	180	242	181	243
rect	181	242	182	243
rect	182	242	183	243
rect	183	242	184	243
rect	184	242	185	243
rect	186	242	187	243
rect	187	242	188	243
rect	189	242	190	243
rect	190	242	191	243
rect	191	242	192	243
rect	192	242	193	243
rect	193	242	194	243
rect	194	242	195	243
rect	195	242	196	243
rect	196	242	197	243
rect	198	242	199	243
rect	199	242	200	243
rect	200	242	201	243
rect	201	242	202	243
rect	202	242	203	243
rect	203	242	204	243
rect	204	242	205	243
rect	205	242	206	243
rect	206	242	207	243
rect	207	242	208	243
rect	208	242	209	243
rect	209	242	210	243
rect	211	242	212	243
rect	212	242	213	243
rect	213	242	214	243
rect	215	242	216	243
rect	216	242	217	243
rect	217	242	218	243
rect	218	242	219	243
rect	219	242	220	243
rect	221	242	222	243
rect	222	242	223	243
rect	223	242	224	243
rect	224	242	225	243
rect	225	242	226	243
rect	226	242	227	243
rect	228	242	229	243
rect	229	242	230	243
rect	230	242	231	243
rect	231	242	232	243
rect	233	242	234	243
rect	234	242	235	243
rect	235	242	236	243
rect	236	242	237	243
rect	237	242	238	243
rect	238	242	239	243
rect	239	242	240	243
rect	240	242	241	243
rect	241	242	242	243
rect	242	242	243	243
rect	243	242	244	243
rect	244	242	245	243
rect	245	242	246	243
rect	246	242	247	243
rect	247	242	248	243
rect	249	242	250	243
rect	250	242	251	243
rect	252	242	253	243
rect	253	242	254	243
rect	254	242	255	243
rect	255	242	256	243
rect	256	242	257	243
rect	257	242	258	243
rect	258	242	259	243
rect	259	242	260	243
rect	261	242	262	243
rect	262	242	263	243
rect	263	242	264	243
rect	265	242	266	243
rect	267	242	268	243
rect	268	242	269	243
rect	269	242	270	243
rect	271	242	272	243
rect	273	242	274	243
rect	274	242	275	243
rect	276	242	277	243
rect	277	242	278	243
rect	278	242	279	243
rect	279	242	280	243
rect	280	242	281	243
rect	281	242	282	243
rect	283	242	284	243
rect	284	242	285	243
rect	285	242	286	243
rect	286	242	287	243
rect	287	242	288	243
rect	288	242	289	243
rect	289	242	290	243
rect	290	242	291	243
rect	291	242	292	243
rect	292	242	293	243
rect	293	242	294	243
rect	294	242	295	243
rect	295	242	296	243
rect	296	242	297	243
rect	297	242	298	243
rect	298	242	299	243
rect	299	242	300	243
rect	300	242	301	243
rect	302	242	303	243
rect	303	242	304	243
rect	305	242	306	243
rect	306	242	307	243
rect	308	242	309	243
rect	309	242	310	243
rect	311	242	312	243
rect	312	242	313	243
rect	313	242	314	243
rect	314	242	315	243
rect	315	242	316	243
rect	317	242	318	243
rect	318	242	319	243
rect	319	242	320	243
rect	320	242	321	243
rect	321	242	322	243
rect	323	242	324	243
rect	325	242	326	243
rect	326	242	327	243
rect	328	242	329	243
rect	329	242	330	243
rect	330	242	331	243
rect	331	242	332	243
rect	332	242	333	243
rect	344	242	345	243
rect	345	242	346	243
rect	346	242	347	243
rect	347	242	348	243
rect	348	242	349	243
rect	361	242	362	243
rect	362	242	363	243
rect	363	242	364	243
rect	364	242	365	243
rect	365	242	366	243
rect	366	242	367	243
rect	367	242	368	243
rect	372	242	373	243
rect	373	242	374	243
rect	374	242	375	243
rect	375	242	376	243
rect	15	244	16	245
rect	16	244	17	245
rect	17	244	18	245
rect	18	244	19	245
rect	19	244	20	245
rect	20	244	21	245
rect	37	244	38	245
rect	38	244	39	245
rect	67	244	68	245
rect	68	244	69	245
rect	69	244	70	245
rect	70	244	71	245
rect	71	244	72	245
rect	72	244	73	245
rect	73	244	74	245
rect	74	244	75	245
rect	75	244	76	245
rect	76	244	77	245
rect	77	244	78	245
rect	78	244	79	245
rect	79	244	80	245
rect	81	244	82	245
rect	82	244	83	245
rect	84	244	85	245
rect	85	244	86	245
rect	86	244	87	245
rect	87	244	88	245
rect	88	244	89	245
rect	89	244	90	245
rect	90	244	91	245
rect	91	244	92	245
rect	92	244	93	245
rect	93	244	94	245
rect	94	244	95	245
rect	95	244	96	245
rect	96	244	97	245
rect	97	244	98	245
rect	98	244	99	245
rect	99	244	100	245
rect	100	244	101	245
rect	101	244	102	245
rect	102	244	103	245
rect	103	244	104	245
rect	104	244	105	245
rect	105	244	106	245
rect	107	244	108	245
rect	108	244	109	245
rect	110	244	111	245
rect	111	244	112	245
rect	112	244	113	245
rect	113	244	114	245
rect	114	244	115	245
rect	115	244	116	245
rect	116	244	117	245
rect	117	244	118	245
rect	119	244	120	245
rect	120	244	121	245
rect	121	244	122	245
rect	122	244	123	245
rect	123	244	124	245
rect	124	244	125	245
rect	125	244	126	245
rect	126	244	127	245
rect	127	244	128	245
rect	128	244	129	245
rect	129	244	130	245
rect	130	244	131	245
rect	131	244	132	245
rect	132	244	133	245
rect	133	244	134	245
rect	135	244	136	245
rect	136	244	137	245
rect	138	244	139	245
rect	139	244	140	245
rect	141	244	142	245
rect	142	244	143	245
rect	143	244	144	245
rect	144	244	145	245
rect	145	244	146	245
rect	146	244	147	245
rect	147	244	148	245
rect	148	244	149	245
rect	150	244	151	245
rect	151	244	152	245
rect	152	244	153	245
rect	153	244	154	245
rect	154	244	155	245
rect	155	244	156	245
rect	156	244	157	245
rect	157	244	158	245
rect	159	244	160	245
rect	160	244	161	245
rect	162	244	163	245
rect	163	244	164	245
rect	164	244	165	245
rect	165	244	166	245
rect	166	244	167	245
rect	167	244	168	245
rect	168	244	169	245
rect	169	244	170	245
rect	171	244	172	245
rect	172	244	173	245
rect	174	244	175	245
rect	175	244	176	245
rect	177	244	178	245
rect	178	244	179	245
rect	180	244	181	245
rect	181	244	182	245
rect	182	244	183	245
rect	183	244	184	245
rect	184	244	185	245
rect	186	244	187	245
rect	187	244	188	245
rect	189	244	190	245
rect	190	244	191	245
rect	191	244	192	245
rect	192	244	193	245
rect	193	244	194	245
rect	194	244	195	245
rect	195	244	196	245
rect	196	244	197	245
rect	198	244	199	245
rect	199	244	200	245
rect	200	244	201	245
rect	201	244	202	245
rect	202	244	203	245
rect	203	244	204	245
rect	204	244	205	245
rect	205	244	206	245
rect	206	244	207	245
rect	207	244	208	245
rect	208	244	209	245
rect	209	244	210	245
rect	211	244	212	245
rect	212	244	213	245
rect	213	244	214	245
rect	215	244	216	245
rect	216	244	217	245
rect	217	244	218	245
rect	218	244	219	245
rect	219	244	220	245
rect	221	244	222	245
rect	222	244	223	245
rect	228	244	229	245
rect	229	244	230	245
rect	230	244	231	245
rect	231	244	232	245
rect	233	244	234	245
rect	234	244	235	245
rect	235	244	236	245
rect	236	244	237	245
rect	237	244	238	245
rect	238	244	239	245
rect	239	244	240	245
rect	240	244	241	245
rect	241	244	242	245
rect	242	244	243	245
rect	243	244	244	245
rect	244	244	245	245
rect	245	244	246	245
rect	246	244	247	245
rect	247	244	248	245
rect	249	244	250	245
rect	250	244	251	245
rect	252	244	253	245
rect	253	244	254	245
rect	271	244	272	245
rect	273	244	274	245
rect	274	244	275	245
rect	276	244	277	245
rect	277	244	278	245
rect	278	244	279	245
rect	279	244	280	245
rect	280	244	281	245
rect	281	244	282	245
rect	283	244	284	245
rect	284	244	285	245
rect	285	244	286	245
rect	286	244	287	245
rect	317	244	318	245
rect	318	244	319	245
rect	319	244	320	245
rect	320	244	321	245
rect	321	244	322	245
rect	323	244	324	245
rect	325	244	326	245
rect	326	244	327	245
rect	328	244	329	245
rect	329	244	330	245
rect	330	244	331	245
rect	331	244	332	245
rect	332	244	333	245
rect	334	244	335	245
rect	335	244	336	245
rect	337	244	338	245
rect	338	244	339	245
rect	340	244	341	245
rect	341	244	342	245
rect	342	244	343	245
rect	343	244	344	245
rect	344	244	345	245
rect	345	244	346	245
rect	346	244	347	245
rect	347	244	348	245
rect	348	244	349	245
rect	349	244	350	245
rect	350	244	351	245
rect	351	244	352	245
rect	353	244	354	245
rect	354	244	355	245
rect	355	244	356	245
rect	356	244	357	245
rect	357	244	358	245
rect	358	244	359	245
rect	359	244	360	245
rect	361	244	362	245
rect	362	244	363	245
rect	363	244	364	245
rect	364	244	365	245
rect	365	244	366	245
rect	366	244	367	245
rect	367	244	368	245
rect	368	244	369	245
rect	369	244	370	245
rect	370	244	371	245
rect	371	244	372	245
rect	372	244	373	245
rect	373	244	374	245
rect	374	244	375	245
rect	375	244	376	245
rect	377	244	378	245
rect	378	244	379	245
rect	379	244	380	245
rect	380	244	381	245
rect	5	246	6	247
rect	6	246	7	247
rect	7	246	8	247
rect	8	246	9	247
rect	9	246	10	247
rect	10	246	11	247
rect	11	246	12	247
rect	12	246	13	247
rect	13	246	14	247
rect	14	246	15	247
rect	15	246	16	247
rect	16	246	17	247
rect	17	246	18	247
rect	18	246	19	247
rect	19	246	20	247
rect	20	246	21	247
rect	22	246	23	247
rect	23	246	24	247
rect	25	246	26	247
rect	26	246	27	247
rect	28	246	29	247
rect	29	246	30	247
rect	31	246	32	247
rect	32	246	33	247
rect	33	246	34	247
rect	34	246	35	247
rect	35	246	36	247
rect	37	246	38	247
rect	38	246	39	247
rect	40	246	41	247
rect	41	246	42	247
rect	42	246	43	247
rect	43	246	44	247
rect	44	246	45	247
rect	45	246	46	247
rect	46	246	47	247
rect	47	246	48	247
rect	49	246	50	247
rect	50	246	51	247
rect	52	246	53	247
rect	53	246	54	247
rect	55	246	56	247
rect	56	246	57	247
rect	58	246	59	247
rect	59	246	60	247
rect	61	246	62	247
rect	62	246	63	247
rect	63	246	64	247
rect	64	246	65	247
rect	65	246	66	247
rect	66	246	67	247
rect	67	246	68	247
rect	68	246	69	247
rect	69	246	70	247
rect	70	246	71	247
rect	71	246	72	247
rect	72	246	73	247
rect	73	246	74	247
rect	74	246	75	247
rect	75	246	76	247
rect	76	246	77	247
rect	77	246	78	247
rect	78	246	79	247
rect	79	246	80	247
rect	81	246	82	247
rect	82	246	83	247
rect	84	246	85	247
rect	85	246	86	247
rect	86	246	87	247
rect	87	246	88	247
rect	88	246	89	247
rect	89	246	90	247
rect	90	246	91	247
rect	91	246	92	247
rect	92	246	93	247
rect	93	246	94	247
rect	94	246	95	247
rect	95	246	96	247
rect	96	246	97	247
rect	97	246	98	247
rect	98	246	99	247
rect	99	246	100	247
rect	100	246	101	247
rect	101	246	102	247
rect	102	246	103	247
rect	103	246	104	247
rect	104	246	105	247
rect	105	246	106	247
rect	107	246	108	247
rect	108	246	109	247
rect	110	246	111	247
rect	111	246	112	247
rect	112	246	113	247
rect	113	246	114	247
rect	114	246	115	247
rect	115	246	116	247
rect	116	246	117	247
rect	117	246	118	247
rect	119	246	120	247
rect	120	246	121	247
rect	121	246	122	247
rect	122	246	123	247
rect	123	246	124	247
rect	124	246	125	247
rect	125	246	126	247
rect	126	246	127	247
rect	127	246	128	247
rect	128	246	129	247
rect	129	246	130	247
rect	130	246	131	247
rect	131	246	132	247
rect	132	246	133	247
rect	133	246	134	247
rect	135	246	136	247
rect	136	246	137	247
rect	138	246	139	247
rect	139	246	140	247
rect	141	246	142	247
rect	142	246	143	247
rect	143	246	144	247
rect	144	246	145	247
rect	145	246	146	247
rect	146	246	147	247
rect	147	246	148	247
rect	148	246	149	247
rect	150	246	151	247
rect	151	246	152	247
rect	152	246	153	247
rect	153	246	154	247
rect	154	246	155	247
rect	155	246	156	247
rect	156	246	157	247
rect	157	246	158	247
rect	159	246	160	247
rect	160	246	161	247
rect	162	246	163	247
rect	163	246	164	247
rect	164	246	165	247
rect	165	246	166	247
rect	166	246	167	247
rect	167	246	168	247
rect	168	246	169	247
rect	169	246	170	247
rect	171	246	172	247
rect	172	246	173	247
rect	174	246	175	247
rect	175	246	176	247
rect	177	246	178	247
rect	178	246	179	247
rect	180	246	181	247
rect	181	246	182	247
rect	182	246	183	247
rect	183	246	184	247
rect	184	246	185	247
rect	186	246	187	247
rect	187	246	188	247
rect	189	246	190	247
rect	190	246	191	247
rect	191	246	192	247
rect	192	246	193	247
rect	193	246	194	247
rect	194	246	195	247
rect	195	246	196	247
rect	196	246	197	247
rect	198	246	199	247
rect	199	246	200	247
rect	200	246	201	247
rect	201	246	202	247
rect	202	246	203	247
rect	203	246	204	247
rect	204	246	205	247
rect	205	246	206	247
rect	206	246	207	247
rect	207	246	208	247
rect	208	246	209	247
rect	209	246	210	247
rect	211	246	212	247
rect	212	246	213	247
rect	213	246	214	247
rect	215	246	216	247
rect	216	246	217	247
rect	217	246	218	247
rect	218	246	219	247
rect	219	246	220	247
rect	221	246	222	247
rect	222	246	223	247
rect	224	246	225	247
rect	225	246	226	247
rect	226	246	227	247
rect	227	246	228	247
rect	228	246	229	247
rect	229	246	230	247
rect	230	246	231	247
rect	231	246	232	247
rect	233	246	234	247
rect	234	246	235	247
rect	235	246	236	247
rect	236	246	237	247
rect	237	246	238	247
rect	238	246	239	247
rect	239	246	240	247
rect	240	246	241	247
rect	241	246	242	247
rect	242	246	243	247
rect	243	246	244	247
rect	244	246	245	247
rect	245	246	246	247
rect	246	246	247	247
rect	247	246	248	247
rect	249	246	250	247
rect	250	246	251	247
rect	252	246	253	247
rect	253	246	254	247
rect	255	246	256	247
rect	256	246	257	247
rect	265	246	266	247
rect	267	246	268	247
rect	268	246	269	247
rect	283	246	284	247
rect	297	246	298	247
rect	298	246	299	247
rect	299	246	300	247
rect	300	246	301	247
rect	311	246	312	247
rect	312	246	313	247
rect	313	246	314	247
rect	314	246	315	247
rect	315	246	316	247
rect	316	246	317	247
rect	317	246	318	247
rect	318	246	319	247
rect	319	246	320	247
rect	320	246	321	247
rect	321	246	322	247
rect	349	246	350	247
rect	350	246	351	247
rect	351	246	352	247
rect	358	246	359	247
rect	359	246	360	247
rect	361	246	362	247
rect	362	246	363	247
rect	371	246	372	247
rect	372	246	373	247
rect	380	246	381	247
rect	381	246	382	247
rect	382	246	383	247
rect	383	246	384	247
rect	384	246	385	247
rect	385	246	386	247
rect	386	246	387	247
rect	282	255	283	256
rect	283	255	284	256
rect	285	255	286	256
rect	286	255	287	256
rect	288	255	289	256
rect	289	255	290	256
rect	290	255	291	256
rect	291	255	292	256
rect	292	255	293	256
rect	293	255	294	256
rect	294	255	295	256
rect	295	255	296	256
rect	297	255	298	256
rect	298	255	299	256
rect	299	255	300	256
rect	300	255	301	256
rect	301	255	302	256
rect	302	255	303	256
rect	303	255	304	256
rect	304	255	305	256
rect	306	255	307	256
rect	307	255	308	256
rect	309	255	310	256
rect	310	255	311	256
rect	311	255	312	256
rect	312	255	313	256
rect	313	255	314	256
rect	315	255	316	256
rect	316	255	317	256
rect	317	255	318	256
rect	318	255	319	256
rect	319	255	320	256
rect	320	255	321	256
rect	321	255	322	256
rect	322	255	323	256
rect	323	255	324	256
rect	325	255	326	256
rect	326	255	327	256
rect	327	255	328	256
rect	328	255	329	256
rect	329	255	330	256
rect	330	255	331	256
rect	331	255	332	256
rect	332	255	333	256
rect	334	255	335	256
rect	335	255	336	256
rect	337	255	338	256
rect	338	255	339	256
rect	340	255	341	256
rect	341	255	342	256
rect	342	255	343	256
rect	343	255	344	256
rect	344	255	345	256
rect	345	255	346	256
rect	346	255	347	256
rect	347	255	348	256
rect	349	255	350	256
rect	350	255	351	256
rect	351	255	352	256
rect	352	255	353	256
rect	353	255	354	256
rect	354	255	355	256
rect	355	255	356	256
rect	356	255	357	256
rect	358	255	359	256
rect	359	255	360	256
rect	360	255	361	256
rect	361	255	362	256
rect	362	255	363	256
rect	363	255	364	256
rect	364	255	365	256
rect	365	255	366	256
rect	180	257	181	258
rect	181	257	182	258
rect	182	257	183	258
rect	183	257	184	258
rect	184	257	185	258
rect	276	257	277	258
rect	277	257	278	258
rect	278	257	279	258
rect	279	257	280	258
rect	58	259	59	260
rect	59	259	60	260
rect	61	259	62	260
rect	62	259	63	260
rect	159	259	160	260
rect	160	259	161	260
rect	162	259	163	260
rect	163	259	164	260
rect	174	259	175	260
rect	175	259	176	260
rect	177	259	178	260
rect	178	259	179	260
rect	179	259	180	260
rect	180	259	181	260
rect	181	259	182	260
rect	182	259	183	260
rect	183	259	184	260
rect	184	259	185	260
rect	185	259	186	260
rect	186	259	187	260
rect	187	259	188	260
rect	189	259	190	260
rect	190	259	191	260
rect	191	259	192	260
rect	192	259	193	260
rect	193	259	194	260
rect	195	259	196	260
rect	196	259	197	260
rect	198	259	199	260
rect	199	259	200	260
rect	258	259	259	260
rect	259	259	260	260
rect	260	259	261	260
rect	261	259	262	260
rect	267	259	268	260
rect	268	259	269	260
rect	270	259	271	260
rect	271	259	272	260
rect	273	259	274	260
rect	274	259	275	260
rect	275	259	276	260
rect	276	259	277	260
rect	277	259	278	260
rect	278	259	279	260
rect	279	259	280	260
rect	281	259	282	260
rect	282	259	283	260
rect	283	259	284	260
rect	285	259	286	260
rect	286	259	287	260
rect	288	259	289	260
rect	380	259	381	260
rect	22	261	23	262
rect	23	261	24	262
rect	25	261	26	262
rect	26	261	27	262
rect	28	261	29	262
rect	29	261	30	262
rect	31	261	32	262
rect	32	261	33	262
rect	55	261	56	262
rect	56	261	57	262
rect	141	261	142	262
rect	142	261	143	262
rect	143	261	144	262
rect	144	261	145	262
rect	145	261	146	262
rect	146	261	147	262
rect	147	261	148	262
rect	148	261	149	262
rect	150	261	151	262
rect	164	261	165	262
rect	165	261	166	262
rect	166	261	167	262
rect	167	261	168	262
rect	168	261	169	262
rect	169	261	170	262
rect	171	261	172	262
rect	177	261	178	262
rect	178	261	179	262
rect	179	261	180	262
rect	180	261	181	262
rect	181	261	182	262
rect	182	261	183	262
rect	183	261	184	262
rect	184	261	185	262
rect	255	261	256	262
rect	256	261	257	262
rect	257	261	258	262
rect	258	261	259	262
rect	259	261	260	262
rect	260	261	261	262
rect	261	261	262	262
rect	263	261	264	262
rect	264	261	265	262
rect	273	261	274	262
rect	274	261	275	262
rect	275	261	276	262
rect	276	261	277	262
rect	285	261	286	262
rect	286	261	287	262
rect	288	261	289	262
rect	290	261	291	262
rect	291	261	292	262
rect	292	261	293	262
rect	293	261	294	262
rect	294	261	295	262
rect	295	261	296	262
rect	297	261	298	262
rect	334	261	335	262
rect	335	261	336	262
rect	337	261	338	262
rect	338	261	339	262
rect	340	261	341	262
rect	358	261	359	262
rect	359	261	360	262
rect	360	261	361	262
rect	361	261	362	262
rect	362	261	363	262
rect	363	261	364	262
rect	364	261	365	262
rect	365	261	366	262
rect	367	261	368	262
rect	368	261	369	262
rect	369	261	370	262
rect	370	261	371	262
rect	371	261	372	262
rect	372	261	373	262
rect	374	261	375	262
rect	375	261	376	262
rect	377	261	378	262
rect	22	263	23	264
rect	23	263	24	264
rect	28	263	29	264
rect	29	263	30	264
rect	31	263	32	264
rect	32	263	33	264
rect	34	263	35	264
rect	35	263	36	264
rect	52	263	53	264
rect	53	263	54	264
rect	61	263	62	264
rect	62	263	63	264
rect	64	263	65	264
rect	65	263	66	264
rect	113	263	114	264
rect	114	263	115	264
rect	115	263	116	264
rect	116	263	117	264
rect	117	263	118	264
rect	119	263	120	264
rect	120	263	121	264
rect	121	263	122	264
rect	122	263	123	264
rect	123	263	124	264
rect	135	263	136	264
rect	136	263	137	264
rect	138	263	139	264
rect	162	263	163	264
rect	164	263	165	264
rect	165	263	166	264
rect	166	263	167	264
rect	167	263	168	264
rect	168	263	169	264
rect	169	263	170	264
rect	171	263	172	264
rect	173	263	174	264
rect	174	263	175	264
rect	195	263	196	264
rect	196	263	197	264
rect	198	263	199	264
rect	199	263	200	264
rect	201	263	202	264
rect	202	263	203	264
rect	203	263	204	264
rect	204	263	205	264
rect	205	263	206	264
rect	206	263	207	264
rect	207	263	208	264
rect	208	263	209	264
rect	209	263	210	264
rect	210	263	211	264
rect	211	263	212	264
rect	212	263	213	264
rect	213	263	214	264
rect	214	263	215	264
rect	215	263	216	264
rect	216	263	217	264
rect	217	263	218	264
rect	218	263	219	264
rect	219	263	220	264
rect	221	263	222	264
rect	222	263	223	264
rect	224	263	225	264
rect	225	263	226	264
rect	226	263	227	264
rect	227	263	228	264
rect	228	263	229	264
rect	229	263	230	264
rect	230	263	231	264
rect	231	263	232	264
rect	233	263	234	264
rect	234	263	235	264
rect	235	263	236	264
rect	236	263	237	264
rect	237	263	238	264
rect	238	263	239	264
rect	239	263	240	264
rect	240	263	241	264
rect	241	263	242	264
rect	242	263	243	264
rect	243	263	244	264
rect	244	263	245	264
rect	245	263	246	264
rect	246	263	247	264
rect	247	263	248	264
rect	249	263	250	264
rect	250	263	251	264
rect	252	263	253	264
rect	253	263	254	264
rect	254	263	255	264
rect	255	263	256	264
rect	256	263	257	264
rect	257	263	258	264
rect	258	263	259	264
rect	259	263	260	264
rect	260	263	261	264
rect	261	263	262	264
rect	263	263	264	264
rect	264	263	265	264
rect	266	263	267	264
rect	267	263	268	264
rect	268	263	269	264
rect	270	263	271	264
rect	271	263	272	264
rect	272	263	273	264
rect	273	263	274	264
rect	274	263	275	264
rect	275	263	276	264
rect	276	263	277	264
rect	278	263	279	264
rect	279	263	280	264
rect	281	263	282	264
rect	282	263	283	264
rect	283	263	284	264
rect	284	263	285	264
rect	285	263	286	264
rect	286	263	287	264
rect	288	263	289	264
rect	290	263	291	264
rect	291	263	292	264
rect	292	263	293	264
rect	293	263	294	264
rect	294	263	295	264
rect	295	263	296	264
rect	297	263	298	264
rect	299	263	300	264
rect	300	263	301	264
rect	301	263	302	264
rect	302	263	303	264
rect	303	263	304	264
rect	304	263	305	264
rect	306	263	307	264
rect	307	263	308	264
rect	309	263	310	264
rect	310	263	311	264
rect	311	263	312	264
rect	312	263	313	264
rect	313	263	314	264
rect	315	263	316	264
rect	316	263	317	264
rect	317	263	318	264
rect	318	263	319	264
rect	319	263	320	264
rect	327	263	328	264
rect	328	263	329	264
rect	329	263	330	264
rect	330	263	331	264
rect	331	263	332	264
rect	332	263	333	264
rect	333	263	334	264
rect	334	263	335	264
rect	335	263	336	264
rect	340	263	341	264
rect	342	263	343	264
rect	343	263	344	264
rect	349	263	350	264
rect	350	263	351	264
rect	351	263	352	264
rect	352	263	353	264
rect	353	263	354	264
rect	354	263	355	264
rect	355	263	356	264
rect	356	263	357	264
rect	357	263	358	264
rect	358	263	359	264
rect	359	263	360	264
rect	25	265	26	266
rect	26	265	27	266
rect	27	265	28	266
rect	28	265	29	266
rect	29	265	30	266
rect	40	265	41	266
rect	41	265	42	266
rect	42	265	43	266
rect	43	265	44	266
rect	44	265	45	266
rect	49	265	50	266
rect	50	265	51	266
rect	51	265	52	266
rect	52	265	53	266
rect	53	265	54	266
rect	55	265	56	266
rect	56	265	57	266
rect	58	265	59	266
rect	59	265	60	266
rect	60	265	61	266
rect	61	265	62	266
rect	62	265	63	266
rect	64	265	65	266
rect	65	265	66	266
rect	67	265	68	266
rect	68	265	69	266
rect	69	265	70	266
rect	70	265	71	266
rect	71	265	72	266
rect	72	265	73	266
rect	73	265	74	266
rect	74	265	75	266
rect	90	265	91	266
rect	104	265	105	266
rect	105	265	106	266
rect	107	265	108	266
rect	108	265	109	266
rect	110	265	111	266
rect	111	265	112	266
rect	134	265	135	266
rect	135	265	136	266
rect	136	265	137	266
rect	138	265	139	266
rect	140	265	141	266
rect	141	265	142	266
rect	161	265	162	266
rect	162	265	163	266
rect	164	265	165	266
rect	165	265	166	266
rect	166	265	167	266
rect	167	265	168	266
rect	168	265	169	266
rect	169	265	170	266
rect	192	265	193	266
rect	193	265	194	266
rect	194	265	195	266
rect	195	265	196	266
rect	196	265	197	266
rect	224	265	225	266
rect	225	265	226	266
rect	226	265	227	266
rect	252	265	253	266
rect	253	265	254	266
rect	254	265	255	266
rect	255	265	256	266
rect	256	265	257	266
rect	257	265	258	266
rect	258	265	259	266
rect	259	265	260	266
rect	260	265	261	266
rect	261	265	262	266
rect	263	265	264	266
rect	264	265	265	266
rect	266	265	267	266
rect	267	265	268	266
rect	268	265	269	266
rect	270	265	271	266
rect	271	265	272	266
rect	272	265	273	266
rect	273	265	274	266
rect	284	265	285	266
rect	285	265	286	266
rect	286	265	287	266
rect	315	265	316	266
rect	316	265	317	266
rect	317	265	318	266
rect	318	265	319	266
rect	319	265	320	266
rect	321	265	322	266
rect	322	265	323	266
rect	323	265	324	266
rect	325	265	326	266
rect	327	265	328	266
rect	328	265	329	266
rect	329	265	330	266
rect	330	265	331	266
rect	331	265	332	266
rect	332	265	333	266
rect	333	265	334	266
rect	334	265	335	266
rect	335	265	336	266
rect	336	265	337	266
rect	337	265	338	266
rect	338	265	339	266
rect	339	265	340	266
rect	340	265	341	266
rect	342	265	343	266
rect	343	265	344	266
rect	345	265	346	266
rect	346	265	347	266
rect	347	265	348	266
rect	348	265	349	266
rect	349	265	350	266
rect	350	265	351	266
rect	351	265	352	266
rect	352	265	353	266
rect	353	265	354	266
rect	354	265	355	266
rect	355	265	356	266
rect	356	265	357	266
rect	357	265	358	266
rect	358	265	359	266
rect	359	265	360	266
rect	361	265	362	266
rect	362	265	363	266
rect	374	265	375	266
rect	375	265	376	266
rect	377	265	378	266
rect	379	265	380	266
rect	380	265	381	266
rect	382	265	383	266
rect	383	265	384	266
rect	384	265	385	266
rect	385	265	386	266
rect	386	265	387	266
rect	5	267	6	268
rect	6	267	7	268
rect	7	267	8	268
rect	8	267	9	268
rect	9	267	10	268
rect	10	267	11	268
rect	11	267	12	268
rect	12	267	13	268
rect	13	267	14	268
rect	14	267	15	268
rect	15	267	16	268
rect	16	267	17	268
rect	17	267	18	268
rect	18	267	19	268
rect	19	267	20	268
rect	20	267	21	268
rect	22	267	23	268
rect	23	267	24	268
rect	25	267	26	268
rect	26	267	27	268
rect	27	267	28	268
rect	28	267	29	268
rect	29	267	30	268
rect	30	267	31	268
rect	31	267	32	268
rect	32	267	33	268
rect	34	267	35	268
rect	35	267	36	268
rect	37	267	38	268
rect	38	267	39	268
rect	39	267	40	268
rect	40	267	41	268
rect	41	267	42	268
rect	42	267	43	268
rect	43	267	44	268
rect	44	267	45	268
rect	46	267	47	268
rect	47	267	48	268
rect	48	267	49	268
rect	49	267	50	268
rect	50	267	51	268
rect	51	267	52	268
rect	52	267	53	268
rect	53	267	54	268
rect	55	267	56	268
rect	56	267	57	268
rect	58	267	59	268
rect	59	267	60	268
rect	84	267	85	268
rect	85	267	86	268
rect	86	267	87	268
rect	87	267	88	268
rect	88	267	89	268
rect	89	267	90	268
rect	90	267	91	268
rect	92	267	93	268
rect	93	267	94	268
rect	94	267	95	268
rect	95	267	96	268
rect	96	267	97	268
rect	97	267	98	268
rect	98	267	99	268
rect	99	267	100	268
rect	104	267	105	268
rect	105	267	106	268
rect	110	267	111	268
rect	111	267	112	268
rect	113	267	114	268
rect	114	267	115	268
rect	119	267	120	268
rect	120	267	121	268
rect	121	267	122	268
rect	122	267	123	268
rect	123	267	124	268
rect	125	267	126	268
rect	126	267	127	268
rect	131	267	132	268
rect	132	267	133	268
rect	134	267	135	268
rect	135	267	136	268
rect	136	267	137	268
rect	150	267	151	268
rect	152	267	153	268
rect	153	267	154	268
rect	154	267	155	268
rect	155	267	156	268
rect	156	267	157	268
rect	157	267	158	268
rect	158	267	159	268
rect	159	267	160	268
rect	161	267	162	268
rect	162	267	163	268
rect	164	267	165	268
rect	165	267	166	268
rect	166	267	167	268
rect	167	267	168	268
rect	168	267	169	268
rect	189	267	190	268
rect	190	267	191	268
rect	192	267	193	268
rect	193	267	194	268
rect	221	267	222	268
rect	222	267	223	268
rect	223	267	224	268
rect	233	267	234	268
rect	234	267	235	268
rect	235	267	236	268
rect	249	267	250	268
rect	250	267	251	268
rect	251	267	252	268
rect	252	267	253	268
rect	253	267	254	268
rect	254	267	255	268
rect	255	267	256	268
rect	256	267	257	268
rect	257	267	258	268
rect	258	267	259	268
rect	270	267	271	268
rect	271	267	272	268
rect	272	267	273	268
rect	273	267	274	268
rect	275	267	276	268
rect	276	267	277	268
rect	278	267	279	268
rect	279	267	280	268
rect	281	267	282	268
rect	282	267	283	268
rect	284	267	285	268
rect	285	267	286	268
rect	286	267	287	268
rect	287	267	288	268
rect	288	267	289	268
rect	290	267	291	268
rect	291	267	292	268
rect	297	267	298	268
rect	299	267	300	268
rect	300	267	301	268
rect	301	267	302	268
rect	306	267	307	268
rect	307	267	308	268
rect	309	267	310	268
rect	310	267	311	268
rect	311	267	312	268
rect	312	267	313	268
rect	313	267	314	268
rect	314	267	315	268
rect	315	267	316	268
rect	316	267	317	268
rect	330	267	331	268
rect	331	267	332	268
rect	332	267	333	268
rect	333	267	334	268
rect	334	267	335	268
rect	339	267	340	268
rect	340	267	341	268
rect	342	267	343	268
rect	343	267	344	268
rect	345	267	346	268
rect	346	267	347	268
rect	347	267	348	268
rect	348	267	349	268
rect	349	267	350	268
rect	350	267	351	268
rect	351	267	352	268
rect	352	267	353	268
rect	353	267	354	268
rect	354	267	355	268
rect	355	267	356	268
rect	356	267	357	268
rect	370	267	371	268
rect	371	267	372	268
rect	372	267	373	268
rect	373	267	374	268
rect	374	267	375	268
rect	375	267	376	268
rect	293	276	294	277
rect	294	276	295	277
rect	295	276	296	277
rect	296	276	297	277
rect	297	276	298	277
rect	298	276	299	277
rect	299	276	300	277
rect	300	276	301	277
rect	301	276	302	277
rect	302	276	303	277
rect	303	276	304	277
rect	304	276	305	277
rect	305	276	306	277
rect	306	276	307	277
rect	307	276	308	277
rect	309	276	310	277
rect	310	276	311	277
rect	382	276	383	277
rect	383	276	384	277
rect	384	276	385	277
rect	385	276	386	277
rect	386	276	387	277
rect	290	278	291	279
rect	291	278	292	279
rect	292	278	293	279
rect	293	278	294	279
rect	294	278	295	279
rect	295	278	296	279
rect	296	278	297	279
rect	297	278	298	279
rect	298	278	299	279
rect	299	278	300	279
rect	300	278	301	279
rect	301	278	302	279
rect	302	278	303	279
rect	303	278	304	279
rect	304	278	305	279
rect	305	278	306	279
rect	306	278	307	279
rect	307	278	308	279
rect	339	278	340	279
rect	340	278	341	279
rect	342	278	343	279
rect	343	278	344	279
rect	345	278	346	279
rect	346	278	347	279
rect	347	278	348	279
rect	348	278	349	279
rect	349	278	350	279
rect	351	278	352	279
rect	352	278	353	279
rect	353	278	354	279
rect	354	278	355	279
rect	355	278	356	279
rect	356	278	357	279
rect	361	278	362	279
rect	362	278	363	279
rect	364	278	365	279
rect	365	278	366	279
rect	367	278	368	279
rect	368	278	369	279
rect	370	278	371	279
rect	371	278	372	279
rect	373	278	374	279
rect	374	278	375	279
rect	375	278	376	279
rect	376	278	377	279
rect	377	278	378	279
rect	379	278	380	279
rect	380	278	381	279
rect	189	280	190	281
rect	190	280	191	281
rect	275	280	276	281
rect	276	280	277	281
rect	278	280	279	281
rect	279	280	280	281
rect	281	280	282	281
rect	282	280	283	281
rect	284	280	285	281
rect	285	280	286	281
rect	286	280	287	281
rect	287	280	288	281
rect	288	280	289	281
rect	290	280	291	281
rect	291	280	292	281
rect	292	280	293	281
rect	293	280	294	281
rect	294	280	295	281
rect	295	280	296	281
rect	296	280	297	281
rect	297	280	298	281
rect	298	280	299	281
rect	299	280	300	281
rect	300	280	301	281
rect	301	280	302	281
rect	302	280	303	281
rect	303	280	304	281
rect	304	280	305	281
rect	305	280	306	281
rect	306	280	307	281
rect	307	280	308	281
rect	336	280	337	281
rect	337	280	338	281
rect	338	280	339	281
rect	339	280	340	281
rect	340	280	341	281
rect	342	280	343	281
rect	343	280	344	281
rect	345	280	346	281
rect	346	280	347	281
rect	347	280	348	281
rect	348	280	349	281
rect	349	280	350	281
rect	351	280	352	281
rect	352	280	353	281
rect	353	280	354	281
rect	354	280	355	281
rect	355	280	356	281
rect	356	280	357	281
rect	358	280	359	281
rect	359	280	360	281
rect	64	282	65	283
rect	65	282	66	283
rect	67	282	68	283
rect	68	282	69	283
rect	108	282	109	283
rect	109	282	110	283
rect	110	282	111	283
rect	111	282	112	283
rect	113	282	114	283
rect	114	282	115	283
rect	131	282	132	283
rect	132	282	133	283
rect	146	282	147	283
rect	147	282	148	283
rect	148	282	149	283
rect	149	282	150	283
rect	150	282	151	283
rect	152	282	153	283
rect	153	282	154	283
rect	155	282	156	283
rect	156	282	157	283
rect	157	282	158	283
rect	158	282	159	283
rect	159	282	160	283
rect	161	282	162	283
rect	162	282	163	283
rect	163	282	164	283
rect	164	282	165	283
rect	165	282	166	283
rect	166	282	167	283
rect	173	282	174	283
rect	174	282	175	283
rect	176	282	177	283
rect	177	282	178	283
rect	178	282	179	283
rect	180	282	181	283
rect	181	282	182	283
rect	186	282	187	283
rect	187	282	188	283
rect	189	282	190	283
rect	190	282	191	283
rect	191	282	192	283
rect	192	282	193	283
rect	193	282	194	283
rect	195	282	196	283
rect	196	282	197	283
rect	198	282	199	283
rect	199	282	200	283
rect	275	282	276	283
rect	276	282	277	283
rect	281	282	282	283
rect	282	282	283	283
rect	284	282	285	283
rect	285	282	286	283
rect	286	282	287	283
rect	287	282	288	283
rect	288	282	289	283
rect	290	282	291	283
rect	291	282	292	283
rect	327	282	328	283
rect	328	282	329	283
rect	329	282	330	283
rect	337	282	338	283
rect	338	282	339	283
rect	339	282	340	283
rect	340	282	341	283
rect	342	282	343	283
rect	343	282	344	283
rect	373	282	374	283
rect	374	282	375	283
rect	375	282	376	283
rect	376	282	377	283
rect	377	282	378	283
rect	379	282	380	283
rect	380	282	381	283
rect	382	282	383	283
rect	383	282	384	283
rect	384	282	385	283
rect	385	282	386	283
rect	386	282	387	283
rect	388	282	389	283
rect	389	282	390	283
rect	390	282	391	283
rect	391	282	392	283
rect	392	282	393	283
rect	61	284	62	285
rect	62	284	63	285
rect	67	284	68	285
rect	68	284	69	285
rect	70	284	71	285
rect	71	284	72	285
rect	110	284	111	285
rect	111	284	112	285
rect	128	284	129	285
rect	129	284	130	285
rect	143	284	144	285
rect	144	284	145	285
rect	145	284	146	285
rect	146	284	147	285
rect	147	284	148	285
rect	161	284	162	285
rect	162	284	163	285
rect	163	284	164	285
rect	170	284	171	285
rect	171	284	172	285
rect	172	284	173	285
rect	173	284	174	285
rect	174	284	175	285
rect	176	284	177	285
rect	177	284	178	285
rect	178	284	179	285
rect	180	284	181	285
rect	181	284	182	285
rect	183	284	184	285
rect	184	284	185	285
rect	185	284	186	285
rect	186	284	187	285
rect	187	284	188	285
rect	189	284	190	285
rect	190	284	191	285
rect	191	284	192	285
rect	192	284	193	285
rect	193	284	194	285
rect	195	284	196	285
rect	196	284	197	285
rect	198	284	199	285
rect	199	284	200	285
rect	201	284	202	285
rect	202	284	203	285
rect	207	284	208	285
rect	208	284	209	285
rect	209	284	210	285
rect	210	284	211	285
rect	211	284	212	285
rect	212	284	213	285
rect	213	284	214	285
rect	214	284	215	285
rect	228	284	229	285
rect	229	284	230	285
rect	237	284	238	285
rect	238	284	239	285
rect	239	284	240	285
rect	240	284	241	285
rect	241	284	242	285
rect	242	284	243	285
rect	243	284	244	285
rect	244	284	245	285
rect	245	284	246	285
rect	260	284	261	285
rect	261	284	262	285
rect	263	284	264	285
rect	264	284	265	285
rect	266	284	267	285
rect	267	284	268	285
rect	268	284	269	285
rect	269	284	270	285
rect	270	284	271	285
rect	278	284	279	285
rect	279	284	280	285
rect	280	284	281	285
rect	281	284	282	285
rect	282	284	283	285
rect	321	284	322	285
rect	322	284	323	285
rect	324	284	325	285
rect	325	284	326	285
rect	326	284	327	285
rect	327	284	328	285
rect	328	284	329	285
rect	329	284	330	285
rect	331	284	332	285
rect	332	284	333	285
rect	333	284	334	285
rect	334	284	335	285
rect	335	284	336	285
rect	337	284	338	285
rect	338	284	339	285
rect	339	284	340	285
rect	340	284	341	285
rect	342	284	343	285
rect	343	284	344	285
rect	344	284	345	285
rect	367	284	368	285
rect	368	284	369	285
rect	370	284	371	285
rect	371	284	372	285
rect	372	284	373	285
rect	373	284	374	285
rect	374	284	375	285
rect	37	286	38	287
rect	38	286	39	287
rect	39	286	40	287
rect	40	286	41	287
rect	41	286	42	287
rect	58	286	59	287
rect	59	286	60	287
rect	60	286	61	287
rect	61	286	62	287
rect	62	286	63	287
rect	64	286	65	287
rect	65	286	66	287
rect	101	286	102	287
rect	102	286	103	287
rect	104	286	105	287
rect	105	286	106	287
rect	106	286	107	287
rect	108	286	109	287
rect	110	286	111	287
rect	111	286	112	287
rect	116	286	117	287
rect	117	286	118	287
rect	125	286	126	287
rect	126	286	127	287
rect	127	286	128	287
rect	128	286	129	287
rect	129	286	130	287
rect	131	286	132	287
rect	132	286	133	287
rect	134	286	135	287
rect	135	286	136	287
rect	136	286	137	287
rect	137	286	138	287
rect	138	286	139	287
rect	140	286	141	287
rect	141	286	142	287
rect	142	286	143	287
rect	143	286	144	287
rect	144	286	145	287
rect	152	286	153	287
rect	153	286	154	287
rect	155	286	156	287
rect	156	286	157	287
rect	157	286	158	287
rect	158	286	159	287
rect	159	286	160	287
rect	160	286	161	287
rect	161	286	162	287
rect	162	286	163	287
rect	163	286	164	287
rect	165	286	166	287
rect	166	286	167	287
rect	168	286	169	287
rect	169	286	170	287
rect	176	286	177	287
rect	177	286	178	287
rect	178	286	179	287
rect	180	286	181	287
rect	181	286	182	287
rect	183	286	184	287
rect	184	286	185	287
rect	185	286	186	287
rect	186	286	187	287
rect	187	286	188	287
rect	189	286	190	287
rect	190	286	191	287
rect	198	286	199	287
rect	199	286	200	287
rect	201	286	202	287
rect	202	286	203	287
rect	204	286	205	287
rect	205	286	206	287
rect	207	286	208	287
rect	208	286	209	287
rect	209	286	210	287
rect	210	286	211	287
rect	211	286	212	287
rect	212	286	213	287
rect	213	286	214	287
rect	214	286	215	287
rect	216	286	217	287
rect	217	286	218	287
rect	228	286	229	287
rect	229	286	230	287
rect	231	286	232	287
rect	232	286	233	287
rect	233	286	234	287
rect	234	286	235	287
rect	235	286	236	287
rect	256	286	257	287
rect	257	286	258	287
rect	258	286	259	287
rect	259	286	260	287
rect	260	286	261	287
rect	261	286	262	287
rect	266	286	267	287
rect	267	286	268	287
rect	268	286	269	287
rect	269	286	270	287
rect	270	286	271	287
rect	272	286	273	287
rect	273	286	274	287
rect	275	286	276	287
rect	276	286	277	287
rect	278	286	279	287
rect	279	286	280	287
rect	334	286	335	287
rect	335	286	336	287
rect	337	286	338	287
rect	338	286	339	287
rect	339	286	340	287
rect	340	286	341	287
rect	351	286	352	287
rect	352	286	353	287
rect	353	286	354	287
rect	364	286	365	287
rect	365	286	366	287
rect	366	286	367	287
rect	367	286	368	287
rect	368	286	369	287
rect	370	286	371	287
rect	371	286	372	287
rect	2	288	3	289
rect	3	288	4	289
rect	4	288	5	289
rect	5	288	6	289
rect	6	288	7	289
rect	7	288	8	289
rect	8	288	9	289
rect	9	288	10	289
rect	10	288	11	289
rect	15	288	16	289
rect	16	288	17	289
rect	17	288	18	289
rect	18	288	19	289
rect	19	288	20	289
rect	20	288	21	289
rect	34	288	35	289
rect	35	288	36	289
rect	36	288	37	289
rect	37	288	38	289
rect	38	288	39	289
rect	46	288	47	289
rect	47	288	48	289
rect	48	288	49	289
rect	49	288	50	289
rect	50	288	51	289
rect	55	288	56	289
rect	56	288	57	289
rect	57	288	58	289
rect	58	288	59	289
rect	59	288	60	289
rect	76	288	77	289
rect	77	288	78	289
rect	78	288	79	289
rect	79	288	80	289
rect	80	288	81	289
rect	92	288	93	289
rect	93	288	94	289
rect	94	288	95	289
rect	95	288	96	289
rect	96	288	97	289
rect	101	288	102	289
rect	102	288	103	289
rect	108	288	109	289
rect	110	288	111	289
rect	111	288	112	289
rect	113	288	114	289
rect	114	288	115	289
rect	116	288	117	289
rect	117	288	118	289
rect	122	288	123	289
rect	123	288	124	289
rect	124	288	125	289
rect	125	288	126	289
rect	126	288	127	289
rect	143	288	144	289
rect	144	288	145	289
rect	146	288	147	289
rect	147	288	148	289
rect	149	288	150	289
rect	150	288	151	289
rect	155	288	156	289
rect	156	288	157	289
rect	157	288	158	289
rect	158	288	159	289
rect	159	288	160	289
rect	160	288	161	289
rect	161	288	162	289
rect	162	288	163	289
rect	163	288	164	289
rect	165	288	166	289
rect	166	288	167	289
rect	168	288	169	289
rect	169	288	170	289
rect	171	288	172	289
rect	172	288	173	289
rect	173	288	174	289
rect	174	288	175	289
rect	175	288	176	289
rect	176	288	177	289
rect	177	288	178	289
rect	178	288	179	289
rect	180	288	181	289
rect	181	288	182	289
rect	183	288	184	289
rect	184	288	185	289
rect	195	288	196	289
rect	196	288	197	289
rect	197	288	198	289
rect	198	288	199	289
rect	199	288	200	289
rect	201	288	202	289
rect	202	288	203	289
rect	204	288	205	289
rect	205	288	206	289
rect	207	288	208	289
rect	208	288	209	289
rect	225	288	226	289
rect	226	288	227	289
rect	228	288	229	289
rect	229	288	230	289
rect	231	288	232	289
rect	232	288	233	289
rect	233	288	234	289
rect	234	288	235	289
rect	235	288	236	289
rect	237	288	238	289
rect	238	288	239	289
rect	239	288	240	289
rect	240	288	241	289
rect	241	288	242	289
rect	242	288	243	289
rect	243	288	244	289
rect	244	288	245	289
rect	245	288	246	289
rect	247	288	248	289
rect	248	288	249	289
rect	249	288	250	289
rect	250	288	251	289
rect	251	288	252	289
rect	252	288	253	289
rect	253	288	254	289
rect	254	288	255	289
rect	256	288	257	289
rect	257	288	258	289
rect	258	288	259	289
rect	259	288	260	289
rect	260	288	261	289
rect	261	288	262	289
rect	262	288	263	289
rect	263	288	264	289
rect	264	288	265	289
rect	265	288	266	289
rect	266	288	267	289
rect	267	288	268	289
rect	268	288	269	289
rect	269	288	270	289
rect	270	288	271	289
rect	272	288	273	289
rect	273	288	274	289
rect	275	288	276	289
rect	276	288	277	289
rect	278	288	279	289
rect	279	288	280	289
rect	281	288	282	289
rect	282	288	283	289
rect	283	288	284	289
rect	284	288	285	289
rect	285	288	286	289
rect	286	288	287	289
rect	287	288	288	289
rect	288	288	289	289
rect	290	288	291	289
rect	291	288	292	289
rect	293	288	294	289
rect	294	288	295	289
rect	295	288	296	289
rect	296	288	297	289
rect	297	288	298	289
rect	298	288	299	289
rect	299	288	300	289
rect	300	288	301	289
rect	301	288	302	289
rect	302	288	303	289
rect	303	288	304	289
rect	304	288	305	289
rect	305	288	306	289
rect	306	288	307	289
rect	307	288	308	289
rect	309	288	310	289
rect	310	288	311	289
rect	312	288	313	289
rect	313	288	314	289
rect	314	288	315	289
rect	315	288	316	289
rect	316	288	317	289
rect	317	288	318	289
rect	319	288	320	289
rect	320	288	321	289
rect	321	288	322	289
rect	322	288	323	289
rect	323	288	324	289
rect	325	288	326	289
rect	326	288	327	289
rect	327	288	328	289
rect	328	288	329	289
rect	329	288	330	289
rect	331	288	332	289
rect	332	288	333	289
rect	334	288	335	289
rect	335	288	336	289
rect	337	288	338	289
rect	338	288	339	289
rect	339	288	340	289
rect	340	288	341	289
rect	341	288	342	289
rect	342	288	343	289
rect	343	288	344	289
rect	344	288	345	289
rect	346	288	347	289
rect	347	288	348	289
rect	348	288	349	289
rect	349	288	350	289
rect	350	288	351	289
rect	364	288	365	289
rect	365	288	366	289
rect	366	288	367	289
rect	367	288	368	289
rect	368	288	369	289
rect	134	297	135	298
rect	135	297	136	298
rect	136	297	137	298
rect	204	297	205	298
rect	205	297	206	298
rect	207	297	208	298
rect	208	297	209	298
rect	210	297	211	298
rect	211	297	212	298
rect	212	297	213	298
rect	213	297	214	298
rect	214	297	215	298
rect	215	297	216	298
rect	216	297	217	298
rect	217	297	218	298
rect	219	297	220	298
rect	220	297	221	298
rect	221	297	222	298
rect	222	297	223	298
rect	223	297	224	298
rect	225	297	226	298
rect	226	297	227	298
rect	228	297	229	298
rect	229	297	230	298
rect	231	297	232	298
rect	232	297	233	298
rect	234	297	235	298
rect	235	297	236	298
rect	236	297	237	298
rect	237	297	238	298
rect	238	297	239	298
rect	239	297	240	298
rect	240	297	241	298
rect	241	297	242	298
rect	247	297	248	298
rect	248	297	249	298
rect	249	297	250	298
rect	250	297	251	298
rect	131	299	132	300
rect	132	299	133	300
rect	133	299	134	300
rect	186	299	187	300
rect	187	299	188	300
rect	189	299	190	300
rect	190	299	191	300
rect	192	299	193	300
rect	193	299	194	300
rect	194	299	195	300
rect	195	299	196	300
rect	196	299	197	300
rect	198	299	199	300
rect	199	299	200	300
rect	201	299	202	300
rect	202	299	203	300
rect	219	299	220	300
rect	220	299	221	300
rect	221	299	222	300
rect	222	299	223	300
rect	223	299	224	300
rect	225	299	226	300
rect	226	299	227	300
rect	228	299	229	300
rect	229	299	230	300
rect	231	299	232	300
rect	232	299	233	300
rect	234	299	235	300
rect	235	299	236	300
rect	236	299	237	300
rect	237	299	238	300
rect	238	299	239	300
rect	239	299	240	300
rect	240	299	241	300
rect	241	299	242	300
rect	243	299	244	300
rect	244	299	245	300
rect	113	301	114	302
rect	114	301	115	302
rect	116	301	117	302
rect	117	301	118	302
rect	119	301	120	302
rect	120	301	121	302
rect	122	301	123	302
rect	123	301	124	302
rect	125	301	126	302
rect	126	301	127	302
rect	128	301	129	302
rect	129	301	130	302
rect	130	301	131	302
rect	177	301	178	302
rect	178	301	179	302
rect	180	301	181	302
rect	181	301	182	302
rect	183	301	184	302
rect	184	301	185	302
rect	207	301	208	302
rect	208	301	209	302
rect	210	301	211	302
rect	211	301	212	302
rect	212	301	213	302
rect	213	301	214	302
rect	214	301	215	302
rect	215	301	216	302
rect	216	301	217	302
rect	217	301	218	302
rect	218	301	219	302
rect	219	301	220	302
rect	220	301	221	302
rect	288	301	289	302
rect	290	301	291	302
rect	291	301	292	302
rect	388	301	389	302
rect	389	301	390	302
rect	391	301	392	302
rect	392	301	393	302
rect	393	301	394	302
rect	114	303	115	304
rect	116	303	117	304
rect	117	303	118	304
rect	119	303	120	304
rect	120	303	121	304
rect	122	303	123	304
rect	123	303	124	304
rect	177	303	178	304
rect	178	303	179	304
rect	180	303	181	304
rect	181	303	182	304
rect	183	303	184	304
rect	184	303	185	304
rect	186	303	187	304
rect	187	303	188	304
rect	201	303	202	304
rect	202	303	203	304
rect	204	303	205	304
rect	205	303	206	304
rect	206	303	207	304
rect	207	303	208	304
rect	208	303	209	304
rect	210	303	211	304
rect	211	303	212	304
rect	212	303	213	304
rect	213	303	214	304
rect	214	303	215	304
rect	215	303	216	304
rect	216	303	217	304
rect	217	303	218	304
rect	270	303	271	304
rect	281	303	282	304
rect	282	303	283	304
rect	283	303	284	304
rect	284	303	285	304
rect	285	303	286	304
rect	286	303	287	304
rect	288	303	289	304
rect	290	303	291	304
rect	291	303	292	304
rect	292	303	293	304
rect	358	303	359	304
rect	359	303	360	304
rect	361	303	362	304
rect	362	303	363	304
rect	364	303	365	304
rect	365	303	366	304
rect	367	303	368	304
rect	368	303	369	304
rect	369	303	370	304
rect	370	303	371	304
rect	371	303	372	304
rect	373	303	374	304
rect	374	303	375	304
rect	376	303	377	304
rect	377	303	378	304
rect	379	303	380	304
rect	380	303	381	304
rect	381	303	382	304
rect	382	303	383	304
rect	383	303	384	304
rect	385	303	386	304
rect	386	303	387	304
rect	387	303	388	304
rect	126	305	127	306
rect	140	305	141	306
rect	141	305	142	306
rect	143	305	144	306
rect	144	305	145	306
rect	146	305	147	306
rect	147	305	148	306
rect	149	305	150	306
rect	150	305	151	306
rect	151	305	152	306
rect	171	305	172	306
rect	172	305	173	306
rect	173	305	174	306
rect	174	305	175	306
rect	175	305	176	306
rect	177	305	178	306
rect	178	305	179	306
rect	180	305	181	306
rect	181	305	182	306
rect	183	305	184	306
rect	184	305	185	306
rect	186	305	187	306
rect	187	305	188	306
rect	198	305	199	306
rect	199	305	200	306
rect	200	305	201	306
rect	201	305	202	306
rect	202	305	203	306
rect	204	305	205	306
rect	205	305	206	306
rect	206	305	207	306
rect	207	305	208	306
rect	208	305	209	306
rect	210	305	211	306
rect	211	305	212	306
rect	212	305	213	306
rect	213	305	214	306
rect	214	305	215	306
rect	234	305	235	306
rect	235	305	236	306
rect	236	305	237	306
rect	237	305	238	306
rect	238	305	239	306
rect	239	305	240	306
rect	240	305	241	306
rect	241	305	242	306
rect	243	305	244	306
rect	244	305	245	306
rect	246	305	247	306
rect	247	305	248	306
rect	248	305	249	306
rect	249	305	250	306
rect	250	305	251	306
rect	252	305	253	306
rect	253	305	254	306
rect	254	305	255	306
rect	256	305	257	306
rect	257	305	258	306
rect	258	305	259	306
rect	259	305	260	306
rect	260	305	261	306
rect	261	305	262	306
rect	262	305	263	306
rect	263	305	264	306
rect	264	305	265	306
rect	265	305	266	306
rect	266	305	267	306
rect	267	305	268	306
rect	268	305	269	306
rect	270	305	271	306
rect	271	305	272	306
rect	272	305	273	306
rect	273	305	274	306
rect	275	305	276	306
rect	276	305	277	306
rect	278	305	279	306
rect	279	305	280	306
rect	280	305	281	306
rect	359	305	360	306
rect	361	305	362	306
rect	362	305	363	306
rect	73	307	74	308
rect	74	307	75	308
rect	75	307	76	308
rect	76	307	77	308
rect	77	307	78	308
rect	78	307	79	308
rect	79	307	80	308
rect	80	307	81	308
rect	82	307	83	308
rect	96	307	97	308
rect	98	307	99	308
rect	99	307	100	308
rect	129	307	130	308
rect	130	307	131	308
rect	132	307	133	308
rect	133	307	134	308
rect	135	307	136	308
rect	136	307	137	308
rect	138	307	139	308
rect	139	307	140	308
rect	140	307	141	308
rect	141	307	142	308
rect	143	307	144	308
rect	144	307	145	308
rect	146	307	147	308
rect	147	307	148	308
rect	165	307	166	308
rect	166	307	167	308
rect	168	307	169	308
rect	169	307	170	308
rect	192	307	193	308
rect	193	307	194	308
rect	194	307	195	308
rect	195	307	196	308
rect	196	307	197	308
rect	197	307	198	308
rect	198	307	199	308
rect	199	307	200	308
rect	200	307	201	308
rect	201	307	202	308
rect	202	307	203	308
rect	204	307	205	308
rect	205	307	206	308
rect	234	307	235	308
rect	235	307	236	308
rect	236	307	237	308
rect	237	307	238	308
rect	238	307	239	308
rect	273	307	274	308
rect	275	307	276	308
rect	276	307	277	308
rect	278	307	279	308
rect	279	307	280	308
rect	280	307	281	308
rect	282	307	283	308
rect	283	307	284	308
rect	284	307	285	308
rect	285	307	286	308
rect	286	307	287	308
rect	288	307	289	308
rect	349	307	350	308
rect	350	307	351	308
rect	351	307	352	308
rect	352	307	353	308
rect	353	307	354	308
rect	355	307	356	308
rect	356	307	357	308
rect	357	307	358	308
rect	359	307	360	308
rect	67	309	68	310
rect	68	309	69	310
rect	70	309	71	310
rect	71	309	72	310
rect	72	309	73	310
rect	73	309	74	310
rect	74	309	75	310
rect	75	309	76	310
rect	76	309	77	310
rect	102	309	103	310
rect	103	309	104	310
rect	104	309	105	310
rect	105	309	106	310
rect	106	309	107	310
rect	107	309	108	310
rect	108	309	109	310
rect	122	309	123	310
rect	123	309	124	310
rect	124	309	125	310
rect	126	309	127	310
rect	127	309	128	310
rect	129	309	130	310
rect	130	309	131	310
rect	132	309	133	310
rect	133	309	134	310
rect	135	309	136	310
rect	136	309	137	310
rect	138	309	139	310
rect	139	309	140	310
rect	140	309	141	310
rect	141	309	142	310
rect	143	309	144	310
rect	144	309	145	310
rect	146	309	147	310
rect	147	309	148	310
rect	148	309	149	310
rect	149	309	150	310
rect	150	309	151	310
rect	151	309	152	310
rect	153	309	154	310
rect	154	309	155	310
rect	155	309	156	310
rect	156	309	157	310
rect	157	309	158	310
rect	159	309	160	310
rect	160	309	161	310
rect	161	309	162	310
rect	162	309	163	310
rect	163	309	164	310
rect	164	309	165	310
rect	165	309	166	310
rect	166	309	167	310
rect	168	309	169	310
rect	169	309	170	310
rect	171	309	172	310
rect	172	309	173	310
rect	173	309	174	310
rect	174	309	175	310
rect	175	309	176	310
rect	177	309	178	310
rect	178	309	179	310
rect	180	309	181	310
rect	181	309	182	310
rect	183	309	184	310
rect	184	309	185	310
rect	186	309	187	310
rect	187	309	188	310
rect	189	309	190	310
rect	190	309	191	310
rect	191	309	192	310
rect	192	309	193	310
rect	193	309	194	310
rect	194	309	195	310
rect	195	309	196	310
rect	196	309	197	310
rect	197	309	198	310
rect	198	309	199	310
rect	199	309	200	310
rect	200	309	201	310
rect	201	309	202	310
rect	202	309	203	310
rect	204	309	205	310
rect	205	309	206	310
rect	207	309	208	310
rect	208	309	209	310
rect	210	309	211	310
rect	211	309	212	310
rect	212	309	213	310
rect	213	309	214	310
rect	214	309	215	310
rect	216	309	217	310
rect	217	309	218	310
rect	219	309	220	310
rect	220	309	221	310
rect	222	309	223	310
rect	223	309	224	310
rect	225	309	226	310
rect	226	309	227	310
rect	228	309	229	310
rect	229	309	230	310
rect	231	309	232	310
rect	232	309	233	310
rect	234	309	235	310
rect	235	309	236	310
rect	236	309	237	310
rect	237	309	238	310
rect	238	309	239	310
rect	240	309	241	310
rect	241	309	242	310
rect	243	309	244	310
rect	244	309	245	310
rect	246	309	247	310
rect	247	309	248	310
rect	248	309	249	310
rect	249	309	250	310
rect	250	309	251	310
rect	252	309	253	310
rect	253	309	254	310
rect	254	309	255	310
rect	256	309	257	310
rect	257	309	258	310
rect	258	309	259	310
rect	259	309	260	310
rect	260	309	261	310
rect	261	309	262	310
rect	262	309	263	310
rect	263	309	264	310
rect	264	309	265	310
rect	265	309	266	310
rect	266	309	267	310
rect	267	309	268	310
rect	268	309	269	310
rect	270	309	271	310
rect	271	309	272	310
rect	273	309	274	310
rect	275	309	276	310
rect	276	309	277	310
rect	278	309	279	310
rect	279	309	280	310
rect	280	309	281	310
rect	282	309	283	310
rect	283	309	284	310
rect	284	309	285	310
rect	285	309	286	310
rect	286	309	287	310
rect	288	309	289	310
rect	289	309	290	310
rect	290	309	291	310
rect	291	309	292	310
rect	292	309	293	310
rect	294	309	295	310
rect	295	309	296	310
rect	296	309	297	310
rect	297	309	298	310
rect	298	309	299	310
rect	299	309	300	310
rect	300	309	301	310
rect	301	309	302	310
rect	302	309	303	310
rect	303	309	304	310
rect	304	309	305	310
rect	305	309	306	310
rect	306	309	307	310
rect	307	309	308	310
rect	309	309	310	310
rect	310	309	311	310
rect	312	309	313	310
rect	313	309	314	310
rect	314	309	315	310
rect	315	309	316	310
rect	316	309	317	310
rect	317	309	318	310
rect	318	309	319	310
rect	319	309	320	310
rect	320	309	321	310
rect	321	309	322	310
rect	322	309	323	310
rect	323	309	324	310
rect	325	309	326	310
rect	326	309	327	310
rect	327	309	328	310
rect	328	309	329	310
rect	329	309	330	310
rect	330	309	331	310
rect	331	309	332	310
rect	332	309	333	310
rect	334	309	335	310
rect	335	309	336	310
rect	337	309	338	310
rect	338	309	339	310
rect	339	309	340	310
rect	340	309	341	310
rect	341	309	342	310
rect	342	309	343	310
rect	343	309	344	310
rect	344	309	345	310
rect	346	309	347	310
rect	347	309	348	310
rect	348	309	349	310
rect	349	309	350	310
rect	350	309	351	310
rect	351	309	352	310
rect	352	309	353	310
rect	353	309	354	310
rect	355	309	356	310
rect	356	309	357	310
rect	357	309	358	310
rect	359	309	360	310
rect	360	309	361	310
rect	361	309	362	310
rect	362	309	363	310
rect	363	309	364	310
rect	364	309	365	310
rect	365	309	366	310
rect	367	309	368	310
rect	368	309	369	310
rect	369	309	370	310
rect	370	309	371	310
rect	371	309	372	310
rect	373	309	374	310
rect	374	309	375	310
rect	376	309	377	310
rect	377	309	378	310
rect	379	309	380	310
rect	380	309	381	310
rect	381	309	382	310
rect	382	309	383	310
rect	383	309	384	310
rect	385	309	386	310
rect	386	309	387	310
rect	387	309	388	310
rect	389	309	390	310
rect	391	309	392	310
rect	392	309	393	310
rect	393	309	394	310
rect	395	309	396	310
rect	396	309	397	310
rect	397	309	398	310
rect	398	309	399	310
rect	399	309	400	310
rect	401	309	402	310
rect	402	309	403	310
rect	403	309	404	310
rect	404	309	405	310
rect	405	309	406	310
rect	406	309	407	310
rect	407	309	408	310
rect	408	309	409	310
rect	409	309	410	310
rect	410	309	411	310
rect	411	309	412	310
rect	412	309	413	310
rect	2	311	3	312
rect	3	311	4	312
rect	5	311	6	312
rect	6	311	7	312
rect	7	311	8	312
rect	9	311	10	312
rect	10	311	11	312
rect	11	311	12	312
rect	12	311	13	312
rect	13	311	14	312
rect	43	311	44	312
rect	44	311	45	312
rect	45	311	46	312
rect	46	311	47	312
rect	64	311	65	312
rect	65	311	66	312
rect	66	311	67	312
rect	67	311	68	312
rect	68	311	69	312
rect	70	311	71	312
rect	71	311	72	312
rect	72	311	73	312
rect	73	311	74	312
rect	82	311	83	312
rect	84	311	85	312
rect	85	311	86	312
rect	86	311	87	312
rect	87	311	88	312
rect	88	311	89	312
rect	89	311	90	312
rect	90	311	91	312
rect	91	311	92	312
rect	96	311	97	312
rect	98	311	99	312
rect	99	311	100	312
rect	100	311	101	312
rect	102	311	103	312
rect	103	311	104	312
rect	104	311	105	312
rect	105	311	106	312
rect	106	311	107	312
rect	107	311	108	312
rect	108	311	109	312
rect	109	311	110	312
rect	123	311	124	312
rect	124	311	125	312
rect	126	311	127	312
rect	127	311	128	312
rect	129	311	130	312
rect	130	311	131	312
rect	132	311	133	312
rect	133	311	134	312
rect	135	311	136	312
rect	136	311	137	312
rect	138	311	139	312
rect	139	311	140	312
rect	140	311	141	312
rect	141	311	142	312
rect	146	311	147	312
rect	147	311	148	312
rect	148	311	149	312
rect	149	311	150	312
rect	150	311	151	312
rect	151	311	152	312
rect	153	311	154	312
rect	154	311	155	312
rect	162	311	163	312
rect	163	311	164	312
rect	183	311	184	312
rect	184	311	185	312
rect	186	311	187	312
rect	187	311	188	312
rect	189	311	190	312
rect	190	311	191	312
rect	191	311	192	312
rect	192	311	193	312
rect	193	311	194	312
rect	194	311	195	312
rect	195	311	196	312
rect	196	311	197	312
rect	197	311	198	312
rect	198	311	199	312
rect	199	311	200	312
rect	225	311	226	312
rect	226	311	227	312
rect	228	311	229	312
rect	229	311	230	312
rect	231	311	232	312
rect	232	311	233	312
rect	234	311	235	312
rect	235	311	236	312
rect	236	311	237	312
rect	237	311	238	312
rect	238	311	239	312
rect	240	311	241	312
rect	241	311	242	312
rect	243	311	244	312
rect	244	311	245	312
rect	246	311	247	312
rect	247	311	248	312
rect	248	311	249	312
rect	249	311	250	312
rect	250	311	251	312
rect	252	311	253	312
rect	253	311	254	312
rect	254	311	255	312
rect	256	311	257	312
rect	257	311	258	312
rect	258	311	259	312
rect	259	311	260	312
rect	260	311	261	312
rect	261	311	262	312
rect	262	311	263	312
rect	263	311	264	312
rect	264	311	265	312
rect	265	311	266	312
rect	266	311	267	312
rect	267	311	268	312
rect	268	311	269	312
rect	270	311	271	312
rect	271	311	272	312
rect	273	311	274	312
rect	275	311	276	312
rect	276	311	277	312
rect	278	311	279	312
rect	279	311	280	312
rect	280	311	281	312
rect	282	311	283	312
rect	283	311	284	312
rect	284	311	285	312
rect	285	311	286	312
rect	286	311	287	312
rect	288	311	289	312
rect	289	311	290	312
rect	290	311	291	312
rect	291	311	292	312
rect	292	311	293	312
rect	294	311	295	312
rect	295	311	296	312
rect	296	311	297	312
rect	297	311	298	312
rect	298	311	299	312
rect	299	311	300	312
rect	300	311	301	312
rect	301	311	302	312
rect	302	311	303	312
rect	303	311	304	312
rect	304	311	305	312
rect	305	311	306	312
rect	306	311	307	312
rect	307	311	308	312
rect	309	311	310	312
rect	310	311	311	312
rect	312	311	313	312
rect	313	311	314	312
rect	314	311	315	312
rect	315	311	316	312
rect	316	311	317	312
rect	317	311	318	312
rect	318	311	319	312
rect	319	311	320	312
rect	320	311	321	312
rect	321	311	322	312
rect	322	311	323	312
rect	323	311	324	312
rect	325	311	326	312
rect	326	311	327	312
rect	327	311	328	312
rect	328	311	329	312
rect	329	311	330	312
rect	330	311	331	312
rect	331	311	332	312
rect	332	311	333	312
rect	334	311	335	312
rect	335	311	336	312
rect	337	311	338	312
rect	338	311	339	312
rect	339	311	340	312
rect	340	311	341	312
rect	341	311	342	312
rect	342	311	343	312
rect	343	311	344	312
rect	344	311	345	312
rect	346	311	347	312
rect	347	311	348	312
rect	348	311	349	312
rect	349	311	350	312
rect	350	311	351	312
rect	351	311	352	312
rect	352	311	353	312
rect	353	311	354	312
rect	355	311	356	312
rect	356	311	357	312
rect	357	311	358	312
rect	359	311	360	312
rect	360	311	361	312
rect	5	313	6	314
rect	6	313	7	314
rect	7	313	8	314
rect	15	313	16	314
rect	16	313	17	314
rect	17	313	18	314
rect	18	313	19	314
rect	19	313	20	314
rect	20	313	21	314
rect	21	313	22	314
rect	22	313	23	314
rect	40	313	41	314
rect	41	313	42	314
rect	42	313	43	314
rect	43	313	44	314
rect	52	313	53	314
rect	53	313	54	314
rect	54	313	55	314
rect	55	313	56	314
rect	61	313	62	314
rect	62	313	63	314
rect	63	313	64	314
rect	64	313	65	314
rect	70	313	71	314
rect	71	313	72	314
rect	72	313	73	314
rect	73	313	74	314
rect	75	313	76	314
rect	76	313	77	314
rect	78	313	79	314
rect	79	313	80	314
rect	98	313	99	314
rect	99	313	100	314
rect	100	313	101	314
rect	102	313	103	314
rect	103	313	104	314
rect	108	313	109	314
rect	109	313	110	314
rect	111	313	112	314
rect	112	313	113	314
rect	114	313	115	314
rect	119	313	120	314
rect	120	313	121	314
rect	121	313	122	314
rect	123	313	124	314
rect	124	313	125	314
rect	126	313	127	314
rect	127	313	128	314
rect	129	313	130	314
rect	130	313	131	314
rect	132	313	133	314
rect	133	313	134	314
rect	135	313	136	314
rect	136	313	137	314
rect	138	313	139	314
rect	139	313	140	314
rect	147	313	148	314
rect	148	313	149	314
rect	159	313	160	314
rect	160	313	161	314
rect	162	313	163	314
rect	163	313	164	314
rect	165	313	166	314
rect	166	313	167	314
rect	168	313	169	314
rect	169	313	170	314
rect	171	313	172	314
rect	172	313	173	314
rect	180	313	181	314
rect	181	313	182	314
rect	182	313	183	314
rect	183	313	184	314
rect	184	313	185	314
rect	186	313	187	314
rect	187	313	188	314
rect	189	313	190	314
rect	190	313	191	314
rect	191	313	192	314
rect	192	313	193	314
rect	193	313	194	314
rect	194	313	195	314
rect	195	313	196	314
rect	196	313	197	314
rect	210	313	211	314
rect	211	313	212	314
rect	212	313	213	314
rect	213	313	214	314
rect	214	313	215	314
rect	216	313	217	314
rect	217	313	218	314
rect	219	313	220	314
rect	220	313	221	314
rect	222	313	223	314
rect	223	313	224	314
rect	231	313	232	314
rect	232	313	233	314
rect	234	313	235	314
rect	235	313	236	314
rect	278	313	279	314
rect	279	313	280	314
rect	280	313	281	314
rect	282	313	283	314
rect	283	313	284	314
rect	284	313	285	314
rect	285	313	286	314
rect	286	313	287	314
rect	288	313	289	314
rect	289	313	290	314
rect	355	313	356	314
rect	356	313	357	314
rect	357	313	358	314
rect	359	313	360	314
rect	360	313	361	314
rect	362	313	363	314
rect	363	313	364	314
rect	364	313	365	314
rect	365	313	366	314
rect	373	313	374	314
rect	374	313	375	314
rect	376	313	377	314
rect	377	313	378	314
rect	378	313	379	314
rect	380	313	381	314
rect	381	313	382	314
rect	382	313	383	314
rect	383	313	384	314
rect	391	313	392	314
rect	392	313	393	314
rect	393	313	394	314
rect	395	313	396	314
rect	396	313	397	314
rect	397	313	398	314
rect	398	313	399	314
rect	399	313	400	314
rect	401	313	402	314
rect	402	313	403	314
rect	403	313	404	314
rect	404	313	405	314
rect	405	313	406	314
rect	406	313	407	314
rect	407	313	408	314
rect	408	313	409	314
rect	409	313	410	314
rect	5	315	6	316
rect	6	315	7	316
rect	7	315	8	316
rect	8	315	9	316
rect	9	315	10	316
rect	10	315	11	316
rect	11	315	12	316
rect	12	315	13	316
rect	13	315	14	316
rect	15	315	16	316
rect	16	315	17	316
rect	17	315	18	316
rect	18	315	19	316
rect	19	315	20	316
rect	20	315	21	316
rect	21	315	22	316
rect	22	315	23	316
rect	23	315	24	316
rect	24	315	25	316
rect	25	315	26	316
rect	26	315	27	316
rect	27	315	28	316
rect	28	315	29	316
rect	29	315	30	316
rect	30	315	31	316
rect	31	315	32	316
rect	32	315	33	316
rect	33	315	34	316
rect	34	315	35	316
rect	35	315	36	316
rect	36	315	37	316
rect	37	315	38	316
rect	38	315	39	316
rect	39	315	40	316
rect	40	315	41	316
rect	41	315	42	316
rect	42	315	43	316
rect	43	315	44	316
rect	45	315	46	316
rect	46	315	47	316
rect	48	315	49	316
rect	49	315	50	316
rect	50	315	51	316
rect	51	315	52	316
rect	52	315	53	316
rect	53	315	54	316
rect	54	315	55	316
rect	55	315	56	316
rect	57	315	58	316
rect	58	315	59	316
rect	59	315	60	316
rect	60	315	61	316
rect	61	315	62	316
rect	62	315	63	316
rect	63	315	64	316
rect	64	315	65	316
rect	66	315	67	316
rect	67	315	68	316
rect	68	315	69	316
rect	69	315	70	316
rect	70	315	71	316
rect	71	315	72	316
rect	72	315	73	316
rect	73	315	74	316
rect	75	315	76	316
rect	76	315	77	316
rect	78	315	79	316
rect	79	315	80	316
rect	81	315	82	316
rect	82	315	83	316
rect	84	315	85	316
rect	85	315	86	316
rect	86	315	87	316
rect	87	315	88	316
rect	88	315	89	316
rect	89	315	90	316
rect	90	315	91	316
rect	91	315	92	316
rect	93	315	94	316
rect	94	315	95	316
rect	95	315	96	316
rect	96	315	97	316
rect	97	315	98	316
rect	98	315	99	316
rect	99	315	100	316
rect	100	315	101	316
rect	102	315	103	316
rect	103	315	104	316
rect	105	315	106	316
rect	106	315	107	316
rect	108	315	109	316
rect	109	315	110	316
rect	111	315	112	316
rect	112	315	113	316
rect	114	315	115	316
rect	115	315	116	316
rect	116	315	117	316
rect	117	315	118	316
rect	118	315	119	316
rect	119	315	120	316
rect	120	315	121	316
rect	121	315	122	316
rect	123	315	124	316
rect	124	315	125	316
rect	126	315	127	316
rect	127	315	128	316
rect	129	315	130	316
rect	130	315	131	316
rect	132	315	133	316
rect	133	315	134	316
rect	135	315	136	316
rect	136	315	137	316
rect	138	315	139	316
rect	139	315	140	316
rect	141	315	142	316
rect	142	315	143	316
rect	143	315	144	316
rect	144	315	145	316
rect	145	315	146	316
rect	147	315	148	316
rect	148	315	149	316
rect	150	315	151	316
rect	151	315	152	316
rect	153	315	154	316
rect	154	315	155	316
rect	156	315	157	316
rect	157	315	158	316
rect	158	315	159	316
rect	159	315	160	316
rect	160	315	161	316
rect	162	315	163	316
rect	163	315	164	316
rect	165	315	166	316
rect	166	315	167	316
rect	168	315	169	316
rect	169	315	170	316
rect	171	315	172	316
rect	172	315	173	316
rect	174	315	175	316
rect	175	315	176	316
rect	177	315	178	316
rect	178	315	179	316
rect	179	315	180	316
rect	180	315	181	316
rect	181	315	182	316
rect	182	315	183	316
rect	183	315	184	316
rect	184	315	185	316
rect	186	315	187	316
rect	187	315	188	316
rect	189	315	190	316
rect	190	315	191	316
rect	191	315	192	316
rect	192	315	193	316
rect	193	315	194	316
rect	194	315	195	316
rect	195	315	196	316
rect	196	315	197	316
rect	198	315	199	316
rect	199	315	200	316
rect	201	315	202	316
rect	202	315	203	316
rect	204	315	205	316
rect	205	315	206	316
rect	207	315	208	316
rect	208	315	209	316
rect	209	315	210	316
rect	210	315	211	316
rect	211	315	212	316
rect	228	315	229	316
rect	229	315	230	316
rect	230	315	231	316
rect	231	315	232	316
rect	232	315	233	316
rect	234	315	235	316
rect	235	315	236	316
rect	237	315	238	316
rect	238	315	239	316
rect	240	315	241	316
rect	241	315	242	316
rect	243	315	244	316
rect	244	315	245	316
rect	246	315	247	316
rect	247	315	248	316
rect	256	315	257	316
rect	257	315	258	316
rect	258	315	259	316
rect	259	315	260	316
rect	275	315	276	316
rect	276	315	277	316
rect	277	315	278	316
rect	278	315	279	316
rect	279	315	280	316
rect	280	315	281	316
rect	282	315	283	316
rect	283	315	284	316
rect	309	315	310	316
rect	310	315	311	316
rect	346	315	347	316
rect	347	315	348	316
rect	348	315	349	316
rect	349	315	350	316
rect	350	315	351	316
rect	351	315	352	316
rect	352	315	353	316
rect	353	315	354	316
rect	354	315	355	316
rect	355	315	356	316
rect	356	315	357	316
rect	357	315	358	316
rect	359	315	360	316
rect	360	315	361	316
rect	362	315	363	316
rect	363	315	364	316
rect	364	315	365	316
rect	365	315	366	316
rect	366	315	367	316
rect	367	315	368	316
rect	368	315	369	316
rect	369	315	370	316
rect	376	315	377	316
rect	377	315	378	316
rect	378	315	379	316
rect	380	315	381	316
rect	381	315	382	316
rect	382	315	383	316
rect	383	315	384	316
rect	384	315	385	316
rect	385	315	386	316
rect	386	315	387	316
rect	387	315	388	316
rect	389	315	390	316
rect	390	315	391	316
rect	401	315	402	316
rect	402	315	403	316
rect	403	315	404	316
rect	404	315	405	316
rect	405	315	406	316
rect	406	315	407	316
rect	407	315	408	316
rect	408	315	409	316
rect	409	315	410	316
rect	411	315	412	316
rect	412	315	413	316
rect	414	315	415	316
rect	415	315	416	316
rect	416	315	417	316
rect	417	315	418	316
rect	418	315	419	316
rect	214	324	215	325
rect	216	324	217	325
rect	217	324	218	325
rect	219	324	220	325
rect	220	324	221	325
rect	222	324	223	325
rect	223	324	224	325
rect	225	324	226	325
rect	226	324	227	325
rect	227	324	228	325
rect	228	324	229	325
rect	229	324	230	325
rect	230	326	231	327
rect	231	326	232	327
rect	232	326	233	327
rect	234	326	235	327
rect	235	326	236	327
rect	148	328	149	329
rect	150	328	151	329
rect	151	328	152	329
rect	153	328	154	329
rect	154	328	155	329
rect	156	328	157	329
rect	157	328	158	329
rect	158	328	159	329
rect	159	328	160	329
rect	160	328	161	329
rect	161	328	162	329
rect	162	328	163	329
rect	163	328	164	329
rect	165	328	166	329
rect	166	328	167	329
rect	168	328	169	329
rect	169	328	170	329
rect	171	328	172	329
rect	172	328	173	329
rect	214	328	215	329
rect	216	328	217	329
rect	217	328	218	329
rect	219	328	220	329
rect	220	328	221	329
rect	222	328	223	329
rect	223	328	224	329
rect	225	328	226	329
rect	226	328	227	329
rect	227	328	228	329
rect	228	328	229	329
rect	230	328	231	329
rect	231	328	232	329
rect	232	328	233	329
rect	234	328	235	329
rect	294	328	295	329
rect	295	328	296	329
rect	296	328	297	329
rect	297	328	298	329
rect	298	328	299	329
rect	299	328	300	329
rect	300	328	301	329
rect	301	328	302	329
rect	302	328	303	329
rect	303	328	304	329
rect	304	328	305	329
rect	305	328	306	329
rect	306	328	307	329
rect	307	328	308	329
rect	308	328	309	329
rect	309	328	310	329
rect	310	328	311	329
rect	311	328	312	329
rect	312	328	313	329
rect	313	328	314	329
rect	314	328	315	329
rect	315	328	316	329
rect	316	328	317	329
rect	317	328	318	329
rect	318	328	319	329
rect	319	328	320	329
rect	320	328	321	329
rect	321	328	322	329
rect	322	328	323	329
rect	324	328	325	329
rect	325	328	326	329
rect	326	328	327	329
rect	327	328	328	329
rect	328	328	329	329
rect	329	328	330	329
rect	330	328	331	329
rect	331	328	332	329
rect	333	328	334	329
rect	334	328	335	329
rect	336	328	337	329
rect	337	328	338	329
rect	339	328	340	329
rect	340	328	341	329
rect	341	328	342	329
rect	342	328	343	329
rect	343	328	344	329
rect	344	328	345	329
rect	345	328	346	329
rect	346	328	347	329
rect	347	328	348	329
rect	175	330	176	331
rect	177	330	178	331
rect	178	330	179	331
rect	180	330	181	331
rect	181	330	182	331
rect	182	330	183	331
rect	183	330	184	331
rect	184	330	185	331
rect	186	330	187	331
rect	187	330	188	331
rect	189	330	190	331
rect	190	330	191	331
rect	227	330	228	331
rect	228	330	229	331
rect	230	330	231	331
rect	231	330	232	331
rect	232	330	233	331
rect	306	330	307	331
rect	307	330	308	331
rect	308	330	309	331
rect	309	330	310	331
rect	310	330	311	331
rect	311	330	312	331
rect	312	330	313	331
rect	313	330	314	331
rect	314	330	315	331
rect	315	330	316	331
rect	316	330	317	331
rect	317	330	318	331
rect	318	330	319	331
rect	319	330	320	331
rect	320	330	321	331
rect	321	330	322	331
rect	322	330	323	331
rect	350	330	351	331
rect	351	330	352	331
rect	352	330	353	331
rect	353	330	354	331
rect	354	330	355	331
rect	355	330	356	331
rect	356	330	357	331
rect	357	330	358	331
rect	359	330	360	331
rect	360	330	361	331
rect	193	332	194	333
rect	194	332	195	333
rect	195	332	196	333
rect	196	332	197	333
rect	198	332	199	333
rect	199	332	200	333
rect	233	332	234	333
rect	234	332	235	333
rect	236	332	237	333
rect	237	332	238	333
rect	238	332	239	333
rect	239	332	240	333
rect	240	332	241	333
rect	241	332	242	333
rect	242	332	243	333
rect	243	332	244	333
rect	244	332	245	333
rect	246	332	247	333
rect	247	332	248	333
rect	257	332	258	333
rect	258	332	259	333
rect	259	332	260	333
rect	324	332	325	333
rect	325	332	326	333
rect	326	332	327	333
rect	327	332	328	333
rect	328	332	329	333
rect	329	332	330	333
rect	330	332	331	333
rect	331	332	332	333
rect	333	332	334	333
rect	334	332	335	333
rect	336	332	337	333
rect	337	332	338	333
rect	339	332	340	333
rect	340	332	341	333
rect	341	332	342	333
rect	342	332	343	333
rect	343	332	344	333
rect	344	332	345	333
rect	345	332	346	333
rect	346	332	347	333
rect	347	332	348	333
rect	348	332	349	333
rect	350	332	351	333
rect	351	332	352	333
rect	352	332	353	333
rect	353	332	354	333
rect	354	332	355	333
rect	355	332	356	333
rect	356	332	357	333
rect	357	332	358	333
rect	359	332	360	333
rect	360	332	361	333
rect	202	334	203	335
rect	204	334	205	335
rect	205	334	206	335
rect	207	334	208	335
rect	208	334	209	335
rect	209	334	210	335
rect	210	334	211	335
rect	211	334	212	335
rect	212	334	213	335
rect	213	334	214	335
rect	214	334	215	335
rect	246	334	247	335
rect	260	334	261	335
rect	261	334	262	335
rect	262	334	263	335
rect	263	334	264	335
rect	264	334	265	335
rect	265	334	266	335
rect	266	334	267	335
rect	267	334	268	335
rect	268	334	269	335
rect	278	334	279	335
rect	279	334	280	335
rect	280	334	281	335
rect	321	334	322	335
rect	322	334	323	335
rect	324	334	325	335
rect	325	334	326	335
rect	326	334	327	335
rect	327	334	328	335
rect	328	334	329	335
rect	329	334	330	335
rect	330	334	331	335
rect	331	334	332	335
rect	347	334	348	335
rect	348	334	349	335
rect	350	334	351	335
rect	351	334	352	335
rect	352	334	353	335
rect	353	334	354	335
rect	354	334	355	335
rect	355	334	356	335
rect	356	334	357	335
rect	357	334	358	335
rect	132	336	133	337
rect	133	336	134	337
rect	135	336	136	337
rect	136	336	137	337
rect	138	336	139	337
rect	139	336	140	337
rect	141	336	142	337
rect	142	336	143	337
rect	143	336	144	337
rect	144	336	145	337
rect	145	336	146	337
rect	146	336	147	337
rect	148	336	149	337
rect	150	336	151	337
rect	151	336	152	337
rect	153	336	154	337
rect	154	336	155	337
rect	156	336	157	337
rect	157	336	158	337
rect	158	336	159	337
rect	159	336	160	337
rect	160	336	161	337
rect	161	336	162	337
rect	162	336	163	337
rect	163	336	164	337
rect	165	336	166	337
rect	166	336	167	337
rect	168	336	169	337
rect	169	336	170	337
rect	171	336	172	337
rect	172	336	173	337
rect	173	336	174	337
rect	175	336	176	337
rect	177	336	178	337
rect	178	336	179	337
rect	180	336	181	337
rect	181	336	182	337
rect	182	336	183	337
rect	183	336	184	337
rect	184	336	185	337
rect	186	336	187	337
rect	187	336	188	337
rect	189	336	190	337
rect	190	336	191	337
rect	191	336	192	337
rect	193	336	194	337
rect	194	336	195	337
rect	195	336	196	337
rect	196	336	197	337
rect	198	336	199	337
rect	199	336	200	337
rect	200	336	201	337
rect	202	336	203	337
rect	204	336	205	337
rect	205	336	206	337
rect	207	336	208	337
rect	208	336	209	337
rect	209	336	210	337
rect	210	336	211	337
rect	211	336	212	337
rect	212	336	213	337
rect	213	336	214	337
rect	214	336	215	337
rect	215	336	216	337
rect	216	336	217	337
rect	217	336	218	337
rect	219	336	220	337
rect	220	336	221	337
rect	222	336	223	337
rect	223	336	224	337
rect	225	336	226	337
rect	227	336	228	337
rect	228	336	229	337
rect	230	336	231	337
rect	231	336	232	337
rect	233	336	234	337
rect	234	336	235	337
rect	236	336	237	337
rect	237	336	238	337
rect	238	336	239	337
rect	239	336	240	337
rect	240	336	241	337
rect	241	336	242	337
rect	242	336	243	337
rect	243	336	244	337
rect	244	336	245	337
rect	245	336	246	337
rect	246	336	247	337
rect	248	336	249	337
rect	249	336	250	337
rect	250	336	251	337
rect	252	336	253	337
rect	253	336	254	337
rect	254	336	255	337
rect	255	336	256	337
rect	257	336	258	337
rect	258	336	259	337
rect	260	336	261	337
rect	261	336	262	337
rect	262	336	263	337
rect	263	336	264	337
rect	264	336	265	337
rect	265	336	266	337
rect	266	336	267	337
rect	267	336	268	337
rect	268	336	269	337
rect	269	336	270	337
rect	270	336	271	337
rect	271	336	272	337
rect	273	336	274	337
rect	274	336	275	337
rect	275	336	276	337
rect	276	336	277	337
rect	278	336	279	337
rect	279	336	280	337
rect	280	336	281	337
rect	281	336	282	337
rect	282	336	283	337
rect	283	336	284	337
rect	285	336	286	337
rect	286	336	287	337
rect	288	336	289	337
rect	289	336	290	337
rect	291	336	292	337
rect	292	336	293	337
rect	293	336	294	337
rect	294	336	295	337
rect	295	336	296	337
rect	296	336	297	337
rect	297	336	298	337
rect	298	336	299	337
rect	299	336	300	337
rect	300	336	301	337
rect	301	336	302	337
rect	302	336	303	337
rect	303	336	304	337
rect	304	336	305	337
rect	306	336	307	337
rect	307	336	308	337
rect	308	336	309	337
rect	309	336	310	337
rect	310	336	311	337
rect	311	336	312	337
rect	312	336	313	337
rect	313	336	314	337
rect	314	336	315	337
rect	315	336	316	337
rect	316	336	317	337
rect	317	336	318	337
rect	318	336	319	337
rect	319	336	320	337
rect	321	336	322	337
rect	322	336	323	337
rect	324	336	325	337
rect	325	336	326	337
rect	326	336	327	337
rect	327	336	328	337
rect	328	336	329	337
rect	329	336	330	337
rect	330	336	331	337
rect	331	336	332	337
rect	332	336	333	337
rect	359	336	360	337
rect	360	336	361	337
rect	362	336	363	337
rect	363	336	364	337
rect	364	336	365	337
rect	365	336	366	337
rect	366	336	367	337
rect	367	336	368	337
rect	368	336	369	337
rect	369	336	370	337
rect	371	336	372	337
rect	372	336	373	337
rect	373	336	374	337
rect	374	336	375	337
rect	375	336	376	337
rect	377	336	378	337
rect	378	336	379	337
rect	383	336	384	337
rect	384	336	385	337
rect	385	336	386	337
rect	386	336	387	337
rect	387	336	388	337
rect	84	338	85	339
rect	85	338	86	339
rect	86	338	87	339
rect	133	338	134	339
rect	135	338	136	339
rect	136	338	137	339
rect	138	338	139	339
rect	139	338	140	339
rect	141	338	142	339
rect	142	338	143	339
rect	143	338	144	339
rect	144	338	145	339
rect	145	338	146	339
rect	146	338	147	339
rect	148	338	149	339
rect	150	338	151	339
rect	151	338	152	339
rect	171	338	172	339
rect	172	338	173	339
rect	173	338	174	339
rect	175	338	176	339
rect	177	338	178	339
rect	178	338	179	339
rect	180	338	181	339
rect	181	338	182	339
rect	182	338	183	339
rect	196	338	197	339
rect	198	338	199	339
rect	199	338	200	339
rect	200	338	201	339
rect	202	338	203	339
rect	207	338	208	339
rect	208	338	209	339
rect	209	338	210	339
rect	217	338	218	339
rect	219	338	220	339
rect	220	338	221	339
rect	222	338	223	339
rect	223	338	224	339
rect	225	338	226	339
rect	227	338	228	339
rect	228	338	229	339
rect	230	338	231	339
rect	231	338	232	339
rect	233	338	234	339
rect	234	338	235	339
rect	236	338	237	339
rect	237	338	238	339
rect	238	338	239	339
rect	239	338	240	339
rect	240	338	241	339
rect	241	338	242	339
rect	242	338	243	339
rect	243	338	244	339
rect	244	338	245	339
rect	245	338	246	339
rect	246	338	247	339
rect	248	338	249	339
rect	249	338	250	339
rect	250	338	251	339
rect	252	338	253	339
rect	253	338	254	339
rect	254	338	255	339
rect	255	338	256	339
rect	257	338	258	339
rect	258	338	259	339
rect	260	338	261	339
rect	261	338	262	339
rect	262	338	263	339
rect	263	338	264	339
rect	264	338	265	339
rect	265	338	266	339
rect	266	338	267	339
rect	267	338	268	339
rect	268	338	269	339
rect	269	338	270	339
rect	270	338	271	339
rect	271	338	272	339
rect	273	338	274	339
rect	274	338	275	339
rect	275	338	276	339
rect	276	338	277	339
rect	278	338	279	339
rect	279	338	280	339
rect	280	338	281	339
rect	281	338	282	339
rect	282	338	283	339
rect	283	338	284	339
rect	285	338	286	339
rect	286	338	287	339
rect	288	338	289	339
rect	289	338	290	339
rect	291	338	292	339
rect	292	338	293	339
rect	293	338	294	339
rect	294	338	295	339
rect	295	338	296	339
rect	296	338	297	339
rect	297	338	298	339
rect	298	338	299	339
rect	299	338	300	339
rect	300	338	301	339
rect	301	338	302	339
rect	302	338	303	339
rect	303	338	304	339
rect	304	338	305	339
rect	306	338	307	339
rect	307	338	308	339
rect	308	338	309	339
rect	309	338	310	339
rect	310	338	311	339
rect	311	338	312	339
rect	312	338	313	339
rect	313	338	314	339
rect	314	338	315	339
rect	315	338	316	339
rect	316	338	317	339
rect	317	338	318	339
rect	318	338	319	339
rect	319	338	320	339
rect	321	338	322	339
rect	322	338	323	339
rect	324	338	325	339
rect	325	338	326	339
rect	326	338	327	339
rect	327	338	328	339
rect	328	338	329	339
rect	329	338	330	339
rect	330	338	331	339
rect	331	338	332	339
rect	332	338	333	339
rect	334	338	335	339
rect	336	338	337	339
rect	337	338	338	339
rect	339	338	340	339
rect	340	338	341	339
rect	341	338	342	339
rect	342	338	343	339
rect	343	338	344	339
rect	344	338	345	339
rect	345	338	346	339
rect	347	338	348	339
rect	348	338	349	339
rect	350	338	351	339
rect	351	338	352	339
rect	352	338	353	339
rect	353	338	354	339
rect	354	338	355	339
rect	355	338	356	339
rect	356	338	357	339
rect	357	338	358	339
rect	359	338	360	339
rect	360	338	361	339
rect	362	338	363	339
rect	363	338	364	339
rect	364	338	365	339
rect	365	338	366	339
rect	366	338	367	339
rect	367	338	368	339
rect	368	338	369	339
rect	369	338	370	339
rect	371	338	372	339
rect	372	338	373	339
rect	373	338	374	339
rect	374	338	375	339
rect	375	338	376	339
rect	377	338	378	339
rect	378	338	379	339
rect	379	338	380	339
rect	380	338	381	339
rect	381	338	382	339
rect	382	338	383	339
rect	383	338	384	339
rect	384	338	385	339
rect	385	338	386	339
rect	386	338	387	339
rect	387	338	388	339
rect	388	338	389	339
rect	389	338	390	339
rect	390	338	391	339
rect	392	338	393	339
rect	393	338	394	339
rect	395	338	396	339
rect	396	338	397	339
rect	397	338	398	339
rect	398	338	399	339
rect	399	338	400	339
rect	401	338	402	339
rect	402	338	403	339
rect	403	338	404	339
rect	404	338	405	339
rect	405	338	406	339
rect	406	338	407	339
rect	407	338	408	339
rect	408	338	409	339
rect	409	338	410	339
rect	81	340	82	341
rect	82	340	83	341
rect	83	340	84	341
rect	100	340	101	341
rect	102	340	103	341
rect	103	340	104	341
rect	145	340	146	341
rect	146	340	147	341
rect	148	340	149	341
rect	154	340	155	341
rect	172	340	173	341
rect	173	340	174	341
rect	175	340	176	341
rect	177	340	178	341
rect	178	340	179	341
rect	180	340	181	341
rect	181	340	182	341
rect	182	340	183	341
rect	184	340	185	341
rect	186	340	187	341
rect	187	340	188	341
rect	189	340	190	341
rect	190	340	191	341
rect	191	340	192	341
rect	193	340	194	341
rect	194	340	195	341
rect	196	340	197	341
rect	208	340	209	341
rect	209	340	210	341
rect	211	340	212	341
rect	212	340	213	341
rect	213	340	214	341
rect	214	340	215	341
rect	215	340	216	341
rect	217	340	218	341
rect	219	340	220	341
rect	220	340	221	341
rect	245	340	246	341
rect	246	340	247	341
rect	248	340	249	341
rect	249	340	250	341
rect	250	340	251	341
rect	269	340	270	341
rect	270	340	271	341
rect	271	340	272	341
rect	273	340	274	341
rect	274	340	275	341
rect	275	340	276	341
rect	276	340	277	341
rect	278	340	279	341
rect	279	340	280	341
rect	280	340	281	341
rect	281	340	282	341
rect	282	340	283	341
rect	283	340	284	341
rect	285	340	286	341
rect	286	340	287	341
rect	312	340	313	341
rect	313	340	314	341
rect	314	340	315	341
rect	315	340	316	341
rect	316	340	317	341
rect	317	340	318	341
rect	318	340	319	341
rect	319	340	320	341
rect	321	340	322	341
rect	322	340	323	341
rect	324	340	325	341
rect	325	340	326	341
rect	326	340	327	341
rect	327	340	328	341
rect	328	340	329	341
rect	329	340	330	341
rect	330	340	331	341
rect	331	340	332	341
rect	332	340	333	341
rect	334	340	335	341
rect	336	340	337	341
rect	337	340	338	341
rect	339	340	340	341
rect	340	340	341	341
rect	341	340	342	341
rect	342	340	343	341
rect	343	340	344	341
rect	344	340	345	341
rect	345	340	346	341
rect	347	340	348	341
rect	348	340	349	341
rect	350	340	351	341
rect	351	340	352	341
rect	352	340	353	341
rect	353	340	354	341
rect	354	340	355	341
rect	355	340	356	341
rect	356	340	357	341
rect	357	340	358	341
rect	359	340	360	341
rect	360	340	361	341
rect	362	340	363	341
rect	363	340	364	341
rect	364	340	365	341
rect	365	340	366	341
rect	366	340	367	341
rect	367	340	368	341
rect	368	340	369	341
rect	369	340	370	341
rect	371	340	372	341
rect	372	340	373	341
rect	373	340	374	341
rect	374	340	375	341
rect	375	340	376	341
rect	377	340	378	341
rect	378	340	379	341
rect	379	340	380	341
rect	380	340	381	341
rect	381	340	382	341
rect	73	342	74	343
rect	75	342	76	343
rect	76	342	77	343
rect	78	342	79	343
rect	79	342	80	343
rect	80	342	81	343
rect	81	342	82	343
rect	82	342	83	343
rect	83	342	84	343
rect	85	342	86	343
rect	86	342	87	343
rect	88	342	89	343
rect	89	342	90	343
rect	90	342	91	343
rect	91	342	92	343
rect	93	342	94	343
rect	94	342	95	343
rect	95	342	96	343
rect	96	342	97	343
rect	97	342	98	343
rect	98	342	99	343
rect	100	342	101	343
rect	106	342	107	343
rect	108	342	109	343
rect	109	342	110	343
rect	111	342	112	343
rect	112	342	113	343
rect	113	342	114	343
rect	115	342	116	343
rect	117	342	118	343
rect	118	342	119	343
rect	119	342	120	343
rect	120	342	121	343
rect	121	342	122	343
rect	135	342	136	343
rect	136	342	137	343
rect	138	342	139	343
rect	139	342	140	343
rect	141	342	142	343
rect	142	342	143	343
rect	143	342	144	343
rect	145	342	146	343
rect	146	342	147	343
rect	148	342	149	343
rect	149	342	150	343
rect	150	342	151	343
rect	151	342	152	343
rect	152	342	153	343
rect	154	342	155	343
rect	155	342	156	343
rect	156	342	157	343
rect	157	342	158	343
rect	158	342	159	343
rect	159	342	160	343
rect	160	342	161	343
rect	161	342	162	343
rect	162	342	163	343
rect	163	342	164	343
rect	165	342	166	343
rect	166	342	167	343
rect	168	342	169	343
rect	169	342	170	343
rect	170	342	171	343
rect	172	342	173	343
rect	173	342	174	343
rect	175	342	176	343
rect	177	342	178	343
rect	178	342	179	343
rect	180	342	181	343
rect	181	342	182	343
rect	182	342	183	343
rect	184	342	185	343
rect	186	342	187	343
rect	187	342	188	343
rect	189	342	190	343
rect	190	342	191	343
rect	191	342	192	343
rect	193	342	194	343
rect	194	342	195	343
rect	196	342	197	343
rect	197	342	198	343
rect	198	342	199	343
rect	199	342	200	343
rect	200	342	201	343
rect	202	342	203	343
rect	203	342	204	343
rect	204	342	205	343
rect	205	342	206	343
rect	206	342	207	343
rect	208	342	209	343
rect	209	342	210	343
rect	211	342	212	343
rect	212	342	213	343
rect	213	342	214	343
rect	214	342	215	343
rect	215	342	216	343
rect	217	342	218	343
rect	219	342	220	343
rect	220	342	221	343
rect	221	342	222	343
rect	222	342	223	343
rect	223	342	224	343
rect	225	342	226	343
rect	227	342	228	343
rect	228	342	229	343
rect	230	342	231	343
rect	231	342	232	343
rect	233	342	234	343
rect	234	342	235	343
rect	236	342	237	343
rect	237	342	238	343
rect	238	342	239	343
rect	239	342	240	343
rect	240	342	241	343
rect	241	342	242	343
rect	242	342	243	343
rect	243	342	244	343
rect	245	342	246	343
rect	246	342	247	343
rect	248	342	249	343
rect	249	342	250	343
rect	250	342	251	343
rect	251	342	252	343
rect	252	342	253	343
rect	253	342	254	343
rect	254	342	255	343
rect	255	342	256	343
rect	257	342	258	343
rect	258	342	259	343
rect	260	342	261	343
rect	261	342	262	343
rect	262	342	263	343
rect	263	342	264	343
rect	264	342	265	343
rect	265	342	266	343
rect	266	342	267	343
rect	267	342	268	343
rect	269	342	270	343
rect	270	342	271	343
rect	271	342	272	343
rect	273	342	274	343
rect	274	342	275	343
rect	275	342	276	343
rect	276	342	277	343
rect	278	342	279	343
rect	279	342	280	343
rect	280	342	281	343
rect	281	342	282	343
rect	282	342	283	343
rect	283	342	284	343
rect	285	342	286	343
rect	286	342	287	343
rect	287	342	288	343
rect	288	342	289	343
rect	289	342	290	343
rect	291	342	292	343
rect	292	342	293	343
rect	293	342	294	343
rect	294	342	295	343
rect	295	342	296	343
rect	296	342	297	343
rect	297	342	298	343
rect	298	342	299	343
rect	299	342	300	343
rect	300	342	301	343
rect	301	342	302	343
rect	302	342	303	343
rect	303	342	304	343
rect	304	342	305	343
rect	306	342	307	343
rect	307	342	308	343
rect	308	342	309	343
rect	309	342	310	343
rect	310	342	311	343
rect	312	342	313	343
rect	313	342	314	343
rect	314	342	315	343
rect	315	342	316	343
rect	316	342	317	343
rect	317	342	318	343
rect	318	342	319	343
rect	319	342	320	343
rect	321	342	322	343
rect	322	342	323	343
rect	324	342	325	343
rect	325	342	326	343
rect	326	342	327	343
rect	327	342	328	343
rect	328	342	329	343
rect	329	342	330	343
rect	330	342	331	343
rect	331	342	332	343
rect	332	342	333	343
rect	334	342	335	343
rect	336	342	337	343
rect	337	342	338	343
rect	339	342	340	343
rect	340	342	341	343
rect	341	342	342	343
rect	342	342	343	343
rect	343	342	344	343
rect	344	342	345	343
rect	345	342	346	343
rect	347	342	348	343
rect	348	342	349	343
rect	350	342	351	343
rect	351	342	352	343
rect	352	342	353	343
rect	353	342	354	343
rect	354	342	355	343
rect	355	342	356	343
rect	356	342	357	343
rect	357	342	358	343
rect	359	342	360	343
rect	360	342	361	343
rect	362	342	363	343
rect	363	342	364	343
rect	364	342	365	343
rect	365	342	366	343
rect	366	342	367	343
rect	367	342	368	343
rect	368	342	369	343
rect	369	342	370	343
rect	371	342	372	343
rect	372	342	373	343
rect	373	342	374	343
rect	374	342	375	343
rect	375	342	376	343
rect	377	342	378	343
rect	78	344	79	345
rect	79	344	80	345
rect	80	344	81	345
rect	103	344	104	345
rect	104	344	105	345
rect	106	344	107	345
rect	111	344	112	345
rect	112	344	113	345
rect	113	344	114	345
rect	115	344	116	345
rect	117	344	118	345
rect	118	344	119	345
rect	119	344	120	345
rect	120	344	121	345
rect	121	344	122	345
rect	122	344	123	345
rect	129	344	130	345
rect	130	344	131	345
rect	131	344	132	345
rect	133	344	134	345
rect	134	344	135	345
rect	151	344	152	345
rect	152	344	153	345
rect	154	344	155	345
rect	155	344	156	345
rect	156	344	157	345
rect	157	344	158	345
rect	158	344	159	345
rect	159	344	160	345
rect	160	344	161	345
rect	161	344	162	345
rect	162	344	163	345
rect	163	344	164	345
rect	165	344	166	345
rect	166	344	167	345
rect	168	344	169	345
rect	169	344	170	345
rect	170	344	171	345
rect	172	344	173	345
rect	173	344	174	345
rect	175	344	176	345
rect	205	344	206	345
rect	206	344	207	345
rect	208	344	209	345
rect	209	344	210	345
rect	211	344	212	345
rect	212	344	213	345
rect	213	344	214	345
rect	214	344	215	345
rect	215	344	216	345
rect	217	344	218	345
rect	225	344	226	345
rect	227	344	228	345
rect	228	344	229	345
rect	230	344	231	345
rect	231	344	232	345
rect	233	344	234	345
rect	234	344	235	345
rect	236	344	237	345
rect	237	344	238	345
rect	238	344	239	345
rect	239	344	240	345
rect	240	344	241	345
rect	241	344	242	345
rect	242	344	243	345
rect	243	344	244	345
rect	245	344	246	345
rect	246	344	247	345
rect	248	344	249	345
rect	249	344	250	345
rect	250	344	251	345
rect	251	344	252	345
rect	252	344	253	345
rect	253	344	254	345
rect	254	344	255	345
rect	255	344	256	345
rect	257	344	258	345
rect	258	344	259	345
rect	260	344	261	345
rect	261	344	262	345
rect	262	344	263	345
rect	263	344	264	345
rect	264	344	265	345
rect	265	344	266	345
rect	266	344	267	345
rect	267	344	268	345
rect	269	344	270	345
rect	270	344	271	345
rect	271	344	272	345
rect	273	344	274	345
rect	274	344	275	345
rect	275	344	276	345
rect	276	344	277	345
rect	278	344	279	345
rect	279	344	280	345
rect	280	344	281	345
rect	281	344	282	345
rect	282	344	283	345
rect	283	344	284	345
rect	285	344	286	345
rect	286	344	287	345
rect	287	344	288	345
rect	288	344	289	345
rect	289	344	290	345
rect	291	344	292	345
rect	292	344	293	345
rect	293	344	294	345
rect	294	344	295	345
rect	295	344	296	345
rect	296	344	297	345
rect	297	344	298	345
rect	298	344	299	345
rect	299	344	300	345
rect	300	344	301	345
rect	301	344	302	345
rect	302	344	303	345
rect	303	344	304	345
rect	304	344	305	345
rect	306	344	307	345
rect	307	344	308	345
rect	308	344	309	345
rect	309	344	310	345
rect	310	344	311	345
rect	312	344	313	345
rect	313	344	314	345
rect	314	344	315	345
rect	315	344	316	345
rect	316	344	317	345
rect	317	344	318	345
rect	318	344	319	345
rect	319	344	320	345
rect	321	344	322	345
rect	322	344	323	345
rect	324	344	325	345
rect	325	344	326	345
rect	326	344	327	345
rect	327	344	328	345
rect	328	344	329	345
rect	329	344	330	345
rect	330	344	331	345
rect	331	344	332	345
rect	332	344	333	345
rect	334	344	335	345
rect	336	344	337	345
rect	337	344	338	345
rect	339	344	340	345
rect	340	344	341	345
rect	341	344	342	345
rect	342	344	343	345
rect	48	346	49	347
rect	49	346	50	347
rect	50	346	51	347
rect	51	346	52	347
rect	52	346	53	347
rect	53	346	54	347
rect	66	346	67	347
rect	67	346	68	347
rect	68	346	69	347
rect	69	346	70	347
rect	70	346	71	347
rect	71	346	72	347
rect	73	346	74	347
rect	75	346	76	347
rect	76	346	77	347
rect	77	346	78	347
rect	97	346	98	347
rect	98	346	99	347
rect	100	346	101	347
rect	101	346	102	347
rect	103	346	104	347
rect	104	346	105	347
rect	106	346	107	347
rect	107	346	108	347
rect	108	346	109	347
rect	109	346	110	347
rect	110	346	111	347
rect	111	346	112	347
rect	112	346	113	347
rect	113	346	114	347
rect	115	346	116	347
rect	141	346	142	347
rect	142	346	143	347
rect	143	346	144	347
rect	145	346	146	347
rect	146	346	147	347
rect	148	346	149	347
rect	149	346	150	347
rect	151	346	152	347
rect	152	346	153	347
rect	154	346	155	347
rect	155	346	156	347
rect	199	346	200	347
rect	200	346	201	347
rect	202	346	203	347
rect	203	346	204	347
rect	205	346	206	347
rect	206	346	207	347
rect	208	346	209	347
rect	209	346	210	347
rect	211	346	212	347
rect	212	346	213	347
rect	213	346	214	347
rect	214	346	215	347
rect	215	346	216	347
rect	217	346	218	347
rect	218	346	219	347
rect	219	346	220	347
rect	220	346	221	347
rect	221	346	222	347
rect	222	346	223	347
rect	223	346	224	347
rect	224	346	225	347
rect	225	346	226	347
rect	227	346	228	347
rect	228	346	229	347
rect	230	346	231	347
rect	231	346	232	347
rect	233	346	234	347
rect	234	346	235	347
rect	236	346	237	347
rect	237	346	238	347
rect	238	346	239	347
rect	239	346	240	347
rect	240	346	241	347
rect	241	346	242	347
rect	242	346	243	347
rect	243	346	244	347
rect	245	346	246	347
rect	246	346	247	347
rect	248	346	249	347
rect	249	346	250	347
rect	250	346	251	347
rect	251	346	252	347
rect	252	346	253	347
rect	253	346	254	347
rect	254	346	255	347
rect	255	346	256	347
rect	257	346	258	347
rect	258	346	259	347
rect	260	346	261	347
rect	261	346	262	347
rect	262	346	263	347
rect	263	346	264	347
rect	264	346	265	347
rect	265	346	266	347
rect	266	346	267	347
rect	267	346	268	347
rect	269	346	270	347
rect	270	346	271	347
rect	271	346	272	347
rect	281	346	282	347
rect	282	346	283	347
rect	283	346	284	347
rect	309	346	310	347
rect	310	346	311	347
rect	312	346	313	347
rect	313	346	314	347
rect	314	346	315	347
rect	315	346	316	347
rect	316	346	317	347
rect	317	346	318	347
rect	318	346	319	347
rect	319	346	320	347
rect	321	346	322	347
rect	322	346	323	347
rect	324	346	325	347
rect	325	346	326	347
rect	326	346	327	347
rect	327	346	328	347
rect	328	346	329	347
rect	329	346	330	347
rect	330	346	331	347
rect	331	346	332	347
rect	332	346	333	347
rect	334	346	335	347
rect	8	348	9	349
rect	9	348	10	349
rect	10	348	11	349
rect	11	348	12	349
rect	12	348	13	349
rect	13	348	14	349
rect	45	348	46	349
rect	46	348	47	349
rect	47	348	48	349
rect	48	348	49	349
rect	49	348	50	349
rect	50	348	51	349
rect	57	348	58	349
rect	58	348	59	349
rect	59	348	60	349
rect	60	348	61	349
rect	61	348	62	349
rect	62	348	63	349
rect	93	348	94	349
rect	94	348	95	349
rect	95	348	96	349
rect	97	348	98	349
rect	98	348	99	349
rect	100	348	101	349
rect	101	348	102	349
rect	103	348	104	349
rect	104	348	105	349
rect	106	348	107	349
rect	107	348	108	349
rect	108	348	109	349
rect	109	348	110	349
rect	110	348	111	349
rect	111	348	112	349
rect	112	348	113	349
rect	113	348	114	349
rect	115	348	116	349
rect	116	348	117	349
rect	117	348	118	349
rect	118	348	119	349
rect	119	348	120	349
rect	120	348	121	349
rect	121	348	122	349
rect	122	348	123	349
rect	124	348	125	349
rect	125	348	126	349
rect	127	348	128	349
rect	128	348	129	349
rect	178	348	179	349
rect	179	348	180	349
rect	181	348	182	349
rect	182	348	183	349
rect	184	348	185	349
rect	189	348	190	349
rect	190	348	191	349
rect	191	348	192	349
rect	193	348	194	349
rect	194	348	195	349
rect	196	348	197	349
rect	197	348	198	349
rect	199	348	200	349
rect	200	348	201	349
rect	202	348	203	349
rect	203	348	204	349
rect	205	348	206	349
rect	206	348	207	349
rect	208	348	209	349
rect	209	348	210	349
rect	211	348	212	349
rect	212	348	213	349
rect	213	348	214	349
rect	214	348	215	349
rect	215	348	216	349
rect	217	348	218	349
rect	218	348	219	349
rect	219	348	220	349
rect	220	348	221	349
rect	221	348	222	349
rect	222	348	223	349
rect	223	348	224	349
rect	224	348	225	349
rect	225	348	226	349
rect	227	348	228	349
rect	228	348	229	349
rect	230	348	231	349
rect	231	348	232	349
rect	233	348	234	349
rect	234	348	235	349
rect	236	348	237	349
rect	237	348	238	349
rect	238	348	239	349
rect	239	348	240	349
rect	240	348	241	349
rect	241	348	242	349
rect	242	348	243	349
rect	243	348	244	349
rect	245	348	246	349
rect	246	348	247	349
rect	248	348	249	349
rect	249	348	250	349
rect	250	348	251	349
rect	251	348	252	349
rect	252	348	253	349
rect	253	348	254	349
rect	254	348	255	349
rect	255	348	256	349
rect	257	348	258	349
rect	258	348	259	349
rect	260	348	261	349
rect	261	348	262	349
rect	262	348	263	349
rect	263	348	264	349
rect	264	348	265	349
rect	265	348	266	349
rect	266	348	267	349
rect	267	348	268	349
rect	269	348	270	349
rect	270	348	271	349
rect	271	348	272	349
rect	272	348	273	349
rect	273	348	274	349
rect	274	348	275	349
rect	275	348	276	349
rect	276	348	277	349
rect	278	348	279	349
rect	279	348	280	349
rect	281	348	282	349
rect	282	348	283	349
rect	283	348	284	349
rect	284	348	285	349
rect	285	348	286	349
rect	286	348	287	349
rect	287	348	288	349
rect	288	348	289	349
rect	290	348	291	349
rect	291	348	292	349
rect	292	348	293	349
rect	293	348	294	349
rect	294	348	295	349
rect	295	348	296	349
rect	296	348	297	349
rect	297	348	298	349
rect	298	348	299	349
rect	299	348	300	349
rect	300	348	301	349
rect	301	348	302	349
rect	302	348	303	349
rect	303	348	304	349
rect	304	348	305	349
rect	306	348	307	349
rect	307	348	308	349
rect	309	348	310	349
rect	310	348	311	349
rect	312	348	313	349
rect	313	348	314	349
rect	314	348	315	349
rect	315	348	316	349
rect	316	348	317	349
rect	317	348	318	349
rect	318	348	319	349
rect	319	348	320	349
rect	321	348	322	349
rect	322	348	323	349
rect	324	348	325	349
rect	325	348	326	349
rect	326	348	327	349
rect	327	348	328	349
rect	328	348	329	349
rect	329	348	330	349
rect	330	348	331	349
rect	331	348	332	349
rect	332	348	333	349
rect	334	348	335	349
rect	335	348	336	349
rect	336	348	337	349
rect	337	348	338	349
rect	371	348	372	349
rect	372	348	373	349
rect	373	348	374	349
rect	374	348	375	349
rect	375	348	376	349
rect	392	348	393	349
rect	393	348	394	349
rect	394	348	395	349
rect	396	348	397	349
rect	397	348	398	349
rect	398	348	399	349
rect	399	348	400	349
rect	417	348	418	349
rect	418	348	419	349
rect	160	357	161	358
rect	161	357	162	358
rect	162	357	163	358
rect	163	357	164	358
rect	164	357	165	358
rect	157	359	158	360
rect	158	359	159	360
rect	159	359	160	360
rect	160	359	161	360
rect	161	359	162	360
rect	162	359	163	360
rect	163	359	164	360
rect	164	359	165	360
rect	165	359	166	360
rect	166	359	167	360
rect	167	359	168	360
rect	169	359	170	360
rect	170	359	171	360
rect	172	359	173	360
rect	173	359	174	360
rect	175	359	176	360
rect	176	359	177	360
rect	178	359	179	360
rect	179	359	180	360
rect	181	359	182	360
rect	182	359	183	360
rect	184	359	185	360
rect	185	359	186	360
rect	187	359	188	360
rect	188	359	189	360
rect	189	359	190	360
rect	190	359	191	360
rect	191	359	192	360
rect	193	359	194	360
rect	194	359	195	360
rect	196	359	197	360
rect	197	359	198	360
rect	198	359	199	360
rect	199	359	200	360
rect	200	359	201	360
rect	201	359	202	360
rect	202	359	203	360
rect	203	359	204	360
rect	205	359	206	360
rect	206	359	207	360
rect	208	359	209	360
rect	209	359	210	360
rect	211	359	212	360
rect	212	359	213	360
rect	214	359	215	360
rect	215	359	216	360
rect	216	359	217	360
rect	217	359	218	360
rect	218	359	219	360
rect	219	359	220	360
rect	220	359	221	360
rect	221	359	222	360
rect	222	359	223	360
rect	224	359	225	360
rect	225	359	226	360
rect	227	359	228	360
rect	228	359	229	360
rect	230	359	231	360
rect	231	359	232	360
rect	233	359	234	360
rect	234	359	235	360
rect	236	359	237	360
rect	237	359	238	360
rect	238	359	239	360
rect	239	359	240	360
rect	240	359	241	360
rect	241	359	242	360
rect	242	359	243	360
rect	243	359	244	360
rect	245	359	246	360
rect	246	359	247	360
rect	248	359	249	360
rect	249	359	250	360
rect	250	359	251	360
rect	251	359	252	360
rect	252	359	253	360
rect	253	359	254	360
rect	254	359	255	360
rect	255	359	256	360
rect	257	359	258	360
rect	258	359	259	360
rect	260	359	261	360
rect	261	359	262	360
rect	262	359	263	360
rect	263	359	264	360
rect	264	359	265	360
rect	265	359	266	360
rect	266	359	267	360
rect	267	359	268	360
rect	269	359	270	360
rect	270	359	271	360
rect	271	359	272	360
rect	272	359	273	360
rect	273	359	274	360
rect	92	361	93	362
rect	93	361	94	362
rect	94	361	95	362
rect	95	361	96	362
rect	97	361	98	362
rect	98	361	99	362
rect	119	361	120	362
rect	120	361	121	362
rect	121	361	122	362
rect	122	361	123	362
rect	124	361	125	362
rect	125	361	126	362
rect	126	361	127	362
rect	127	361	128	362
rect	128	361	129	362
rect	129	361	130	362
rect	130	361	131	362
rect	131	361	132	362
rect	158	361	159	362
rect	159	361	160	362
rect	160	361	161	362
rect	161	361	162	362
rect	162	361	163	362
rect	163	361	164	362
rect	164	361	165	362
rect	165	361	166	362
rect	166	361	167	362
rect	167	361	168	362
rect	169	361	170	362
rect	170	361	171	362
rect	172	361	173	362
rect	173	361	174	362
rect	175	361	176	362
rect	176	361	177	362
rect	178	361	179	362
rect	179	361	180	362
rect	181	361	182	362
rect	182	361	183	362
rect	79	363	80	364
rect	80	363	81	364
rect	82	363	83	364
rect	83	363	84	364
rect	85	363	86	364
rect	86	363	87	364
rect	88	363	89	364
rect	89	363	90	364
rect	90	363	91	364
rect	92	363	93	364
rect	93	363	94	364
rect	94	363	95	364
rect	95	363	96	364
rect	97	363	98	364
rect	98	363	99	364
rect	99	363	100	364
rect	100	363	101	364
rect	101	363	102	364
rect	103	363	104	364
rect	104	363	105	364
rect	106	363	107	364
rect	107	363	108	364
rect	108	363	109	364
rect	109	363	110	364
rect	110	363	111	364
rect	111	363	112	364
rect	112	363	113	364
rect	113	363	114	364
rect	115	363	116	364
rect	116	363	117	364
rect	117	363	118	364
rect	119	363	120	364
rect	120	363	121	364
rect	121	363	122	364
rect	122	363	123	364
rect	124	363	125	364
rect	125	363	126	364
rect	126	363	127	364
rect	127	363	128	364
rect	128	363	129	364
rect	129	363	130	364
rect	130	363	131	364
rect	131	363	132	364
rect	132	363	133	364
rect	133	363	134	364
rect	134	363	135	364
rect	136	363	137	364
rect	137	363	138	364
rect	139	363	140	364
rect	140	363	141	364
rect	141	363	142	364
rect	142	363	143	364
rect	143	363	144	364
rect	144	363	145	364
rect	145	363	146	364
rect	146	363	147	364
rect	148	363	149	364
rect	149	363	150	364
rect	151	363	152	364
rect	152	363	153	364
rect	154	363	155	364
rect	155	363	156	364
rect	156	363	157	364
rect	158	363	159	364
rect	159	363	160	364
rect	160	363	161	364
rect	161	363	162	364
rect	162	363	163	364
rect	163	363	164	364
rect	164	363	165	364
rect	165	363	166	364
rect	166	363	167	364
rect	167	363	168	364
rect	169	363	170	364
rect	170	363	171	364
rect	172	363	173	364
rect	173	363	174	364
rect	175	363	176	364
rect	176	363	177	364
rect	178	363	179	364
rect	179	363	180	364
rect	181	363	182	364
rect	182	363	183	364
rect	183	363	184	364
rect	184	363	185	364
rect	185	363	186	364
rect	187	363	188	364
rect	188	363	189	364
rect	189	363	190	364
rect	190	363	191	364
rect	191	363	192	364
rect	193	363	194	364
rect	194	363	195	364
rect	196	363	197	364
rect	197	363	198	364
rect	198	363	199	364
rect	199	363	200	364
rect	200	363	201	364
rect	201	363	202	364
rect	202	363	203	364
rect	203	363	204	364
rect	205	363	206	364
rect	206	363	207	364
rect	208	363	209	364
rect	209	363	210	364
rect	211	363	212	364
rect	212	363	213	364
rect	242	363	243	364
rect	243	363	244	364
rect	245	363	246	364
rect	246	363	247	364
rect	248	363	249	364
rect	249	363	250	364
rect	250	363	251	364
rect	251	363	252	364
rect	252	363	253	364
rect	253	363	254	364
rect	254	363	255	364
rect	255	363	256	364
rect	257	363	258	364
rect	258	363	259	364
rect	260	363	261	364
rect	261	363	262	364
rect	262	363	263	364
rect	263	363	264	364
rect	264	363	265	364
rect	265	363	266	364
rect	266	363	267	364
rect	267	363	268	364
rect	269	363	270	364
rect	270	363	271	364
rect	271	363	272	364
rect	272	363	273	364
rect	273	363	274	364
rect	275	363	276	364
rect	276	363	277	364
rect	278	363	279	364
rect	279	363	280	364
rect	296	363	297	364
rect	297	363	298	364
rect	298	363	299	364
rect	299	363	300	364
rect	300	363	301	364
rect	301	363	302	364
rect	302	363	303	364
rect	303	363	304	364
rect	304	363	305	364
rect	306	363	307	364
rect	307	363	308	364
rect	309	363	310	364
rect	310	363	311	364
rect	312	363	313	364
rect	313	363	314	364
rect	314	363	315	364
rect	315	363	316	364
rect	316	363	317	364
rect	317	363	318	364
rect	318	363	319	364
rect	319	363	320	364
rect	321	363	322	364
rect	322	363	323	364
rect	73	365	74	366
rect	74	365	75	366
rect	76	365	77	366
rect	77	365	78	366
rect	78	365	79	366
rect	85	365	86	366
rect	86	365	87	366
rect	88	365	89	366
rect	89	365	90	366
rect	90	365	91	366
rect	92	365	93	366
rect	93	365	94	366
rect	134	365	135	366
rect	136	365	137	366
rect	137	365	138	366
rect	139	365	140	366
rect	140	365	141	366
rect	141	365	142	366
rect	142	365	143	366
rect	143	365	144	366
rect	144	365	145	366
rect	145	365	146	366
rect	146	365	147	366
rect	148	365	149	366
rect	149	365	150	366
rect	151	365	152	366
rect	152	365	153	366
rect	154	365	155	366
rect	155	365	156	366
rect	156	365	157	366
rect	158	365	159	366
rect	159	365	160	366
rect	160	365	161	366
rect	161	365	162	366
rect	162	365	163	366
rect	163	365	164	366
rect	164	365	165	366
rect	165	365	166	366
rect	166	365	167	366
rect	167	365	168	366
rect	190	365	191	366
rect	191	365	192	366
rect	193	365	194	366
rect	194	365	195	366
rect	196	365	197	366
rect	197	365	198	366
rect	198	365	199	366
rect	199	365	200	366
rect	200	365	201	366
rect	201	365	202	366
rect	202	365	203	366
rect	203	365	204	366
rect	205	365	206	366
rect	206	365	207	366
rect	208	365	209	366
rect	209	365	210	366
rect	211	365	212	366
rect	212	365	213	366
rect	213	365	214	366
rect	214	365	215	366
rect	215	365	216	366
rect	216	365	217	366
rect	217	365	218	366
rect	218	365	219	366
rect	219	365	220	366
rect	220	365	221	366
rect	221	365	222	366
rect	222	365	223	366
rect	224	365	225	366
rect	225	365	226	366
rect	227	365	228	366
rect	228	365	229	366
rect	230	365	231	366
rect	231	365	232	366
rect	233	365	234	366
rect	234	365	235	366
rect	236	365	237	366
rect	237	365	238	366
rect	238	365	239	366
rect	239	365	240	366
rect	240	365	241	366
rect	242	365	243	366
rect	243	365	244	366
rect	284	365	285	366
rect	285	365	286	366
rect	286	365	287	366
rect	287	365	288	366
rect	288	365	289	366
rect	290	365	291	366
rect	291	365	292	366
rect	292	365	293	366
rect	293	365	294	366
rect	294	365	295	366
rect	296	365	297	366
rect	297	365	298	366
rect	298	365	299	366
rect	299	365	300	366
rect	300	365	301	366
rect	301	365	302	366
rect	302	365	303	366
rect	303	365	304	366
rect	304	365	305	366
rect	306	365	307	366
rect	307	365	308	366
rect	309	365	310	366
rect	310	365	311	366
rect	74	367	75	368
rect	82	367	83	368
rect	83	367	84	368
rect	84	367	85	368
rect	85	367	86	368
rect	86	367	87	368
rect	88	367	89	368
rect	89	367	90	368
rect	90	367	91	368
rect	92	367	93	368
rect	93	367	94	368
rect	95	367	96	368
rect	97	367	98	368
rect	98	367	99	368
rect	99	367	100	368
rect	100	367	101	368
rect	101	367	102	368
rect	103	367	104	368
rect	104	367	105	368
rect	106	367	107	368
rect	107	367	108	368
rect	108	367	109	368
rect	109	367	110	368
rect	110	367	111	368
rect	111	367	112	368
rect	112	367	113	368
rect	113	367	114	368
rect	115	367	116	368
rect	116	367	117	368
rect	117	367	118	368
rect	119	367	120	368
rect	120	367	121	368
rect	121	367	122	368
rect	122	367	123	368
rect	124	367	125	368
rect	125	367	126	368
rect	126	367	127	368
rect	127	367	128	368
rect	128	367	129	368
rect	129	367	130	368
rect	130	367	131	368
rect	131	367	132	368
rect	132	367	133	368
rect	134	367	135	368
rect	136	367	137	368
rect	137	367	138	368
rect	139	367	140	368
rect	140	367	141	368
rect	141	367	142	368
rect	142	367	143	368
rect	143	367	144	368
rect	144	367	145	368
rect	145	367	146	368
rect	146	367	147	368
rect	148	367	149	368
rect	149	367	150	368
rect	151	367	152	368
rect	152	367	153	368
rect	154	367	155	368
rect	155	367	156	368
rect	156	367	157	368
rect	158	367	159	368
rect	159	367	160	368
rect	160	367	161	368
rect	161	367	162	368
rect	162	367	163	368
rect	163	367	164	368
rect	164	367	165	368
rect	165	367	166	368
rect	166	367	167	368
rect	167	367	168	368
rect	168	367	169	368
rect	169	367	170	368
rect	170	367	171	368
rect	172	367	173	368
rect	173	367	174	368
rect	175	367	176	368
rect	176	367	177	368
rect	178	367	179	368
rect	179	367	180	368
rect	181	367	182	368
rect	182	367	183	368
rect	183	367	184	368
rect	184	367	185	368
rect	185	367	186	368
rect	187	367	188	368
rect	188	367	189	368
rect	190	367	191	368
rect	191	367	192	368
rect	193	367	194	368
rect	194	367	195	368
rect	196	367	197	368
rect	197	367	198	368
rect	198	367	199	368
rect	199	367	200	368
rect	200	367	201	368
rect	201	367	202	368
rect	202	367	203	368
rect	203	367	204	368
rect	205	367	206	368
rect	206	367	207	368
rect	208	367	209	368
rect	209	367	210	368
rect	211	367	212	368
rect	212	367	213	368
rect	213	367	214	368
rect	214	367	215	368
rect	215	367	216	368
rect	216	367	217	368
rect	217	367	218	368
rect	218	367	219	368
rect	219	367	220	368
rect	220	367	221	368
rect	221	367	222	368
rect	222	367	223	368
rect	224	367	225	368
rect	225	367	226	368
rect	227	367	228	368
rect	228	367	229	368
rect	230	367	231	368
rect	231	367	232	368
rect	233	367	234	368
rect	234	367	235	368
rect	236	367	237	368
rect	237	367	238	368
rect	238	367	239	368
rect	239	367	240	368
rect	240	367	241	368
rect	242	367	243	368
rect	243	367	244	368
rect	244	367	245	368
rect	245	367	246	368
rect	246	367	247	368
rect	248	367	249	368
rect	249	367	250	368
rect	250	367	251	368
rect	251	367	252	368
rect	252	367	253	368
rect	253	367	254	368
rect	254	367	255	368
rect	255	367	256	368
rect	257	367	258	368
rect	258	367	259	368
rect	260	367	261	368
rect	261	367	262	368
rect	262	367	263	368
rect	263	367	264	368
rect	264	367	265	368
rect	265	367	266	368
rect	266	367	267	368
rect	267	367	268	368
rect	269	367	270	368
rect	270	367	271	368
rect	271	367	272	368
rect	272	367	273	368
rect	273	367	274	368
rect	275	367	276	368
rect	276	367	277	368
rect	278	367	279	368
rect	279	367	280	368
rect	280	367	281	368
rect	281	367	282	368
rect	282	367	283	368
rect	284	367	285	368
rect	285	367	286	368
rect	286	367	287	368
rect	287	367	288	368
rect	288	367	289	368
rect	290	367	291	368
rect	291	367	292	368
rect	292	367	293	368
rect	293	367	294	368
rect	294	367	295	368
rect	296	367	297	368
rect	297	367	298	368
rect	298	367	299	368
rect	299	367	300	368
rect	300	367	301	368
rect	301	367	302	368
rect	302	367	303	368
rect	303	367	304	368
rect	304	367	305	368
rect	306	367	307	368
rect	307	367	308	368
rect	309	367	310	368
rect	310	367	311	368
rect	311	367	312	368
rect	312	367	313	368
rect	313	367	314	368
rect	314	367	315	368
rect	315	367	316	368
rect	316	367	317	368
rect	317	367	318	368
rect	318	367	319	368
rect	319	367	320	368
rect	321	367	322	368
rect	322	367	323	368
rect	323	367	324	368
rect	324	367	325	368
rect	325	367	326	368
rect	77	369	78	370
rect	78	369	79	370
rect	80	369	81	370
rect	81	369	82	370
rect	82	369	83	370
rect	83	369	84	370
rect	84	369	85	370
rect	85	369	86	370
rect	86	369	87	370
rect	88	369	89	370
rect	89	369	90	370
rect	90	369	91	370
rect	92	369	93	370
rect	93	369	94	370
rect	95	369	96	370
rect	97	369	98	370
rect	98	369	99	370
rect	99	369	100	370
rect	100	369	101	370
rect	101	369	102	370
rect	103	369	104	370
rect	104	369	105	370
rect	131	369	132	370
rect	132	369	133	370
rect	134	369	135	370
rect	136	369	137	370
rect	137	369	138	370
rect	139	369	140	370
rect	140	369	141	370
rect	141	369	142	370
rect	142	369	143	370
rect	143	369	144	370
rect	144	369	145	370
rect	145	369	146	370
rect	146	369	147	370
rect	148	369	149	370
rect	149	369	150	370
rect	154	369	155	370
rect	155	369	156	370
rect	156	369	157	370
rect	158	369	159	370
rect	159	369	160	370
rect	160	369	161	370
rect	161	369	162	370
rect	162	369	163	370
rect	163	369	164	370
rect	168	369	169	370
rect	169	369	170	370
rect	170	369	171	370
rect	172	369	173	370
rect	173	369	174	370
rect	175	369	176	370
rect	176	369	177	370
rect	178	369	179	370
rect	179	369	180	370
rect	181	369	182	370
rect	182	369	183	370
rect	183	369	184	370
rect	184	369	185	370
rect	185	369	186	370
rect	187	369	188	370
rect	188	369	189	370
rect	190	369	191	370
rect	191	369	192	370
rect	193	369	194	370
rect	194	369	195	370
rect	281	369	282	370
rect	282	369	283	370
rect	284	369	285	370
rect	285	369	286	370
rect	286	369	287	370
rect	287	369	288	370
rect	288	369	289	370
rect	290	369	291	370
rect	291	369	292	370
rect	292	369	293	370
rect	293	369	294	370
rect	294	369	295	370
rect	296	369	297	370
rect	297	369	298	370
rect	298	369	299	370
rect	299	369	300	370
rect	300	369	301	370
rect	301	369	302	370
rect	302	369	303	370
rect	303	369	304	370
rect	304	369	305	370
rect	306	369	307	370
rect	307	369	308	370
rect	309	369	310	370
rect	310	369	311	370
rect	311	369	312	370
rect	312	369	313	370
rect	313	369	314	370
rect	314	369	315	370
rect	315	369	316	370
rect	316	369	317	370
rect	317	369	318	370
rect	318	369	319	370
rect	319	369	320	370
rect	324	369	325	370
rect	325	369	326	370
rect	326	369	327	370
rect	327	369	328	370
rect	328	369	329	370
rect	329	369	330	370
rect	330	369	331	370
rect	331	369	332	370
rect	332	369	333	370
rect	333	369	334	370
rect	334	369	335	370
rect	335	369	336	370
rect	336	369	337	370
rect	337	369	338	370
rect	338	369	339	370
rect	339	369	340	370
rect	340	369	341	370
rect	341	369	342	370
rect	342	369	343	370
rect	343	369	344	370
rect	344	369	345	370
rect	345	369	346	370
rect	347	369	348	370
rect	348	369	349	370
rect	71	371	72	372
rect	72	371	73	372
rect	74	371	75	372
rect	75	371	76	372
rect	77	371	78	372
rect	78	371	79	372
rect	80	371	81	372
rect	81	371	82	372
rect	82	371	83	372
rect	83	371	84	372
rect	84	371	85	372
rect	85	371	86	372
rect	86	371	87	372
rect	88	371	89	372
rect	89	371	90	372
rect	90	371	91	372
rect	92	371	93	372
rect	93	371	94	372
rect	95	371	96	372
rect	97	371	98	372
rect	98	371	99	372
rect	99	371	100	372
rect	100	371	101	372
rect	101	371	102	372
rect	146	371	147	372
rect	152	371	153	372
rect	153	371	154	372
rect	154	371	155	372
rect	155	371	156	372
rect	156	371	157	372
rect	158	371	159	372
rect	159	371	160	372
rect	160	371	161	372
rect	161	371	162	372
rect	162	371	163	372
rect	163	371	164	372
rect	165	371	166	372
rect	166	371	167	372
rect	168	371	169	372
rect	169	371	170	372
rect	170	371	171	372
rect	187	371	188	372
rect	188	371	189	372
rect	190	371	191	372
rect	191	371	192	372
rect	202	371	203	372
rect	203	371	204	372
rect	205	371	206	372
rect	206	371	207	372
rect	208	371	209	372
rect	209	371	210	372
rect	221	371	222	372
rect	222	371	223	372
rect	224	371	225	372
rect	225	371	226	372
rect	227	371	228	372
rect	228	371	229	372
rect	230	371	231	372
rect	231	371	232	372
rect	245	371	246	372
rect	246	371	247	372
rect	248	371	249	372
rect	249	371	250	372
rect	250	371	251	372
rect	251	371	252	372
rect	252	371	253	372
rect	253	371	254	372
rect	254	371	255	372
rect	255	371	256	372
rect	257	371	258	372
rect	258	371	259	372
rect	260	371	261	372
rect	261	371	262	372
rect	262	371	263	372
rect	263	371	264	372
rect	264	371	265	372
rect	265	371	266	372
rect	266	371	267	372
rect	267	371	268	372
rect	272	371	273	372
rect	273	371	274	372
rect	275	371	276	372
rect	276	371	277	372
rect	278	371	279	372
rect	279	371	280	372
rect	281	371	282	372
rect	282	371	283	372
rect	284	371	285	372
rect	285	371	286	372
rect	286	371	287	372
rect	287	371	288	372
rect	288	371	289	372
rect	290	371	291	372
rect	291	371	292	372
rect	292	371	293	372
rect	293	371	294	372
rect	294	371	295	372
rect	296	371	297	372
rect	297	371	298	372
rect	298	371	299	372
rect	299	371	300	372
rect	300	371	301	372
rect	301	371	302	372
rect	302	371	303	372
rect	303	371	304	372
rect	304	371	305	372
rect	306	371	307	372
rect	307	371	308	372
rect	309	371	310	372
rect	310	371	311	372
rect	311	371	312	372
rect	312	371	313	372
rect	313	371	314	372
rect	314	371	315	372
rect	315	371	316	372
rect	316	371	317	372
rect	317	371	318	372
rect	318	371	319	372
rect	319	371	320	372
rect	320	371	321	372
rect	321	371	322	372
rect	322	371	323	372
rect	324	371	325	372
rect	325	371	326	372
rect	349	371	350	372
rect	350	371	351	372
rect	351	371	352	372
rect	352	371	353	372
rect	353	371	354	372
rect	354	371	355	372
rect	355	371	356	372
rect	356	371	357	372
rect	357	371	358	372
rect	5	373	6	374
rect	6	373	7	374
rect	8	373	9	374
rect	9	373	10	374
rect	11	373	12	374
rect	12	373	13	374
rect	13	373	14	374
rect	14	373	15	374
rect	15	373	16	374
rect	16	373	17	374
rect	17	373	18	374
rect	18	373	19	374
rect	19	373	20	374
rect	68	373	69	374
rect	69	373	70	374
rect	71	373	72	374
rect	72	373	73	374
rect	74	373	75	374
rect	75	373	76	374
rect	77	373	78	374
rect	78	373	79	374
rect	80	373	81	374
rect	81	373	82	374
rect	82	373	83	374
rect	83	373	84	374
rect	84	373	85	374
rect	85	373	86	374
rect	86	373	87	374
rect	88	373	89	374
rect	89	373	90	374
rect	90	373	91	374
rect	92	373	93	374
rect	93	373	94	374
rect	95	373	96	374
rect	107	373	108	374
rect	108	373	109	374
rect	109	373	110	374
rect	110	373	111	374
rect	111	373	112	374
rect	112	373	113	374
rect	113	373	114	374
rect	122	373	123	374
rect	124	373	125	374
rect	125	373	126	374
rect	126	373	127	374
rect	127	373	128	374
rect	128	373	129	374
rect	129	373	130	374
rect	131	373	132	374
rect	132	373	133	374
rect	134	373	135	374
rect	149	373	150	374
rect	150	373	151	374
rect	152	373	153	374
rect	153	373	154	374
rect	154	373	155	374
rect	155	373	156	374
rect	156	373	157	374
rect	158	373	159	374
rect	159	373	160	374
rect	160	373	161	374
rect	161	373	162	374
rect	162	373	163	374
rect	163	373	164	374
rect	165	373	166	374
rect	166	373	167	374
rect	168	373	169	374
rect	169	373	170	374
rect	170	373	171	374
rect	171	373	172	374
rect	172	373	173	374
rect	173	373	174	374
rect	175	373	176	374
rect	176	373	177	374
rect	178	373	179	374
rect	179	373	180	374
rect	193	373	194	374
rect	194	373	195	374
rect	195	373	196	374
rect	196	373	197	374
rect	197	373	198	374
rect	198	373	199	374
rect	199	373	200	374
rect	200	373	201	374
rect	202	373	203	374
rect	203	373	204	374
rect	205	373	206	374
rect	206	373	207	374
rect	218	373	219	374
rect	219	373	220	374
rect	221	373	222	374
rect	222	373	223	374
rect	224	373	225	374
rect	225	373	226	374
rect	227	373	228	374
rect	228	373	229	374
rect	233	373	234	374
rect	234	373	235	374
rect	236	373	237	374
rect	237	373	238	374
rect	238	373	239	374
rect	239	373	240	374
rect	240	373	241	374
rect	242	373	243	374
rect	243	373	244	374
rect	245	373	246	374
rect	246	373	247	374
rect	254	373	255	374
rect	255	373	256	374
rect	269	373	270	374
rect	270	373	271	374
rect	272	373	273	374
rect	273	373	274	374
rect	275	373	276	374
rect	276	373	277	374
rect	278	373	279	374
rect	279	373	280	374
rect	281	373	282	374
rect	282	373	283	374
rect	284	373	285	374
rect	285	373	286	374
rect	286	373	287	374
rect	287	373	288	374
rect	288	373	289	374
rect	290	373	291	374
rect	291	373	292	374
rect	292	373	293	374
rect	293	373	294	374
rect	294	373	295	374
rect	296	373	297	374
rect	297	373	298	374
rect	298	373	299	374
rect	299	373	300	374
rect	300	373	301	374
rect	301	373	302	374
rect	302	373	303	374
rect	303	373	304	374
rect	304	373	305	374
rect	306	373	307	374
rect	307	373	308	374
rect	333	373	334	374
rect	334	373	335	374
rect	335	373	336	374
rect	336	373	337	374
rect	337	373	338	374
rect	338	373	339	374
rect	339	373	340	374
rect	340	373	341	374
rect	341	373	342	374
rect	342	373	343	374
rect	343	373	344	374
rect	344	373	345	374
rect	345	373	346	374
rect	347	373	348	374
rect	349	373	350	374
rect	350	373	351	374
rect	351	373	352	374
rect	352	373	353	374
rect	353	373	354	374
rect	354	373	355	374
rect	355	373	356	374
rect	356	373	357	374
rect	357	373	358	374
rect	358	373	359	374
rect	359	373	360	374
rect	360	373	361	374
rect	361	373	362	374
rect	362	373	363	374
rect	363	373	364	374
rect	364	373	365	374
rect	365	373	366	374
rect	366	373	367	374
rect	367	373	368	374
rect	368	373	369	374
rect	369	373	370	374
rect	370	373	371	374
rect	372	373	373	374
rect	373	373	374	374
rect	374	373	375	374
rect	5	375	6	376
rect	6	375	7	376
rect	55	375	56	376
rect	56	375	57	376
rect	57	375	58	376
rect	58	375	59	376
rect	59	375	60	376
rect	60	375	61	376
rect	61	375	62	376
rect	62	375	63	376
rect	64	375	65	376
rect	65	375	66	376
rect	66	375	67	376
rect	68	375	69	376
rect	69	375	70	376
rect	71	375	72	376
rect	72	375	73	376
rect	74	375	75	376
rect	75	375	76	376
rect	77	375	78	376
rect	78	375	79	376
rect	80	375	81	376
rect	81	375	82	376
rect	82	375	83	376
rect	83	375	84	376
rect	84	375	85	376
rect	85	375	86	376
rect	86	375	87	376
rect	88	375	89	376
rect	89	375	90	376
rect	90	375	91	376
rect	92	375	93	376
rect	93	375	94	376
rect	95	375	96	376
rect	96	375	97	376
rect	97	375	98	376
rect	98	375	99	376
rect	99	375	100	376
rect	100	375	101	376
rect	101	375	102	376
rect	102	375	103	376
rect	103	375	104	376
rect	104	375	105	376
rect	105	375	106	376
rect	107	375	108	376
rect	108	375	109	376
rect	109	375	110	376
rect	110	375	111	376
rect	111	375	112	376
rect	112	375	113	376
rect	113	375	114	376
rect	114	375	115	376
rect	115	375	116	376
rect	116	375	117	376
rect	117	375	118	376
rect	119	375	120	376
rect	120	375	121	376
rect	122	375	123	376
rect	124	375	125	376
rect	125	375	126	376
rect	126	375	127	376
rect	127	375	128	376
rect	128	375	129	376
rect	129	375	130	376
rect	131	375	132	376
rect	132	375	133	376
rect	134	375	135	376
rect	135	375	136	376
rect	136	375	137	376
rect	137	375	138	376
rect	139	375	140	376
rect	140	375	141	376
rect	141	375	142	376
rect	142	375	143	376
rect	143	375	144	376
rect	144	375	145	376
rect	146	375	147	376
rect	147	375	148	376
rect	149	375	150	376
rect	150	375	151	376
rect	152	375	153	376
rect	153	375	154	376
rect	154	375	155	376
rect	155	375	156	376
rect	156	375	157	376
rect	158	375	159	376
rect	159	375	160	376
rect	160	375	161	376
rect	161	375	162	376
rect	162	375	163	376
rect	163	375	164	376
rect	165	375	166	376
rect	166	375	167	376
rect	168	375	169	376
rect	169	375	170	376
rect	170	375	171	376
rect	171	375	172	376
rect	172	375	173	376
rect	173	375	174	376
rect	175	375	176	376
rect	176	375	177	376
rect	178	375	179	376
rect	179	375	180	376
rect	180	375	181	376
rect	181	375	182	376
rect	182	375	183	376
rect	183	375	184	376
rect	184	375	185	376
rect	185	375	186	376
rect	186	375	187	376
rect	187	375	188	376
rect	188	375	189	376
rect	190	375	191	376
rect	191	375	192	376
rect	193	375	194	376
rect	194	375	195	376
rect	195	375	196	376
rect	196	375	197	376
rect	197	375	198	376
rect	198	375	199	376
rect	199	375	200	376
rect	200	375	201	376
rect	202	375	203	376
rect	203	375	204	376
rect	205	375	206	376
rect	206	375	207	376
rect	207	375	208	376
rect	208	375	209	376
rect	209	375	210	376
rect	210	375	211	376
rect	211	375	212	376
rect	212	375	213	376
rect	213	375	214	376
rect	214	375	215	376
rect	215	375	216	376
rect	216	375	217	376
rect	218	375	219	376
rect	219	375	220	376
rect	221	375	222	376
rect	222	375	223	376
rect	224	375	225	376
rect	225	375	226	376
rect	227	375	228	376
rect	228	375	229	376
rect	229	375	230	376
rect	230	375	231	376
rect	231	375	232	376
rect	233	375	234	376
rect	234	375	235	376
rect	236	375	237	376
rect	237	375	238	376
rect	238	375	239	376
rect	239	375	240	376
rect	240	375	241	376
rect	242	375	243	376
rect	243	375	244	376
rect	245	375	246	376
rect	246	375	247	376
rect	247	375	248	376
rect	248	375	249	376
rect	249	375	250	376
rect	250	375	251	376
rect	251	375	252	376
rect	252	375	253	376
rect	254	375	255	376
rect	255	375	256	376
rect	256	375	257	376
rect	257	375	258	376
rect	258	375	259	376
rect	260	375	261	376
rect	261	375	262	376
rect	262	375	263	376
rect	263	375	264	376
rect	264	375	265	376
rect	265	375	266	376
rect	266	375	267	376
rect	267	375	268	376
rect	269	375	270	376
rect	270	375	271	376
rect	272	375	273	376
rect	273	375	274	376
rect	275	375	276	376
rect	276	375	277	376
rect	278	375	279	376
rect	279	375	280	376
rect	281	375	282	376
rect	282	375	283	376
rect	284	375	285	376
rect	285	375	286	376
rect	286	375	287	376
rect	287	375	288	376
rect	288	375	289	376
rect	290	375	291	376
rect	291	375	292	376
rect	292	375	293	376
rect	293	375	294	376
rect	294	375	295	376
rect	296	375	297	376
rect	297	375	298	376
rect	298	375	299	376
rect	299	375	300	376
rect	300	375	301	376
rect	301	375	302	376
rect	302	375	303	376
rect	303	375	304	376
rect	304	375	305	376
rect	306	375	307	376
rect	307	375	308	376
rect	308	375	309	376
rect	309	375	310	376
rect	310	375	311	376
rect	311	375	312	376
rect	312	375	313	376
rect	313	375	314	376
rect	314	375	315	376
rect	315	375	316	376
rect	316	375	317	376
rect	317	375	318	376
rect	318	375	319	376
rect	319	375	320	376
rect	320	375	321	376
rect	321	375	322	376
rect	322	375	323	376
rect	324	375	325	376
rect	325	375	326	376
rect	327	375	328	376
rect	328	375	329	376
rect	329	375	330	376
rect	330	375	331	376
rect	331	375	332	376
rect	333	375	334	376
rect	334	375	335	376
rect	335	375	336	376
rect	336	375	337	376
rect	337	375	338	376
rect	338	375	339	376
rect	339	375	340	376
rect	340	375	341	376
rect	341	375	342	376
rect	342	375	343	376
rect	343	375	344	376
rect	344	375	345	376
rect	345	375	346	376
rect	347	375	348	376
rect	349	375	350	376
rect	350	375	351	376
rect	365	375	366	376
rect	366	375	367	376
rect	367	375	368	376
rect	368	375	369	376
rect	369	375	370	376
rect	370	375	371	376
rect	372	375	373	376
rect	373	375	374	376
rect	374	375	375	376
rect	375	375	376	376
rect	376	375	377	376
rect	377	375	378	376
rect	378	375	379	376
rect	379	375	380	376
rect	380	375	381	376
rect	381	375	382	376
rect	382	375	383	376
rect	383	375	384	376
rect	384	375	385	376
rect	385	375	386	376
rect	386	375	387	376
rect	387	375	388	376
rect	388	375	389	376
rect	389	375	390	376
rect	390	375	391	376
rect	391	375	392	376
rect	393	375	394	376
rect	394	375	395	376
rect	9	377	10	378
rect	11	377	12	378
rect	12	377	13	378
rect	13	377	14	378
rect	14	377	15	378
rect	15	377	16	378
rect	16	377	17	378
rect	17	377	18	378
rect	18	377	19	378
rect	19	377	20	378
rect	20	377	21	378
rect	21	377	22	378
rect	22	377	23	378
rect	23	377	24	378
rect	24	377	25	378
rect	25	377	26	378
rect	26	377	27	378
rect	27	377	28	378
rect	28	377	29	378
rect	29	377	30	378
rect	30	377	31	378
rect	31	377	32	378
rect	32	377	33	378
rect	33	377	34	378
rect	34	377	35	378
rect	35	377	36	378
rect	36	377	37	378
rect	37	377	38	378
rect	38	377	39	378
rect	39	377	40	378
rect	40	377	41	378
rect	41	377	42	378
rect	42	377	43	378
rect	43	377	44	378
rect	44	377	45	378
rect	45	377	46	378
rect	46	377	47	378
rect	47	377	48	378
rect	48	377	49	378
rect	49	377	50	378
rect	50	377	51	378
rect	52	377	53	378
rect	53	377	54	378
rect	54	377	55	378
rect	55	377	56	378
rect	56	377	57	378
rect	57	377	58	378
rect	58	377	59	378
rect	59	377	60	378
rect	60	377	61	378
rect	61	377	62	378
rect	62	377	63	378
rect	64	377	65	378
rect	65	377	66	378
rect	66	377	67	378
rect	68	377	69	378
rect	69	377	70	378
rect	71	377	72	378
rect	72	377	73	378
rect	74	377	75	378
rect	75	377	76	378
rect	77	377	78	378
rect	78	377	79	378
rect	80	377	81	378
rect	81	377	82	378
rect	82	377	83	378
rect	83	377	84	378
rect	84	377	85	378
rect	85	377	86	378
rect	86	377	87	378
rect	88	377	89	378
rect	89	377	90	378
rect	90	377	91	378
rect	92	377	93	378
rect	93	377	94	378
rect	95	377	96	378
rect	96	377	97	378
rect	97	377	98	378
rect	98	377	99	378
rect	99	377	100	378
rect	100	377	101	378
rect	101	377	102	378
rect	102	377	103	378
rect	103	377	104	378
rect	104	377	105	378
rect	105	377	106	378
rect	107	377	108	378
rect	108	377	109	378
rect	109	377	110	378
rect	110	377	111	378
rect	111	377	112	378
rect	112	377	113	378
rect	113	377	114	378
rect	114	377	115	378
rect	115	377	116	378
rect	116	377	117	378
rect	117	377	118	378
rect	119	377	120	378
rect	120	377	121	378
rect	122	377	123	378
rect	124	377	125	378
rect	125	377	126	378
rect	126	377	127	378
rect	127	377	128	378
rect	128	377	129	378
rect	129	377	130	378
rect	131	377	132	378
rect	132	377	133	378
rect	134	377	135	378
rect	135	377	136	378
rect	136	377	137	378
rect	137	377	138	378
rect	143	377	144	378
rect	144	377	145	378
rect	146	377	147	378
rect	147	377	148	378
rect	149	377	150	378
rect	150	377	151	378
rect	152	377	153	378
rect	153	377	154	378
rect	154	377	155	378
rect	155	377	156	378
rect	156	377	157	378
rect	158	377	159	378
rect	159	377	160	378
rect	160	377	161	378
rect	161	377	162	378
rect	162	377	163	378
rect	163	377	164	378
rect	165	377	166	378
rect	166	377	167	378
rect	168	377	169	378
rect	169	377	170	378
rect	170	377	171	378
rect	171	377	172	378
rect	172	377	173	378
rect	173	377	174	378
rect	175	377	176	378
rect	176	377	177	378
rect	187	377	188	378
rect	188	377	189	378
rect	190	377	191	378
rect	191	377	192	378
rect	193	377	194	378
rect	194	377	195	378
rect	195	377	196	378
rect	196	377	197	378
rect	197	377	198	378
rect	198	377	199	378
rect	199	377	200	378
rect	200	377	201	378
rect	202	377	203	378
rect	203	377	204	378
rect	205	377	206	378
rect	206	377	207	378
rect	207	377	208	378
rect	208	377	209	378
rect	209	377	210	378
rect	210	377	211	378
rect	211	377	212	378
rect	212	377	213	378
rect	213	377	214	378
rect	214	377	215	378
rect	215	377	216	378
rect	216	377	217	378
rect	218	377	219	378
rect	219	377	220	378
rect	221	377	222	378
rect	222	377	223	378
rect	224	377	225	378
rect	225	377	226	378
rect	227	377	228	378
rect	228	377	229	378
rect	229	377	230	378
rect	230	377	231	378
rect	231	377	232	378
rect	233	377	234	378
rect	234	377	235	378
rect	236	377	237	378
rect	237	377	238	378
rect	238	377	239	378
rect	239	377	240	378
rect	240	377	241	378
rect	242	377	243	378
rect	243	377	244	378
rect	245	377	246	378
rect	246	377	247	378
rect	247	377	248	378
rect	248	377	249	378
rect	249	377	250	378
rect	250	377	251	378
rect	251	377	252	378
rect	252	377	253	378
rect	254	377	255	378
rect	255	377	256	378
rect	256	377	257	378
rect	257	377	258	378
rect	258	377	259	378
rect	266	377	267	378
rect	267	377	268	378
rect	269	377	270	378
rect	270	377	271	378
rect	272	377	273	378
rect	273	377	274	378
rect	275	377	276	378
rect	276	377	277	378
rect	278	377	279	378
rect	279	377	280	378
rect	281	377	282	378
rect	282	377	283	378
rect	284	377	285	378
rect	285	377	286	378
rect	286	377	287	378
rect	287	377	288	378
rect	288	377	289	378
rect	290	377	291	378
rect	291	377	292	378
rect	292	377	293	378
rect	293	377	294	378
rect	294	377	295	378
rect	296	377	297	378
rect	297	377	298	378
rect	298	377	299	378
rect	299	377	300	378
rect	300	377	301	378
rect	301	377	302	378
rect	302	377	303	378
rect	303	377	304	378
rect	304	377	305	378
rect	312	377	313	378
rect	313	377	314	378
rect	314	377	315	378
rect	315	377	316	378
rect	316	377	317	378
rect	321	377	322	378
rect	322	377	323	378
rect	324	377	325	378
rect	325	377	326	378
rect	327	377	328	378
rect	328	377	329	378
rect	329	377	330	378
rect	330	377	331	378
rect	331	377	332	378
rect	333	377	334	378
rect	334	377	335	378
rect	335	377	336	378
rect	336	377	337	378
rect	337	377	338	378
rect	338	377	339	378
rect	339	377	340	378
rect	340	377	341	378
rect	341	377	342	378
rect	342	377	343	378
rect	343	377	344	378
rect	344	377	345	378
rect	345	377	346	378
rect	347	377	348	378
rect	349	377	350	378
rect	350	377	351	378
rect	352	377	353	378
rect	353	377	354	378
rect	354	377	355	378
rect	355	377	356	378
rect	356	377	357	378
rect	357	377	358	378
rect	358	377	359	378
rect	359	377	360	378
rect	360	377	361	378
rect	361	377	362	378
rect	362	377	363	378
rect	363	377	364	378
rect	365	377	366	378
rect	366	377	367	378
rect	367	377	368	378
rect	368	377	369	378
rect	369	377	370	378
rect	370	377	371	378
rect	11	379	12	380
rect	12	379	13	380
rect	13	379	14	380
rect	52	379	53	380
rect	53	379	54	380
rect	54	379	55	380
rect	55	379	56	380
rect	56	379	57	380
rect	57	379	58	380
rect	64	379	65	380
rect	65	379	66	380
rect	66	379	67	380
rect	68	379	69	380
rect	69	379	70	380
rect	71	379	72	380
rect	72	379	73	380
rect	74	379	75	380
rect	75	379	76	380
rect	77	379	78	380
rect	78	379	79	380
rect	80	379	81	380
rect	81	379	82	380
rect	88	379	89	380
rect	89	379	90	380
rect	90	379	91	380
rect	92	379	93	380
rect	93	379	94	380
rect	95	379	96	380
rect	96	379	97	380
rect	116	379	117	380
rect	117	379	118	380
rect	119	379	120	380
rect	120	379	121	380
rect	122	379	123	380
rect	140	379	141	380
rect	141	379	142	380
rect	143	379	144	380
rect	144	379	145	380
rect	146	379	147	380
rect	147	379	148	380
rect	149	379	150	380
rect	150	379	151	380
rect	152	379	153	380
rect	153	379	154	380
rect	154	379	155	380
rect	155	379	156	380
rect	156	379	157	380
rect	158	379	159	380
rect	159	379	160	380
rect	160	379	161	380
rect	161	379	162	380
rect	162	379	163	380
rect	163	379	164	380
rect	165	379	166	380
rect	166	379	167	380
rect	168	379	169	380
rect	169	379	170	380
rect	170	379	171	380
rect	171	379	172	380
rect	172	379	173	380
rect	173	379	174	380
rect	184	379	185	380
rect	185	379	186	380
rect	187	379	188	380
rect	188	379	189	380
rect	190	379	191	380
rect	191	379	192	380
rect	193	379	194	380
rect	194	379	195	380
rect	195	379	196	380
rect	196	379	197	380
rect	197	379	198	380
rect	198	379	199	380
rect	199	379	200	380
rect	200	379	201	380
rect	202	379	203	380
rect	203	379	204	380
rect	224	379	225	380
rect	225	379	226	380
rect	230	379	231	380
rect	231	379	232	380
rect	233	379	234	380
rect	234	379	235	380
rect	257	379	258	380
rect	258	379	259	380
rect	259	379	260	380
rect	260	379	261	380
rect	261	379	262	380
rect	262	379	263	380
rect	263	379	264	380
rect	264	379	265	380
rect	266	379	267	380
rect	267	379	268	380
rect	269	379	270	380
rect	270	379	271	380
rect	272	379	273	380
rect	273	379	274	380
rect	275	379	276	380
rect	276	379	277	380
rect	287	379	288	380
rect	288	379	289	380
rect	299	379	300	380
rect	300	379	301	380
rect	301	379	302	380
rect	302	379	303	380
rect	303	379	304	380
rect	304	379	305	380
rect	305	379	306	380
rect	306	379	307	380
rect	307	379	308	380
rect	308	379	309	380
rect	309	379	310	380
rect	310	379	311	380
rect	312	379	313	380
rect	313	379	314	380
rect	314	379	315	380
rect	315	379	316	380
rect	316	379	317	380
rect	318	379	319	380
rect	319	379	320	380
rect	321	379	322	380
rect	322	379	323	380
rect	324	379	325	380
rect	325	379	326	380
rect	327	379	328	380
rect	328	379	329	380
rect	329	379	330	380
rect	330	379	331	380
rect	331	379	332	380
rect	333	379	334	380
rect	334	379	335	380
rect	335	379	336	380
rect	336	379	337	380
rect	337	379	338	380
rect	338	379	339	380
rect	339	379	340	380
rect	340	379	341	380
rect	341	379	342	380
rect	342	379	343	380
rect	343	379	344	380
rect	344	379	345	380
rect	345	379	346	380
rect	362	379	363	380
rect	363	379	364	380
rect	365	379	366	380
rect	366	379	367	380
rect	367	379	368	380
rect	368	379	369	380
rect	369	379	370	380
rect	370	379	371	380
rect	371	379	372	380
rect	372	379	373	380
rect	373	379	374	380
rect	374	379	375	380
rect	375	379	376	380
rect	376	379	377	380
rect	377	379	378	380
rect	378	379	379	380
rect	379	379	380	380
rect	380	379	381	380
rect	381	379	382	380
rect	382	379	383	380
rect	383	379	384	380
rect	384	379	385	380
rect	385	379	386	380
rect	386	379	387	380
rect	387	379	388	380
rect	388	379	389	380
rect	389	379	390	380
rect	390	379	391	380
rect	391	379	392	380
rect	278	388	279	389
rect	279	388	280	389
rect	281	388	282	389
rect	282	388	283	389
rect	284	388	285	389
rect	285	388	286	389
rect	264	390	265	391
rect	266	390	267	391
rect	267	390	268	391
rect	269	390	270	391
rect	270	390	271	391
rect	272	390	273	391
rect	273	390	274	391
rect	274	390	275	391
rect	275	390	276	391
rect	276	390	277	391
rect	277	390	278	391
rect	278	390	279	391
rect	279	390	280	391
rect	281	390	282	391
rect	282	390	283	391
rect	288	390	289	391
rect	290	390	291	391
rect	291	390	292	391
rect	292	390	293	391
rect	293	390	294	391
rect	294	390	295	391
rect	296	390	297	391
rect	297	390	298	391
rect	298	390	299	391
rect	299	390	300	391
rect	300	390	301	391
rect	301	390	302	391
rect	302	390	303	391
rect	303	390	304	391
rect	304	390	305	391
rect	305	390	306	391
rect	306	390	307	391
rect	307	390	308	391
rect	308	390	309	391
rect	309	390	310	391
rect	310	390	311	391
rect	312	390	313	391
rect	313	390	314	391
rect	314	390	315	391
rect	315	390	316	391
rect	316	390	317	391
rect	317	390	318	391
rect	318	390	319	391
rect	319	390	320	391
rect	321	390	322	391
rect	322	390	323	391
rect	122	392	123	393
rect	123	392	124	393
rect	125	392	126	393
rect	126	392	127	393
rect	213	392	214	393
rect	214	392	215	393
rect	215	392	216	393
rect	216	392	217	393
rect	218	392	219	393
rect	219	392	220	393
rect	221	392	222	393
rect	222	392	223	393
rect	223	392	224	393
rect	224	392	225	393
rect	225	392	226	393
rect	226	392	227	393
rect	227	392	228	393
rect	228	392	229	393
rect	230	392	231	393
rect	231	392	232	393
rect	233	392	234	393
rect	234	392	235	393
rect	235	392	236	393
rect	236	392	237	393
rect	237	392	238	393
rect	238	392	239	393
rect	239	392	240	393
rect	240	392	241	393
rect	261	392	262	393
rect	262	392	263	393
rect	264	392	265	393
rect	266	392	267	393
rect	267	392	268	393
rect	269	392	270	393
rect	270	392	271	393
rect	272	392	273	393
rect	273	392	274	393
rect	274	392	275	393
rect	275	392	276	393
rect	276	392	277	393
rect	277	392	278	393
rect	278	392	279	393
rect	279	392	280	393
rect	281	392	282	393
rect	282	392	283	393
rect	283	392	284	393
rect	284	392	285	393
rect	285	392	286	393
rect	286	392	287	393
rect	288	392	289	393
rect	290	392	291	393
rect	291	392	292	393
rect	292	392	293	393
rect	293	392	294	393
rect	294	392	295	393
rect	296	392	297	393
rect	297	392	298	393
rect	298	392	299	393
rect	299	392	300	393
rect	300	392	301	393
rect	301	392	302	393
rect	302	392	303	393
rect	303	392	304	393
rect	304	392	305	393
rect	305	392	306	393
rect	306	392	307	393
rect	307	392	308	393
rect	308	392	309	393
rect	309	392	310	393
rect	310	392	311	393
rect	122	394	123	395
rect	123	394	124	395
rect	125	394	126	395
rect	126	394	127	395
rect	127	394	128	395
rect	128	394	129	395
rect	129	394	130	395
rect	131	394	132	395
rect	132	394	133	395
rect	133	394	134	395
rect	134	394	135	395
rect	135	394	136	395
rect	136	394	137	395
rect	137	394	138	395
rect	138	394	139	395
rect	243	394	244	395
rect	245	394	246	395
rect	246	394	247	395
rect	247	394	248	395
rect	248	394	249	395
rect	249	394	250	395
rect	250	394	251	395
rect	251	394	252	395
rect	252	394	253	395
rect	254	394	255	395
rect	255	394	256	395
rect	257	394	258	395
rect	258	394	259	395
rect	259	394	260	395
rect	261	394	262	395
rect	262	394	263	395
rect	264	394	265	395
rect	266	394	267	395
rect	267	394	268	395
rect	269	394	270	395
rect	270	394	271	395
rect	285	394	286	395
rect	286	394	287	395
rect	288	394	289	395
rect	290	394	291	395
rect	291	394	292	395
rect	292	394	293	395
rect	293	394	294	395
rect	294	394	295	395
rect	296	394	297	395
rect	297	394	298	395
rect	298	394	299	395
rect	299	394	300	395
rect	300	394	301	395
rect	301	394	302	395
rect	302	394	303	395
rect	303	394	304	395
rect	304	394	305	395
rect	305	394	306	395
rect	306	394	307	395
rect	307	394	308	395
rect	308	394	309	395
rect	309	394	310	395
rect	310	394	311	395
rect	311	394	312	395
rect	312	394	313	395
rect	313	394	314	395
rect	314	394	315	395
rect	315	394	316	395
rect	316	394	317	395
rect	317	394	318	395
rect	318	394	319	395
rect	319	394	320	395
rect	321	394	322	395
rect	322	394	323	395
rect	323	394	324	395
rect	324	394	325	395
rect	325	394	326	395
rect	326	394	327	395
rect	327	394	328	395
rect	328	394	329	395
rect	329	394	330	395
rect	330	394	331	395
rect	331	394	332	395
rect	113	396	114	397
rect	114	396	115	397
rect	116	396	117	397
rect	117	396	118	397
rect	119	396	120	397
rect	120	396	121	397
rect	122	396	123	397
rect	123	396	124	397
rect	125	396	126	397
rect	126	396	127	397
rect	127	396	128	397
rect	128	396	129	397
rect	129	396	130	397
rect	141	396	142	397
rect	143	396	144	397
rect	144	396	145	397
rect	146	396	147	397
rect	147	396	148	397
rect	149	396	150	397
rect	150	396	151	397
rect	152	396	153	397
rect	153	396	154	397
rect	154	396	155	397
rect	155	396	156	397
rect	156	396	157	397
rect	157	396	158	397
rect	158	396	159	397
rect	159	396	160	397
rect	160	396	161	397
rect	161	396	162	397
rect	162	396	163	397
rect	163	396	164	397
rect	164	396	165	397
rect	165	396	166	397
rect	166	396	167	397
rect	168	396	169	397
rect	169	396	170	397
rect	170	396	171	397
rect	171	396	172	397
rect	172	396	173	397
rect	174	396	175	397
rect	175	396	176	397
rect	176	396	177	397
rect	177	396	178	397
rect	178	396	179	397
rect	179	396	180	397
rect	181	396	182	397
rect	182	396	183	397
rect	184	396	185	397
rect	185	396	186	397
rect	186	396	187	397
rect	187	396	188	397
rect	188	396	189	397
rect	189	396	190	397
rect	190	396	191	397
rect	191	396	192	397
rect	193	396	194	397
rect	194	396	195	397
rect	195	396	196	397
rect	196	396	197	397
rect	197	396	198	397
rect	198	396	199	397
rect	199	396	200	397
rect	200	396	201	397
rect	202	396	203	397
rect	203	396	204	397
rect	204	396	205	397
rect	205	396	206	397
rect	206	396	207	397
rect	207	396	208	397
rect	208	396	209	397
rect	209	396	210	397
rect	210	396	211	397
rect	211	396	212	397
rect	213	396	214	397
rect	214	396	215	397
rect	228	396	229	397
rect	230	396	231	397
rect	231	396	232	397
rect	233	396	234	397
rect	234	396	235	397
rect	235	396	236	397
rect	236	396	237	397
rect	237	396	238	397
rect	238	396	239	397
rect	239	396	240	397
rect	240	396	241	397
rect	241	396	242	397
rect	243	396	244	397
rect	245	396	246	397
rect	246	396	247	397
rect	247	396	248	397
rect	248	396	249	397
rect	249	396	250	397
rect	250	396	251	397
rect	251	396	252	397
rect	252	396	253	397
rect	254	396	255	397
rect	255	396	256	397
rect	257	396	258	397
rect	258	396	259	397
rect	259	396	260	397
rect	261	396	262	397
rect	262	396	263	397
rect	264	396	265	397
rect	281	396	282	397
rect	282	396	283	397
rect	283	396	284	397
rect	285	396	286	397
rect	286	396	287	397
rect	288	396	289	397
rect	294	396	295	397
rect	296	396	297	397
rect	297	396	298	397
rect	298	396	299	397
rect	299	396	300	397
rect	300	396	301	397
rect	301	396	302	397
rect	302	396	303	397
rect	303	396	304	397
rect	304	396	305	397
rect	305	396	306	397
rect	306	396	307	397
rect	307	396	308	397
rect	308	396	309	397
rect	309	396	310	397
rect	310	396	311	397
rect	311	396	312	397
rect	312	396	313	397
rect	313	396	314	397
rect	314	396	315	397
rect	315	396	316	397
rect	316	396	317	397
rect	317	396	318	397
rect	318	396	319	397
rect	319	396	320	397
rect	321	396	322	397
rect	322	396	323	397
rect	323	396	324	397
rect	324	396	325	397
rect	325	396	326	397
rect	326	396	327	397
rect	327	396	328	397
rect	328	396	329	397
rect	329	396	330	397
rect	330	396	331	397
rect	331	396	332	397
rect	332	396	333	397
rect	333	396	334	397
rect	334	396	335	397
rect	335	396	336	397
rect	336	396	337	397
rect	337	396	338	397
rect	339	396	340	397
rect	340	396	341	397
rect	341	396	342	397
rect	342	396	343	397
rect	343	396	344	397
rect	344	396	345	397
rect	346	396	347	397
rect	347	396	348	397
rect	349	396	350	397
rect	350	396	351	397
rect	351	396	352	397
rect	352	396	353	397
rect	353	396	354	397
rect	131	398	132	399
rect	132	398	133	399
rect	133	398	134	399
rect	134	398	135	399
rect	135	398	136	399
rect	136	398	137	399
rect	137	398	138	399
rect	138	398	139	399
rect	139	398	140	399
rect	141	398	142	399
rect	143	398	144	399
rect	144	398	145	399
rect	146	398	147	399
rect	147	398	148	399
rect	202	398	203	399
rect	203	398	204	399
rect	204	398	205	399
rect	205	398	206	399
rect	210	398	211	399
rect	211	398	212	399
rect	213	398	214	399
rect	214	398	215	399
rect	216	398	217	399
rect	218	398	219	399
rect	219	398	220	399
rect	221	398	222	399
rect	222	398	223	399
rect	223	398	224	399
rect	224	398	225	399
rect	225	398	226	399
rect	226	398	227	399
rect	228	398	229	399
rect	240	398	241	399
rect	241	398	242	399
rect	243	398	244	399
rect	245	398	246	399
rect	246	398	247	399
rect	247	398	248	399
rect	248	398	249	399
rect	249	398	250	399
rect	250	398	251	399
rect	251	398	252	399
rect	252	398	253	399
rect	257	398	258	399
rect	258	398	259	399
rect	259	398	260	399
rect	261	398	262	399
rect	262	398	263	399
rect	264	398	265	399
rect	265	398	266	399
rect	276	398	277	399
rect	277	398	278	399
rect	278	398	279	399
rect	279	398	280	399
rect	280	398	281	399
rect	281	398	282	399
rect	282	398	283	399
rect	283	398	284	399
rect	285	398	286	399
rect	286	398	287	399
rect	288	398	289	399
rect	289	398	290	399
rect	290	398	291	399
rect	291	398	292	399
rect	292	398	293	399
rect	294	398	295	399
rect	296	398	297	399
rect	297	398	298	399
rect	298	398	299	399
rect	299	398	300	399
rect	300	398	301	399
rect	301	398	302	399
rect	302	398	303	399
rect	303	398	304	399
rect	304	398	305	399
rect	305	398	306	399
rect	306	398	307	399
rect	307	398	308	399
rect	308	398	309	399
rect	309	398	310	399
rect	310	398	311	399
rect	311	398	312	399
rect	312	398	313	399
rect	313	398	314	399
rect	314	398	315	399
rect	315	398	316	399
rect	316	398	317	399
rect	317	398	318	399
rect	318	398	319	399
rect	319	398	320	399
rect	332	398	333	399
rect	333	398	334	399
rect	334	398	335	399
rect	335	398	336	399
rect	336	398	337	399
rect	337	398	338	399
rect	339	398	340	399
rect	340	398	341	399
rect	341	398	342	399
rect	342	398	343	399
rect	343	398	344	399
rect	344	398	345	399
rect	346	398	347	399
rect	347	398	348	399
rect	349	398	350	399
rect	350	398	351	399
rect	351	398	352	399
rect	352	398	353	399
rect	353	398	354	399
rect	354	398	355	399
rect	355	398	356	399
rect	356	398	357	399
rect	357	398	358	399
rect	358	398	359	399
rect	359	398	360	399
rect	360	398	361	399
rect	361	398	362	399
rect	362	398	363	399
rect	363	398	364	399
rect	64	400	65	401
rect	65	400	66	401
rect	66	400	67	401
rect	68	400	69	401
rect	69	400	70	401
rect	98	400	99	401
rect	99	400	100	401
rect	100	400	101	401
rect	101	400	102	401
rect	102	400	103	401
rect	103	400	104	401
rect	104	400	105	401
rect	105	400	106	401
rect	107	400	108	401
rect	108	400	109	401
rect	109	400	110	401
rect	110	400	111	401
rect	111	400	112	401
rect	113	400	114	401
rect	114	400	115	401
rect	116	400	117	401
rect	117	400	118	401
rect	119	400	120	401
rect	120	400	121	401
rect	122	400	123	401
rect	123	400	124	401
rect	125	400	126	401
rect	126	400	127	401
rect	127	400	128	401
rect	128	400	129	401
rect	129	400	130	401
rect	131	400	132	401
rect	132	400	133	401
rect	133	400	134	401
rect	134	400	135	401
rect	135	400	136	401
rect	136	400	137	401
rect	137	400	138	401
rect	138	400	139	401
rect	139	400	140	401
rect	141	400	142	401
rect	143	400	144	401
rect	144	400	145	401
rect	146	400	147	401
rect	147	400	148	401
rect	148	400	149	401
rect	149	400	150	401
rect	150	400	151	401
rect	152	400	153	401
rect	153	400	154	401
rect	154	400	155	401
rect	155	400	156	401
rect	156	400	157	401
rect	157	400	158	401
rect	158	400	159	401
rect	159	400	160	401
rect	160	400	161	401
rect	161	400	162	401
rect	162	400	163	401
rect	163	400	164	401
rect	164	400	165	401
rect	165	400	166	401
rect	166	400	167	401
rect	168	400	169	401
rect	169	400	170	401
rect	170	400	171	401
rect	171	400	172	401
rect	172	400	173	401
rect	174	400	175	401
rect	175	400	176	401
rect	176	400	177	401
rect	177	400	178	401
rect	178	400	179	401
rect	179	400	180	401
rect	181	400	182	401
rect	182	400	183	401
rect	184	400	185	401
rect	185	400	186	401
rect	186	400	187	401
rect	187	400	188	401
rect	188	400	189	401
rect	189	400	190	401
rect	190	400	191	401
rect	191	400	192	401
rect	193	400	194	401
rect	194	400	195	401
rect	195	400	196	401
rect	196	400	197	401
rect	197	400	198	401
rect	198	400	199	401
rect	199	400	200	401
rect	200	400	201	401
rect	201	400	202	401
rect	202	400	203	401
rect	203	400	204	401
rect	204	400	205	401
rect	205	400	206	401
rect	207	400	208	401
rect	208	400	209	401
rect	210	400	211	401
rect	211	400	212	401
rect	213	400	214	401
rect	214	400	215	401
rect	216	400	217	401
rect	218	400	219	401
rect	219	400	220	401
rect	221	400	222	401
rect	222	400	223	401
rect	223	400	224	401
rect	224	400	225	401
rect	225	400	226	401
rect	226	400	227	401
rect	228	400	229	401
rect	229	400	230	401
rect	230	400	231	401
rect	231	400	232	401
rect	233	400	234	401
rect	234	400	235	401
rect	235	400	236	401
rect	236	400	237	401
rect	237	400	238	401
rect	238	400	239	401
rect	240	400	241	401
rect	241	400	242	401
rect	243	400	244	401
rect	245	400	246	401
rect	246	400	247	401
rect	247	400	248	401
rect	248	400	249	401
rect	249	400	250	401
rect	250	400	251	401
rect	251	400	252	401
rect	252	400	253	401
rect	253	400	254	401
rect	254	400	255	401
rect	255	400	256	401
rect	256	400	257	401
rect	257	400	258	401
rect	258	400	259	401
rect	259	400	260	401
rect	261	400	262	401
rect	262	400	263	401
rect	264	400	265	401
rect	265	400	266	401
rect	267	400	268	401
rect	269	400	270	401
rect	270	400	271	401
rect	271	400	272	401
rect	272	400	273	401
rect	273	400	274	401
rect	274	400	275	401
rect	276	400	277	401
rect	277	400	278	401
rect	278	400	279	401
rect	279	400	280	401
rect	280	400	281	401
rect	281	400	282	401
rect	282	400	283	401
rect	283	400	284	401
rect	285	400	286	401
rect	286	400	287	401
rect	288	400	289	401
rect	289	400	290	401
rect	290	400	291	401
rect	291	400	292	401
rect	292	400	293	401
rect	294	400	295	401
rect	296	400	297	401
rect	297	400	298	401
rect	298	400	299	401
rect	299	400	300	401
rect	300	400	301	401
rect	301	400	302	401
rect	302	400	303	401
rect	303	400	304	401
rect	304	400	305	401
rect	305	400	306	401
rect	313	400	314	401
rect	314	400	315	401
rect	315	400	316	401
rect	316	400	317	401
rect	317	400	318	401
rect	329	400	330	401
rect	330	400	331	401
rect	332	400	333	401
rect	333	400	334	401
rect	334	400	335	401
rect	335	400	336	401
rect	336	400	337	401
rect	337	400	338	401
rect	339	400	340	401
rect	340	400	341	401
rect	341	400	342	401
rect	342	400	343	401
rect	343	400	344	401
rect	344	400	345	401
rect	346	400	347	401
rect	347	400	348	401
rect	61	402	62	403
rect	62	402	63	403
rect	64	402	65	403
rect	65	402	66	403
rect	66	402	67	403
rect	77	402	78	403
rect	78	402	79	403
rect	80	402	81	403
rect	82	402	83	403
rect	83	402	84	403
rect	98	402	99	403
rect	99	402	100	403
rect	100	402	101	403
rect	101	402	102	403
rect	102	402	103	403
rect	103	402	104	403
rect	104	402	105	403
rect	105	402	106	403
rect	119	402	120	403
rect	120	402	121	403
rect	122	402	123	403
rect	123	402	124	403
rect	128	402	129	403
rect	129	402	130	403
rect	131	402	132	403
rect	132	402	133	403
rect	133	402	134	403
rect	134	402	135	403
rect	135	402	136	403
rect	136	402	137	403
rect	137	402	138	403
rect	138	402	139	403
rect	139	402	140	403
rect	141	402	142	403
rect	143	402	144	403
rect	144	402	145	403
rect	198	402	199	403
rect	199	402	200	403
rect	200	402	201	403
rect	201	402	202	403
rect	202	402	203	403
rect	203	402	204	403
rect	204	402	205	403
rect	205	402	206	403
rect	207	402	208	403
rect	208	402	209	403
rect	210	402	211	403
rect	211	402	212	403
rect	213	402	214	403
rect	214	402	215	403
rect	216	402	217	403
rect	231	402	232	403
rect	237	402	238	403
rect	238	402	239	403
rect	240	402	241	403
rect	241	402	242	403
rect	243	402	244	403
rect	245	402	246	403
rect	246	402	247	403
rect	247	402	248	403
rect	248	402	249	403
rect	249	402	250	403
rect	250	402	251	403
rect	251	402	252	403
rect	252	402	253	403
rect	253	402	254	403
rect	254	402	255	403
rect	255	402	256	403
rect	256	402	257	403
rect	257	402	258	403
rect	258	402	259	403
rect	259	402	260	403
rect	261	402	262	403
rect	262	402	263	403
rect	264	402	265	403
rect	265	402	266	403
rect	267	402	268	403
rect	273	402	274	403
rect	274	402	275	403
rect	276	402	277	403
rect	277	402	278	403
rect	278	402	279	403
rect	279	402	280	403
rect	280	402	281	403
rect	281	402	282	403
rect	282	402	283	403
rect	283	402	284	403
rect	285	402	286	403
rect	286	402	287	403
rect	288	402	289	403
rect	289	402	290	403
rect	290	402	291	403
rect	291	402	292	403
rect	292	402	293	403
rect	294	402	295	403
rect	296	402	297	403
rect	297	402	298	403
rect	298	402	299	403
rect	299	402	300	403
rect	300	402	301	403
rect	301	402	302	403
rect	302	402	303	403
rect	303	402	304	403
rect	304	402	305	403
rect	305	402	306	403
rect	307	402	308	403
rect	308	402	309	403
rect	309	402	310	403
rect	310	402	311	403
rect	311	402	312	403
rect	313	402	314	403
rect	314	402	315	403
rect	315	402	316	403
rect	316	402	317	403
rect	317	402	318	403
rect	319	402	320	403
rect	320	402	321	403
rect	321	402	322	403
rect	322	402	323	403
rect	323	402	324	403
rect	324	402	325	403
rect	325	402	326	403
rect	326	402	327	403
rect	327	402	328	403
rect	329	402	330	403
rect	330	402	331	403
rect	332	402	333	403
rect	333	402	334	403
rect	334	402	335	403
rect	335	402	336	403
rect	336	402	337	403
rect	337	402	338	403
rect	5	404	6	405
rect	6	404	7	405
rect	7	404	8	405
rect	15	404	16	405
rect	16	404	17	405
rect	17	404	18	405
rect	18	404	19	405
rect	19	404	20	405
rect	59	404	60	405
rect	61	404	62	405
rect	62	404	63	405
rect	64	404	65	405
rect	65	404	66	405
rect	74	404	75	405
rect	95	404	96	405
rect	96	404	97	405
rect	98	404	99	405
rect	99	404	100	405
rect	110	404	111	405
rect	111	404	112	405
rect	113	404	114	405
rect	114	404	115	405
rect	125	404	126	405
rect	126	404	127	405
rect	128	404	129	405
rect	129	404	130	405
rect	131	404	132	405
rect	132	404	133	405
rect	133	404	134	405
rect	134	404	135	405
rect	135	404	136	405
rect	136	404	137	405
rect	137	404	138	405
rect	138	404	139	405
rect	139	404	140	405
rect	141	404	142	405
rect	147	404	148	405
rect	148	404	149	405
rect	149	404	150	405
rect	150	404	151	405
rect	168	404	169	405
rect	169	404	170	405
rect	170	404	171	405
rect	171	404	172	405
rect	172	404	173	405
rect	181	404	182	405
rect	182	404	183	405
rect	193	404	194	405
rect	194	404	195	405
rect	195	404	196	405
rect	196	404	197	405
rect	198	404	199	405
rect	199	404	200	405
rect	219	404	220	405
rect	220	404	221	405
rect	222	404	223	405
rect	223	404	224	405
rect	224	404	225	405
rect	225	404	226	405
rect	226	404	227	405
rect	228	404	229	405
rect	229	404	230	405
rect	231	404	232	405
rect	232	404	233	405
rect	233	404	234	405
rect	234	404	235	405
rect	235	404	236	405
rect	237	404	238	405
rect	238	404	239	405
rect	240	404	241	405
rect	241	404	242	405
rect	243	404	244	405
rect	252	404	253	405
rect	253	404	254	405
rect	254	404	255	405
rect	255	404	256	405
rect	256	404	257	405
rect	257	404	258	405
rect	258	404	259	405
rect	259	404	260	405
rect	261	404	262	405
rect	262	404	263	405
rect	264	404	265	405
rect	265	404	266	405
rect	267	404	268	405
rect	268	404	269	405
rect	269	404	270	405
rect	270	404	271	405
rect	271	404	272	405
rect	273	404	274	405
rect	274	404	275	405
rect	276	404	277	405
rect	277	404	278	405
rect	278	404	279	405
rect	279	404	280	405
rect	280	404	281	405
rect	281	404	282	405
rect	282	404	283	405
rect	283	404	284	405
rect	285	404	286	405
rect	286	404	287	405
rect	288	404	289	405
rect	289	404	290	405
rect	290	404	291	405
rect	291	404	292	405
rect	292	404	293	405
rect	294	404	295	405
rect	304	404	305	405
rect	305	404	306	405
rect	307	404	308	405
rect	308	404	309	405
rect	309	404	310	405
rect	310	404	311	405
rect	311	404	312	405
rect	313	404	314	405
rect	314	404	315	405
rect	315	404	316	405
rect	316	404	317	405
rect	317	404	318	405
rect	319	404	320	405
rect	320	404	321	405
rect	321	404	322	405
rect	322	404	323	405
rect	323	404	324	405
rect	324	404	325	405
rect	325	404	326	405
rect	326	404	327	405
rect	327	404	328	405
rect	329	404	330	405
rect	330	404	331	405
rect	332	404	333	405
rect	333	404	334	405
rect	334	404	335	405
rect	335	404	336	405
rect	336	404	337	405
rect	337	404	338	405
rect	338	404	339	405
rect	339	404	340	405
rect	340	404	341	405
rect	341	404	342	405
rect	342	404	343	405
rect	343	404	344	405
rect	344	404	345	405
rect	73	413	74	414
rect	74	413	75	414
rect	76	413	77	414
rect	77	413	78	414
rect	90	413	91	414
rect	91	413	92	414
rect	92	413	93	414
rect	93	413	94	414
rect	94	413	95	414
rect	95	413	96	414
rect	96	413	97	414
rect	98	413	99	414
rect	99	413	100	414
rect	101	413	102	414
rect	102	413	103	414
rect	104	413	105	414
rect	105	413	106	414
rect	106	413	107	414
rect	107	413	108	414
rect	108	413	109	414
rect	110	413	111	414
rect	111	413	112	414
rect	238	413	239	414
rect	240	413	241	414
rect	241	413	242	414
rect	243	413	244	414
rect	244	413	245	414
rect	245	413	246	414
rect	246	413	247	414
rect	247	413	248	414
rect	248	413	249	414
rect	249	413	250	414
rect	250	413	251	414
rect	252	413	253	414
rect	253	413	254	414
rect	254	413	255	414
rect	255	413	256	414
rect	256	413	257	414
rect	258	413	259	414
rect	259	413	260	414
rect	261	413	262	414
rect	262	413	263	414
rect	269	413	270	414
rect	270	413	271	414
rect	271	413	272	414
rect	272	413	273	414
rect	273	413	274	414
rect	274	413	275	414
rect	276	413	277	414
rect	277	413	278	414
rect	279	413	280	414
rect	280	413	281	414
rect	281	413	282	414
rect	282	413	283	414
rect	283	413	284	414
rect	285	413	286	414
rect	286	413	287	414
rect	288	413	289	414
rect	289	413	290	414
rect	290	413	291	414
rect	291	413	292	414
rect	292	413	293	414
rect	294	413	295	414
rect	295	413	296	414
rect	296	413	297	414
rect	298	413	299	414
rect	299	413	300	414
rect	300	413	301	414
rect	301	413	302	414
rect	302	413	303	414
rect	304	413	305	414
rect	305	413	306	414
rect	307	413	308	414
rect	308	413	309	414
rect	309	413	310	414
rect	310	413	311	414
rect	311	413	312	414
rect	76	415	77	416
rect	110	415	111	416
rect	111	415	112	416
rect	112	415	113	416
rect	119	415	120	416
rect	120	415	121	416
rect	144	415	145	416
rect	145	415	146	416
rect	147	415	148	416
rect	148	415	149	416
rect	149	415	150	416
rect	150	415	151	416
rect	151	415	152	416
rect	152	415	153	416
rect	153	415	154	416
rect	154	415	155	416
rect	155	415	156	416
rect	156	415	157	416
rect	157	415	158	416
rect	158	415	159	416
rect	159	415	160	416
rect	160	415	161	416
rect	161	415	162	416
rect	162	415	163	416
rect	163	415	164	416
rect	164	415	165	416
rect	165	415	166	416
rect	166	415	167	416
rect	167	415	168	416
rect	168	415	169	416
rect	169	415	170	416
rect	170	415	171	416
rect	171	415	172	416
rect	172	415	173	416
rect	173	415	174	416
rect	174	415	175	416
rect	175	415	176	416
rect	176	415	177	416
rect	177	415	178	416
rect	178	415	179	416
rect	179	415	180	416
rect	180	415	181	416
rect	181	415	182	416
rect	182	415	183	416
rect	183	415	184	416
rect	184	415	185	416
rect	185	415	186	416
rect	186	415	187	416
rect	187	415	188	416
rect	188	415	189	416
rect	189	415	190	416
rect	190	415	191	416
rect	191	415	192	416
rect	192	415	193	416
rect	193	415	194	416
rect	194	415	195	416
rect	195	415	196	416
rect	196	415	197	416
rect	198	415	199	416
rect	199	415	200	416
rect	201	415	202	416
rect	202	415	203	416
rect	203	415	204	416
rect	204	415	205	416
rect	205	415	206	416
rect	207	415	208	416
rect	208	415	209	416
rect	210	415	211	416
rect	211	415	212	416
rect	213	415	214	416
rect	214	415	215	416
rect	215	415	216	416
rect	216	415	217	416
rect	217	415	218	416
rect	219	415	220	416
rect	220	415	221	416
rect	222	415	223	416
rect	223	415	224	416
rect	224	415	225	416
rect	225	415	226	416
rect	226	415	227	416
rect	227	415	228	416
rect	228	415	229	416
rect	229	415	230	416
rect	263	415	264	416
rect	264	415	265	416
rect	265	415	266	416
rect	267	415	268	416
rect	269	415	270	416
rect	270	415	271	416
rect	271	415	272	416
rect	272	415	273	416
rect	273	415	274	416
rect	274	415	275	416
rect	276	415	277	416
rect	277	415	278	416
rect	279	415	280	416
rect	280	415	281	416
rect	281	415	282	416
rect	282	415	283	416
rect	283	415	284	416
rect	285	415	286	416
rect	286	415	287	416
rect	288	415	289	416
rect	289	415	290	416
rect	290	415	291	416
rect	291	415	292	416
rect	292	415	293	416
rect	294	415	295	416
rect	295	415	296	416
rect	296	415	297	416
rect	75	417	76	418
rect	76	417	77	418
rect	78	417	79	418
rect	79	417	80	418
rect	80	417	81	418
rect	82	417	83	418
rect	83	417	84	418
rect	84	417	85	418
rect	85	417	86	418
rect	86	417	87	418
rect	87	417	88	418
rect	88	417	89	418
rect	90	417	91	418
rect	91	417	92	418
rect	92	417	93	418
rect	93	417	94	418
rect	94	417	95	418
rect	95	417	96	418
rect	96	417	97	418
rect	98	417	99	418
rect	99	417	100	418
rect	101	417	102	418
rect	102	417	103	418
rect	104	417	105	418
rect	105	417	106	418
rect	106	417	107	418
rect	107	417	108	418
rect	108	417	109	418
rect	109	417	110	418
rect	110	417	111	418
rect	111	417	112	418
rect	112	417	113	418
rect	114	417	115	418
rect	115	417	116	418
rect	116	417	117	418
rect	117	417	118	418
rect	118	417	119	418
rect	119	417	120	418
rect	120	417	121	418
rect	121	417	122	418
rect	122	417	123	418
rect	123	417	124	418
rect	125	417	126	418
rect	126	417	127	418
rect	128	417	129	418
rect	129	417	130	418
rect	131	417	132	418
rect	132	417	133	418
rect	134	417	135	418
rect	135	417	136	418
rect	136	417	137	418
rect	137	417	138	418
rect	138	417	139	418
rect	139	417	140	418
rect	140	417	141	418
rect	141	417	142	418
rect	142	417	143	418
rect	143	417	144	418
rect	144	417	145	418
rect	145	417	146	418
rect	147	417	148	418
rect	148	417	149	418
rect	149	417	150	418
rect	150	417	151	418
rect	151	417	152	418
rect	152	417	153	418
rect	153	417	154	418
rect	154	417	155	418
rect	155	417	156	418
rect	156	417	157	418
rect	157	417	158	418
rect	158	417	159	418
rect	159	417	160	418
rect	160	417	161	418
rect	161	417	162	418
rect	162	417	163	418
rect	163	417	164	418
rect	164	417	165	418
rect	165	417	166	418
rect	166	417	167	418
rect	167	417	168	418
rect	168	417	169	418
rect	169	417	170	418
rect	170	417	171	418
rect	171	417	172	418
rect	172	417	173	418
rect	173	417	174	418
rect	174	417	175	418
rect	175	417	176	418
rect	176	417	177	418
rect	177	417	178	418
rect	178	417	179	418
rect	179	417	180	418
rect	180	417	181	418
rect	181	417	182	418
rect	182	417	183	418
rect	183	417	184	418
rect	184	417	185	418
rect	185	417	186	418
rect	186	417	187	418
rect	187	417	188	418
rect	188	417	189	418
rect	189	417	190	418
rect	190	417	191	418
rect	191	417	192	418
rect	192	417	193	418
rect	193	417	194	418
rect	194	417	195	418
rect	195	417	196	418
rect	196	417	197	418
rect	198	417	199	418
rect	199	417	200	418
rect	201	417	202	418
rect	202	417	203	418
rect	203	417	204	418
rect	204	417	205	418
rect	205	417	206	418
rect	207	417	208	418
rect	208	417	209	418
rect	210	417	211	418
rect	211	417	212	418
rect	213	417	214	418
rect	214	417	215	418
rect	215	417	216	418
rect	216	417	217	418
rect	217	417	218	418
rect	219	417	220	418
rect	220	417	221	418
rect	232	417	233	418
rect	233	417	234	418
rect	234	417	235	418
rect	235	417	236	418
rect	236	417	237	418
rect	238	417	239	418
rect	254	417	255	418
rect	255	417	256	418
rect	256	417	257	418
rect	258	417	259	418
rect	259	417	260	418
rect	261	417	262	418
rect	263	417	264	418
rect	264	417	265	418
rect	265	417	266	418
rect	267	417	268	418
rect	269	417	270	418
rect	270	417	271	418
rect	271	417	272	418
rect	272	417	273	418
rect	273	417	274	418
rect	274	417	275	418
rect	276	417	277	418
rect	277	417	278	418
rect	279	417	280	418
rect	280	417	281	418
rect	281	417	282	418
rect	282	417	283	418
rect	283	417	284	418
rect	285	417	286	418
rect	286	417	287	418
rect	288	417	289	418
rect	289	417	290	418
rect	290	417	291	418
rect	291	417	292	418
rect	292	417	293	418
rect	294	417	295	418
rect	295	417	296	418
rect	296	417	297	418
rect	297	417	298	418
rect	298	417	299	418
rect	299	417	300	418
rect	300	417	301	418
rect	301	417	302	418
rect	302	417	303	418
rect	304	417	305	418
rect	305	417	306	418
rect	67	419	68	420
rect	68	419	69	420
rect	69	419	70	420
rect	70	419	71	420
rect	71	419	72	420
rect	72	419	73	420
rect	73	419	74	420
rect	75	419	76	420
rect	76	419	77	420
rect	78	419	79	420
rect	79	419	80	420
rect	80	419	81	420
rect	82	419	83	420
rect	83	419	84	420
rect	84	419	85	420
rect	85	419	86	420
rect	86	419	87	420
rect	87	419	88	420
rect	88	419	89	420
rect	90	419	91	420
rect	91	419	92	420
rect	92	419	93	420
rect	93	419	94	420
rect	94	419	95	420
rect	95	419	96	420
rect	96	419	97	420
rect	98	419	99	420
rect	99	419	100	420
rect	101	419	102	420
rect	102	419	103	420
rect	104	419	105	420
rect	105	419	106	420
rect	106	419	107	420
rect	107	419	108	420
rect	108	419	109	420
rect	109	419	110	420
rect	110	419	111	420
rect	111	419	112	420
rect	112	419	113	420
rect	114	419	115	420
rect	115	419	116	420
rect	116	419	117	420
rect	117	419	118	420
rect	118	419	119	420
rect	119	419	120	420
rect	120	419	121	420
rect	121	419	122	420
rect	122	419	123	420
rect	123	419	124	420
rect	125	419	126	420
rect	126	419	127	420
rect	128	419	129	420
rect	129	419	130	420
rect	131	419	132	420
rect	132	419	133	420
rect	134	419	135	420
rect	135	419	136	420
rect	136	419	137	420
rect	137	419	138	420
rect	138	419	139	420
rect	139	419	140	420
rect	140	419	141	420
rect	141	419	142	420
rect	142	419	143	420
rect	143	419	144	420
rect	144	419	145	420
rect	145	419	146	420
rect	147	419	148	420
rect	148	419	149	420
rect	149	419	150	420
rect	150	419	151	420
rect	151	419	152	420
rect	152	419	153	420
rect	153	419	154	420
rect	154	419	155	420
rect	155	419	156	420
rect	156	419	157	420
rect	157	419	158	420
rect	158	419	159	420
rect	159	419	160	420
rect	160	419	161	420
rect	161	419	162	420
rect	162	419	163	420
rect	163	419	164	420
rect	164	419	165	420
rect	165	419	166	420
rect	166	419	167	420
rect	167	419	168	420
rect	168	419	169	420
rect	169	419	170	420
rect	170	419	171	420
rect	171	419	172	420
rect	172	419	173	420
rect	173	419	174	420
rect	174	419	175	420
rect	175	419	176	420
rect	176	419	177	420
rect	177	419	178	420
rect	178	419	179	420
rect	179	419	180	420
rect	180	419	181	420
rect	181	419	182	420
rect	182	419	183	420
rect	183	419	184	420
rect	184	419	185	420
rect	185	419	186	420
rect	186	419	187	420
rect	187	419	188	420
rect	188	419	189	420
rect	189	419	190	420
rect	190	419	191	420
rect	191	419	192	420
rect	192	419	193	420
rect	193	419	194	420
rect	194	419	195	420
rect	195	419	196	420
rect	196	419	197	420
rect	198	419	199	420
rect	199	419	200	420
rect	201	419	202	420
rect	202	419	203	420
rect	203	419	204	420
rect	204	419	205	420
rect	205	419	206	420
rect	225	419	226	420
rect	226	419	227	420
rect	227	419	228	420
rect	228	419	229	420
rect	229	419	230	420
rect	230	419	231	420
rect	232	419	233	420
rect	233	419	234	420
rect	234	419	235	420
rect	235	419	236	420
rect	236	419	237	420
rect	238	419	239	420
rect	239	419	240	420
rect	240	419	241	420
rect	241	419	242	420
rect	243	419	244	420
rect	244	419	245	420
rect	245	419	246	420
rect	246	419	247	420
rect	247	419	248	420
rect	248	419	249	420
rect	249	419	250	420
rect	250	419	251	420
rect	252	419	253	420
rect	254	419	255	420
rect	255	419	256	420
rect	256	419	257	420
rect	258	419	259	420
rect	259	419	260	420
rect	261	419	262	420
rect	263	419	264	420
rect	264	419	265	420
rect	265	419	266	420
rect	267	419	268	420
rect	269	419	270	420
rect	270	419	271	420
rect	271	419	272	420
rect	272	419	273	420
rect	273	419	274	420
rect	274	419	275	420
rect	282	419	283	420
rect	283	419	284	420
rect	285	419	286	420
rect	286	419	287	420
rect	288	419	289	420
rect	289	419	290	420
rect	290	419	291	420
rect	291	419	292	420
rect	292	419	293	420
rect	294	419	295	420
rect	295	419	296	420
rect	296	419	297	420
rect	297	419	298	420
rect	298	419	299	420
rect	299	419	300	420
rect	300	419	301	420
rect	301	419	302	420
rect	302	419	303	420
rect	108	421	109	422
rect	109	421	110	422
rect	110	421	111	422
rect	111	421	112	422
rect	112	421	113	422
rect	114	421	115	422
rect	115	421	116	422
rect	116	421	117	422
rect	117	421	118	422
rect	118	421	119	422
rect	119	421	120	422
rect	120	421	121	422
rect	121	421	122	422
rect	122	421	123	422
rect	123	421	124	422
rect	125	421	126	422
rect	126	421	127	422
rect	128	421	129	422
rect	129	421	130	422
rect	187	421	188	422
rect	188	421	189	422
rect	189	421	190	422
rect	190	421	191	422
rect	191	421	192	422
rect	192	421	193	422
rect	193	421	194	422
rect	194	421	195	422
rect	195	421	196	422
rect	196	421	197	422
rect	206	421	207	422
rect	207	421	208	422
rect	208	421	209	422
rect	210	421	211	422
rect	211	421	212	422
rect	213	421	214	422
rect	214	421	215	422
rect	215	421	216	422
rect	216	421	217	422
rect	217	421	218	422
rect	222	421	223	422
rect	223	421	224	422
rect	225	421	226	422
rect	226	421	227	422
rect	227	421	228	422
rect	228	421	229	422
rect	229	421	230	422
rect	230	421	231	422
rect	232	421	233	422
rect	233	421	234	422
rect	234	421	235	422
rect	235	421	236	422
rect	236	421	237	422
rect	238	421	239	422
rect	239	421	240	422
rect	240	421	241	422
rect	241	421	242	422
rect	248	421	249	422
rect	249	421	250	422
rect	250	421	251	422
rect	252	421	253	422
rect	254	421	255	422
rect	255	421	256	422
rect	256	421	257	422
rect	258	421	259	422
rect	259	421	260	422
rect	261	421	262	422
rect	263	421	264	422
rect	264	421	265	422
rect	265	421	266	422
rect	267	421	268	422
rect	269	421	270	422
rect	270	421	271	422
rect	271	421	272	422
rect	272	421	273	422
rect	273	421	274	422
rect	274	421	275	422
rect	275	421	276	422
rect	276	421	277	422
rect	277	421	278	422
rect	279	421	280	422
rect	280	421	281	422
rect	282	421	283	422
rect	283	421	284	422
rect	285	421	286	422
rect	286	421	287	422
rect	288	421	289	422
rect	289	421	290	422
rect	290	421	291	422
rect	291	421	292	422
rect	292	421	293	422
rect	294	421	295	422
rect	295	421	296	422
rect	296	421	297	422
rect	297	421	298	422
rect	298	421	299	422
rect	299	421	300	422
rect	300	421	301	422
rect	301	421	302	422
rect	302	421	303	422
rect	303	421	304	422
rect	304	421	305	422
rect	305	421	306	422
rect	306	421	307	422
rect	307	421	308	422
rect	308	421	309	422
rect	309	421	310	422
rect	310	421	311	422
rect	311	421	312	422
rect	312	421	313	422
rect	313	421	314	422
rect	314	421	315	422
rect	315	421	316	422
rect	316	421	317	422
rect	317	421	318	422
rect	318	421	319	422
rect	319	421	320	422
rect	320	421	321	422
rect	321	421	322	422
rect	322	421	323	422
rect	323	421	324	422
rect	324	421	325	422
rect	104	423	105	424
rect	105	423	106	424
rect	106	423	107	424
rect	108	423	109	424
rect	109	423	110	424
rect	110	423	111	424
rect	111	423	112	424
rect	112	423	113	424
rect	114	423	115	424
rect	115	423	116	424
rect	116	423	117	424
rect	117	423	118	424
rect	118	423	119	424
rect	119	423	120	424
rect	120	423	121	424
rect	121	423	122	424
rect	122	423	123	424
rect	123	423	124	424
rect	125	423	126	424
rect	126	423	127	424
rect	128	423	129	424
rect	129	423	130	424
rect	130	423	131	424
rect	131	423	132	424
rect	132	423	133	424
rect	134	423	135	424
rect	135	423	136	424
rect	136	423	137	424
rect	137	423	138	424
rect	138	423	139	424
rect	139	423	140	424
rect	140	423	141	424
rect	141	423	142	424
rect	142	423	143	424
rect	143	423	144	424
rect	144	423	145	424
rect	145	423	146	424
rect	197	423	198	424
rect	198	423	199	424
rect	199	423	200	424
rect	210	423	211	424
rect	211	423	212	424
rect	219	423	220	424
rect	220	423	221	424
rect	222	423	223	424
rect	223	423	224	424
rect	225	423	226	424
rect	226	423	227	424
rect	227	423	228	424
rect	228	423	229	424
rect	229	423	230	424
rect	230	423	231	424
rect	232	423	233	424
rect	233	423	234	424
rect	234	423	235	424
rect	235	423	236	424
rect	236	423	237	424
rect	238	423	239	424
rect	239	423	240	424
rect	240	423	241	424
rect	241	423	242	424
rect	242	423	243	424
rect	243	423	244	424
rect	244	423	245	424
rect	245	423	246	424
rect	246	423	247	424
rect	248	423	249	424
rect	249	423	250	424
rect	250	423	251	424
rect	258	423	259	424
rect	259	423	260	424
rect	279	423	280	424
rect	280	423	281	424
rect	282	423	283	424
rect	283	423	284	424
rect	288	423	289	424
rect	289	423	290	424
rect	290	423	291	424
rect	291	423	292	424
rect	292	423	293	424
rect	101	425	102	426
rect	102	425	103	426
rect	103	425	104	426
rect	104	425	105	426
rect	105	425	106	426
rect	106	425	107	426
rect	108	425	109	426
rect	109	425	110	426
rect	121	425	122	426
rect	122	425	123	426
rect	123	425	124	426
rect	125	425	126	426
rect	126	425	127	426
rect	128	425	129	426
rect	129	425	130	426
rect	130	425	131	426
rect	131	425	132	426
rect	132	425	133	426
rect	134	425	135	426
rect	135	425	136	426
rect	136	425	137	426
rect	137	425	138	426
rect	138	425	139	426
rect	139	425	140	426
rect	140	425	141	426
rect	141	425	142	426
rect	142	425	143	426
rect	143	425	144	426
rect	144	425	145	426
rect	145	425	146	426
rect	146	425	147	426
rect	147	425	148	426
rect	148	425	149	426
rect	149	425	150	426
rect	150	425	151	426
rect	151	425	152	426
rect	152	425	153	426
rect	153	425	154	426
rect	154	425	155	426
rect	155	425	156	426
rect	156	425	157	426
rect	157	425	158	426
rect	158	425	159	426
rect	159	425	160	426
rect	160	425	161	426
rect	161	425	162	426
rect	162	425	163	426
rect	163	425	164	426
rect	164	425	165	426
rect	165	425	166	426
rect	166	425	167	426
rect	167	425	168	426
rect	168	425	169	426
rect	169	425	170	426
rect	170	425	171	426
rect	171	425	172	426
rect	172	425	173	426
rect	173	425	174	426
rect	174	425	175	426
rect	175	425	176	426
rect	176	425	177	426
rect	177	425	178	426
rect	178	425	179	426
rect	179	425	180	426
rect	180	425	181	426
rect	181	425	182	426
rect	182	425	183	426
rect	183	425	184	426
rect	184	425	185	426
rect	185	425	186	426
rect	187	425	188	426
rect	188	425	189	426
rect	189	425	190	426
rect	190	425	191	426
rect	191	425	192	426
rect	192	425	193	426
rect	193	425	194	426
rect	194	425	195	426
rect	195	425	196	426
rect	197	425	198	426
rect	198	425	199	426
rect	199	425	200	426
rect	200	425	201	426
rect	201	425	202	426
rect	202	425	203	426
rect	203	425	204	426
rect	204	425	205	426
rect	206	425	207	426
rect	207	425	208	426
rect	208	425	209	426
rect	209	425	210	426
rect	210	425	211	426
rect	211	425	212	426
rect	212	425	213	426
rect	213	425	214	426
rect	214	425	215	426
rect	215	425	216	426
rect	216	425	217	426
rect	217	425	218	426
rect	219	425	220	426
rect	220	425	221	426
rect	222	425	223	426
rect	223	425	224	426
rect	225	425	226	426
rect	226	425	227	426
rect	227	425	228	426
rect	228	425	229	426
rect	229	425	230	426
rect	230	425	231	426
rect	232	425	233	426
rect	233	425	234	426
rect	234	425	235	426
rect	235	425	236	426
rect	236	425	237	426
rect	238	425	239	426
rect	239	425	240	426
rect	240	425	241	426
rect	241	425	242	426
rect	242	425	243	426
rect	243	425	244	426
rect	244	425	245	426
rect	245	425	246	426
rect	246	425	247	426
rect	248	425	249	426
rect	249	425	250	426
rect	250	425	251	426
rect	251	425	252	426
rect	252	425	253	426
rect	254	425	255	426
rect	255	425	256	426
rect	256	425	257	426
rect	257	425	258	426
rect	258	425	259	426
rect	259	425	260	426
rect	260	425	261	426
rect	261	425	262	426
rect	263	425	264	426
rect	264	425	265	426
rect	266	425	267	426
rect	267	425	268	426
rect	269	425	270	426
rect	270	425	271	426
rect	271	425	272	426
rect	272	425	273	426
rect	273	425	274	426
rect	274	425	275	426
rect	275	425	276	426
rect	276	425	277	426
rect	277	425	278	426
rect	278	425	279	426
rect	279	425	280	426
rect	280	425	281	426
rect	282	425	283	426
rect	283	425	284	426
rect	284	425	285	426
rect	285	425	286	426
rect	286	425	287	426
rect	287	425	288	426
rect	288	425	289	426
rect	289	425	290	426
rect	290	425	291	426
rect	291	425	292	426
rect	292	425	293	426
rect	293	425	294	426
rect	294	425	295	426
rect	295	425	296	426
rect	296	425	297	426
rect	297	425	298	426
rect	298	425	299	426
rect	299	425	300	426
rect	300	425	301	426
rect	301	425	302	426
rect	302	425	303	426
rect	303	425	304	426
rect	304	425	305	426
rect	305	425	306	426
rect	306	425	307	426
rect	307	425	308	426
rect	308	425	309	426
rect	309	425	310	426
rect	310	425	311	426
rect	311	425	312	426
rect	312	425	313	426
rect	313	425	314	426
rect	314	425	315	426
rect	315	425	316	426
rect	316	425	317	426
rect	317	425	318	426
rect	318	425	319	426
rect	319	425	320	426
rect	320	425	321	426
rect	321	425	322	426
rect	322	425	323	426
rect	323	425	324	426
rect	324	425	325	426
rect	325	425	326	426
rect	326	425	327	426
rect	327	425	328	426
rect	58	427	59	428
rect	59	427	60	428
rect	60	427	61	428
rect	61	427	62	428
rect	62	427	63	428
rect	102	427	103	428
rect	103	427	104	428
rect	104	427	105	428
rect	105	427	106	428
rect	106	427	107	428
rect	108	427	109	428
rect	109	427	110	428
rect	111	427	112	428
rect	112	427	113	428
rect	114	427	115	428
rect	115	427	116	428
rect	116	427	117	428
rect	117	427	118	428
rect	118	427	119	428
rect	119	427	120	428
rect	121	427	122	428
rect	122	427	123	428
rect	123	427	124	428
rect	128	427	129	428
rect	129	427	130	428
rect	130	427	131	428
rect	131	427	132	428
rect	132	427	133	428
rect	191	427	192	428
rect	192	427	193	428
rect	193	427	194	428
rect	194	427	195	428
rect	195	427	196	428
rect	197	427	198	428
rect	198	427	199	428
rect	199	427	200	428
rect	200	427	201	428
rect	201	427	202	428
rect	202	427	203	428
rect	203	427	204	428
rect	204	427	205	428
rect	206	427	207	428
rect	207	427	208	428
rect	208	427	209	428
rect	209	427	210	428
rect	210	427	211	428
rect	211	427	212	428
rect	212	427	213	428
rect	213	427	214	428
rect	214	427	215	428
rect	215	427	216	428
rect	216	427	217	428
rect	217	427	218	428
rect	219	427	220	428
rect	220	427	221	428
rect	222	427	223	428
rect	223	427	224	428
rect	225	427	226	428
rect	226	427	227	428
rect	227	427	228	428
rect	228	427	229	428
rect	229	427	230	428
rect	230	427	231	428
rect	232	427	233	428
rect	233	427	234	428
rect	234	427	235	428
rect	235	427	236	428
rect	236	427	237	428
rect	238	427	239	428
rect	239	427	240	428
rect	240	427	241	428
rect	241	427	242	428
rect	242	427	243	428
rect	243	427	244	428
rect	244	427	245	428
rect	245	427	246	428
rect	246	427	247	428
rect	248	427	249	428
rect	249	427	250	428
rect	250	427	251	428
rect	251	427	252	428
rect	252	427	253	428
rect	254	427	255	428
rect	255	427	256	428
rect	256	427	257	428
rect	257	427	258	428
rect	258	427	259	428
rect	259	427	260	428
rect	260	427	261	428
rect	261	427	262	428
rect	263	427	264	428
rect	264	427	265	428
rect	266	427	267	428
rect	267	427	268	428
rect	269	427	270	428
rect	270	427	271	428
rect	271	427	272	428
rect	272	427	273	428
rect	273	427	274	428
rect	274	427	275	428
rect	275	427	276	428
rect	276	427	277	428
rect	277	427	278	428
rect	278	427	279	428
rect	279	427	280	428
rect	280	427	281	428
rect	282	427	283	428
rect	283	427	284	428
rect	284	427	285	428
rect	285	427	286	428
rect	286	427	287	428
rect	287	427	288	428
rect	288	427	289	428
rect	289	427	290	428
rect	290	427	291	428
rect	291	427	292	428
rect	292	427	293	428
rect	293	427	294	428
rect	294	427	295	428
rect	295	427	296	428
rect	296	427	297	428
rect	297	427	298	428
rect	298	427	299	428
rect	299	427	300	428
rect	300	427	301	428
rect	301	427	302	428
rect	302	427	303	428
rect	303	427	304	428
rect	304	427	305	428
rect	305	427	306	428
rect	306	427	307	428
rect	307	427	308	428
rect	308	427	309	428
rect	309	427	310	428
rect	310	427	311	428
rect	311	427	312	428
rect	312	427	313	428
rect	313	427	314	428
rect	314	427	315	428
rect	315	427	316	428
rect	316	427	317	428
rect	317	427	318	428
rect	318	427	319	428
rect	319	427	320	428
rect	320	427	321	428
rect	321	427	322	428
rect	322	427	323	428
rect	323	427	324	428
rect	324	427	325	428
rect	325	427	326	428
rect	326	427	327	428
rect	327	427	328	428
rect	328	427	329	428
rect	329	427	330	428
rect	330	427	331	428
rect	72	436	73	437
rect	73	436	74	437
rect	74	436	75	437
rect	75	436	76	437
rect	76	436	77	437
rect	78	436	79	437
rect	79	436	80	437
rect	82	438	83	439
rect	83	438	84	439
rect	84	438	85	439
rect	85	438	86	439
rect	87	438	88	439
rect	88	438	89	439
rect	90	438	91	439
rect	91	438	92	439
rect	92	438	93	439
rect	93	438	94	439
rect	94	438	95	439
rect	96	438	97	439
rect	97	438	98	439
rect	99	438	100	439
rect	100	438	101	439
rect	101	438	102	439
rect	102	438	103	439
rect	103	438	104	439
rect	104	438	105	439
rect	105	438	106	439
rect	106	438	107	439
rect	108	438	109	439
rect	109	438	110	439
rect	111	438	112	439
rect	112	438	113	439
rect	113	438	114	439
rect	114	438	115	439
rect	115	438	116	439
rect	117	438	118	439
rect	118	438	119	439
rect	119	438	120	439
rect	120	438	121	439
rect	121	438	122	439
rect	122	438	123	439
rect	123	438	124	439
rect	124	438	125	439
rect	125	438	126	439
rect	126	438	127	439
rect	127	438	128	439
rect	128	438	129	439
rect	129	438	130	439
rect	130	438	131	439
rect	131	438	132	439
rect	132	438	133	439
rect	133	438	134	439
rect	134	438	135	439
rect	135	438	136	439
rect	136	438	137	439
rect	137	438	138	439
rect	138	438	139	439
rect	139	438	140	439
rect	140	438	141	439
rect	141	438	142	439
rect	142	438	143	439
rect	143	438	144	439
rect	144	438	145	439
rect	145	438	146	439
rect	146	438	147	439
rect	147	438	148	439
rect	148	438	149	439
rect	149	438	150	439
rect	150	438	151	439
rect	151	438	152	439
rect	152	438	153	439
rect	153	438	154	439
rect	154	438	155	439
rect	155	438	156	439
rect	156	438	157	439
rect	157	438	158	439
rect	158	438	159	439
rect	159	438	160	439
rect	160	438	161	439
rect	161	438	162	439
rect	162	438	163	439
rect	163	438	164	439
rect	164	438	165	439
rect	165	438	166	439
rect	166	438	167	439
rect	78	440	79	441
rect	79	440	80	441
rect	80	440	81	441
rect	82	440	83	441
rect	83	440	84	441
rect	84	440	85	441
rect	85	440	86	441
rect	99	440	100	441
rect	100	440	101	441
rect	111	440	112	441
rect	112	440	113	441
rect	113	440	114	441
rect	114	440	115	441
rect	115	440	116	441
rect	117	440	118	441
rect	118	440	119	441
rect	119	440	120	441
rect	120	440	121	441
rect	121	440	122	441
rect	122	440	123	441
rect	123	440	124	441
rect	124	440	125	441
rect	125	440	126	441
rect	126	440	127	441
rect	127	440	128	441
rect	128	440	129	441
rect	129	440	130	441
rect	130	440	131	441
rect	131	440	132	441
rect	132	440	133	441
rect	133	440	134	441
rect	134	440	135	441
rect	135	440	136	441
rect	136	440	137	441
rect	137	440	138	441
rect	138	440	139	441
rect	139	440	140	441
rect	140	440	141	441
rect	141	440	142	441
rect	142	440	143	441
rect	143	440	144	441
rect	144	440	145	441
rect	145	440	146	441
rect	146	440	147	441
rect	147	440	148	441
rect	148	440	149	441
rect	149	440	150	441
rect	150	440	151	441
rect	151	440	152	441
rect	152	440	153	441
rect	153	440	154	441
rect	154	440	155	441
rect	155	440	156	441
rect	156	440	157	441
rect	157	440	158	441
rect	158	440	159	441
rect	159	440	160	441
rect	160	440	161	441
rect	161	440	162	441
rect	162	440	163	441
rect	163	440	164	441
rect	164	440	165	441
rect	165	440	166	441
rect	166	440	167	441
rect	168	440	169	441
rect	169	440	170	441
rect	170	440	171	441
rect	171	440	172	441
rect	172	440	173	441
rect	173	440	174	441
rect	174	440	175	441
rect	175	440	176	441
rect	176	440	177	441
rect	177	440	178	441
rect	178	440	179	441
rect	179	440	180	441
rect	180	440	181	441
rect	181	440	182	441
rect	182	440	183	441
rect	183	440	184	441
rect	184	440	185	441
rect	185	440	186	441
rect	186	440	187	441
rect	187	440	188	441
rect	188	440	189	441
rect	189	440	190	441
rect	190	440	191	441
rect	191	440	192	441
rect	192	440	193	441
rect	193	440	194	441
rect	194	440	195	441
rect	195	440	196	441
rect	197	440	198	441
rect	198	440	199	441
rect	199	440	200	441
rect	200	440	201	441
rect	201	440	202	441
rect	203	440	204	441
rect	204	440	205	441
rect	206	440	207	441
rect	207	440	208	441
rect	208	440	209	441
rect	209	440	210	441
rect	210	440	211	441
rect	211	440	212	441
rect	212	440	213	441
rect	213	440	214	441
rect	214	440	215	441
rect	215	440	216	441
rect	216	440	217	441
rect	217	440	218	441
rect	219	440	220	441
rect	220	440	221	441
rect	222	440	223	441
rect	223	440	224	441
rect	251	440	252	441
rect	252	440	253	441
rect	254	440	255	441
rect	255	440	256	441
rect	256	440	257	441
rect	257	440	258	441
rect	258	440	259	441
rect	260	440	261	441
rect	261	440	262	441
rect	263	440	264	441
rect	264	440	265	441
rect	79	442	80	443
rect	80	442	81	443
rect	82	442	83	443
rect	83	442	84	443
rect	84	442	85	443
rect	85	442	86	443
rect	86	442	87	443
rect	87	442	88	443
rect	88	442	89	443
rect	96	442	97	443
rect	97	442	98	443
rect	98	442	99	443
rect	99	442	100	443
rect	100	442	101	443
rect	102	442	103	443
rect	103	442	104	443
rect	104	442	105	443
rect	105	442	106	443
rect	106	442	107	443
rect	108	442	109	443
rect	109	442	110	443
rect	110	442	111	443
rect	111	442	112	443
rect	112	442	113	443
rect	113	442	114	443
rect	114	442	115	443
rect	115	442	116	443
rect	117	442	118	443
rect	118	442	119	443
rect	119	442	120	443
rect	120	442	121	443
rect	121	442	122	443
rect	122	442	123	443
rect	123	442	124	443
rect	124	442	125	443
rect	125	442	126	443
rect	126	442	127	443
rect	127	442	128	443
rect	128	442	129	443
rect	129	442	130	443
rect	130	442	131	443
rect	131	442	132	443
rect	132	442	133	443
rect	133	442	134	443
rect	134	442	135	443
rect	135	442	136	443
rect	136	442	137	443
rect	137	442	138	443
rect	138	442	139	443
rect	139	442	140	443
rect	140	442	141	443
rect	141	442	142	443
rect	142	442	143	443
rect	143	442	144	443
rect	144	442	145	443
rect	145	442	146	443
rect	146	442	147	443
rect	147	442	148	443
rect	148	442	149	443
rect	149	442	150	443
rect	150	442	151	443
rect	151	442	152	443
rect	152	442	153	443
rect	153	442	154	443
rect	154	442	155	443
rect	155	442	156	443
rect	156	442	157	443
rect	157	442	158	443
rect	158	442	159	443
rect	159	442	160	443
rect	160	442	161	443
rect	161	442	162	443
rect	162	442	163	443
rect	163	442	164	443
rect	164	442	165	443
rect	165	442	166	443
rect	166	442	167	443
rect	168	442	169	443
rect	169	442	170	443
rect	170	442	171	443
rect	171	442	172	443
rect	172	442	173	443
rect	173	442	174	443
rect	174	442	175	443
rect	175	442	176	443
rect	176	442	177	443
rect	177	442	178	443
rect	178	442	179	443
rect	179	442	180	443
rect	180	442	181	443
rect	181	442	182	443
rect	182	442	183	443
rect	183	442	184	443
rect	184	442	185	443
rect	185	442	186	443
rect	186	442	187	443
rect	187	442	188	443
rect	188	442	189	443
rect	189	442	190	443
rect	190	442	191	443
rect	191	442	192	443
rect	192	442	193	443
rect	193	442	194	443
rect	194	442	195	443
rect	195	442	196	443
rect	232	442	233	443
rect	233	442	234	443
rect	234	442	235	443
rect	235	442	236	443
rect	236	442	237	443
rect	248	442	249	443
rect	249	442	250	443
rect	250	442	251	443
rect	251	442	252	443
rect	252	442	253	443
rect	260	442	261	443
rect	261	442	262	443
rect	33	444	34	445
rect	34	444	35	445
rect	35	444	36	445
rect	36	444	37	445
rect	37	444	38	445
rect	38	444	39	445
rect	39	444	40	445
rect	40	444	41	445
rect	41	444	42	445
rect	42	444	43	445
rect	43	444	44	445
rect	44	444	45	445
rect	45	444	46	445
rect	46	444	47	445
rect	47	444	48	445
rect	48	444	49	445
rect	49	444	50	445
rect	50	444	51	445
rect	51	444	52	445
rect	52	444	53	445
rect	53	444	54	445
rect	54	444	55	445
rect	55	444	56	445
rect	56	444	57	445
rect	57	444	58	445
rect	58	444	59	445
rect	59	444	60	445
rect	60	444	61	445
rect	61	444	62	445
rect	62	444	63	445
rect	63	444	64	445
rect	64	444	65	445
rect	65	444	66	445
rect	66	444	67	445
rect	67	444	68	445
rect	68	444	69	445
rect	69	444	70	445
rect	70	444	71	445
rect	71	444	72	445
rect	72	444	73	445
rect	73	444	74	445
rect	74	444	75	445
rect	75	444	76	445
rect	76	444	77	445
rect	77	444	78	445
rect	79	444	80	445
rect	80	444	81	445
rect	82	444	83	445
rect	83	444	84	445
rect	84	444	85	445
rect	85	444	86	445
rect	86	444	87	445
rect	87	444	88	445
rect	88	444	89	445
rect	89	444	90	445
rect	90	444	91	445
rect	91	444	92	445
rect	92	444	93	445
rect	93	444	94	445
rect	94	444	95	445
rect	95	444	96	445
rect	96	444	97	445
rect	97	444	98	445
rect	108	444	109	445
rect	109	444	110	445
rect	110	444	111	445
rect	111	444	112	445
rect	112	444	113	445
rect	113	444	114	445
rect	114	444	115	445
rect	115	444	116	445
rect	203	444	204	445
rect	204	444	205	445
rect	219	444	220	445
rect	220	444	221	445
rect	228	444	229	445
rect	229	444	230	445
rect	230	444	231	445
rect	231	444	232	445
rect	232	444	233	445
rect	233	444	234	445
rect	234	444	235	445
rect	235	444	236	445
rect	236	444	237	445
rect	237	444	238	445
rect	238	444	239	445
rect	239	444	240	445
rect	240	444	241	445
rect	241	444	242	445
rect	242	444	243	445
rect	243	444	244	445
rect	244	444	245	445
rect	245	444	246	445
rect	246	444	247	445
rect	247	444	248	445
rect	248	444	249	445
rect	249	444	250	445
rect	250	444	251	445
rect	251	444	252	445
rect	252	444	253	445
rect	253	444	254	445
rect	254	444	255	445
rect	255	444	256	445
rect	256	444	257	445
rect	257	444	258	445
rect	258	444	259	445
rect	259	444	260	445
rect	260	444	261	445
rect	261	444	262	445
rect	262	444	263	445
rect	263	444	264	445
rect	264	444	265	445
rect	265	444	266	445
rect	266	444	267	445
rect	267	444	268	445
rect	268	444	269	445
rect	269	444	270	445
rect	270	444	271	445
rect	271	444	272	445
rect	272	444	273	445
rect	273	444	274	445
rect	274	444	275	445
rect	275	444	276	445
rect	276	444	277	445
rect	277	444	278	445
rect	278	444	279	445
rect	279	444	280	445
rect	280	444	281	445
rect	102	453	103	454
rect	103	453	104	454
rect	105	453	106	454
rect	106	453	107	454
rect	99	455	100	456
rect	100	455	101	456
rect	101	455	102	456
rect	102	455	103	456
rect	103	455	104	456
<< metal2 >>
rect	69	1	70	2
rect	72	1	73	2
rect	69	2	70	3
rect	72	2	73	3
rect	56	3	57	4
rect	69	3	70	4
rect	72	3	73	4
rect	131	3	132	4
rect	190	3	191	4
rect	193	3	194	4
rect	56	4	57	5
rect	69	4	70	5
rect	72	4	73	5
rect	131	4	132	5
rect	190	4	191	5
rect	193	4	194	5
rect	43	5	44	6
rect	56	5	57	6
rect	69	5	70	6
rect	72	5	73	6
rect	109	5	110	6
rect	118	5	119	6
rect	124	5	125	6
rect	131	5	132	6
rect	173	5	174	6
rect	190	5	191	6
rect	193	5	194	6
rect	220	5	221	6
rect	237	5	238	6
rect	243	5	244	6
rect	246	5	247	6
rect	252	5	253	6
rect	262	5	263	6
rect	265	5	266	6
rect	11	12	12	13
rect	29	12	30	13
rect	32	12	33	13
rect	53	12	54	13
rect	56	12	57	13
rect	72	12	73	13
rect	85	12	86	13
rect	109	12	110	13
rect	118	12	119	13
rect	131	12	132	13
rect	142	12	143	13
rect	163	12	164	13
rect	170	12	171	13
rect	177	12	178	13
rect	180	12	181	13
rect	190	12	191	13
rect	200	12	201	13
rect	214	12	215	13
rect	220	12	221	13
rect	243	12	244	13
rect	246	12	247	13
rect	252	12	253	13
rect	262	12	263	13
rect	11	13	12	14
rect	29	13	30	14
rect	53	13	54	14
rect	56	13	57	14
rect	72	13	73	14
rect	85	13	86	14
rect	109	13	110	14
rect	118	13	119	14
rect	131	13	132	14
rect	142	13	143	14
rect	163	13	164	14
rect	170	13	171	14
rect	177	13	178	14
rect	180	13	181	14
rect	190	13	191	14
rect	200	13	201	14
rect	214	13	215	14
rect	220	13	221	14
rect	243	13	244	14
rect	246	13	247	14
rect	262	13	263	14
rect	11	14	12	15
rect	29	14	30	15
rect	53	14	54	15
rect	56	14	57	15
rect	72	14	73	15
rect	85	14	86	15
rect	109	14	110	15
rect	118	14	119	15
rect	131	14	132	15
rect	142	14	143	15
rect	163	14	164	15
rect	170	14	171	15
rect	177	14	178	15
rect	180	14	181	15
rect	190	14	191	15
rect	200	14	201	15
rect	214	14	215	15
rect	220	14	221	15
rect	243	14	244	15
rect	246	14	247	15
rect	262	14	263	15
rect	11	15	12	16
rect	29	15	30	16
rect	53	15	54	16
rect	56	15	57	16
rect	72	15	73	16
rect	85	15	86	16
rect	109	15	110	16
rect	118	15	119	16
rect	131	15	132	16
rect	142	15	143	16
rect	163	15	164	16
rect	170	15	171	16
rect	177	15	178	16
rect	200	15	201	16
rect	214	15	215	16
rect	220	15	221	16
rect	243	15	244	16
rect	262	15	263	16
rect	11	16	12	17
rect	29	16	30	17
rect	53	16	54	17
rect	56	16	57	17
rect	72	16	73	17
rect	85	16	86	17
rect	109	16	110	17
rect	118	16	119	17
rect	131	16	132	17
rect	142	16	143	17
rect	163	16	164	17
rect	170	16	171	17
rect	177	16	178	17
rect	182	16	183	17
rect	191	16	192	17
rect	200	16	201	17
rect	214	16	215	17
rect	220	16	221	17
rect	243	16	244	17
rect	253	16	254	17
rect	262	16	263	17
rect	11	17	12	18
rect	29	17	30	18
rect	53	17	54	18
rect	56	17	57	18
rect	72	17	73	18
rect	85	17	86	18
rect	118	17	119	18
rect	131	17	132	18
rect	142	17	143	18
rect	163	17	164	18
rect	170	17	171	18
rect	177	17	178	18
rect	182	17	183	18
rect	191	17	192	18
rect	214	17	215	18
rect	253	17	254	18
rect	262	17	263	18
rect	11	18	12	19
rect	29	18	30	19
rect	53	18	54	19
rect	56	18	57	19
rect	72	18	73	19
rect	85	18	86	19
rect	108	18	109	19
rect	118	18	119	19
rect	131	18	132	19
rect	142	18	143	19
rect	163	18	164	19
rect	170	18	171	19
rect	177	18	178	19
rect	179	18	180	19
rect	182	18	183	19
rect	191	18	192	19
rect	214	18	215	19
rect	221	18	222	19
rect	253	18	254	19
rect	262	18	263	19
rect	265	18	266	19
rect	11	19	12	20
rect	29	19	30	20
rect	53	19	54	20
rect	56	19	57	20
rect	72	19	73	20
rect	85	19	86	20
rect	108	19	109	20
rect	131	19	132	20
rect	142	19	143	20
rect	163	19	164	20
rect	179	19	180	20
rect	182	19	183	20
rect	191	19	192	20
rect	214	19	215	20
rect	221	19	222	20
rect	253	19	254	20
rect	262	19	263	20
rect	265	19	266	20
rect	11	20	12	21
rect	29	20	30	21
rect	53	20	54	21
rect	56	20	57	21
rect	72	20	73	21
rect	85	20	86	21
rect	95	20	96	21
rect	108	20	109	21
rect	131	20	132	21
rect	142	20	143	21
rect	163	20	164	21
rect	167	20	168	21
rect	179	20	180	21
rect	182	20	183	21
rect	191	20	192	21
rect	200	20	201	21
rect	209	20	210	21
rect	214	20	215	21
rect	221	20	222	21
rect	253	20	254	21
rect	262	20	263	21
rect	265	20	266	21
rect	278	20	279	21
rect	11	21	12	22
rect	29	21	30	22
rect	95	21	96	22
rect	108	21	109	22
rect	142	21	143	22
rect	167	21	168	22
rect	179	21	180	22
rect	182	21	183	22
rect	191	21	192	22
rect	200	21	201	22
rect	209	21	210	22
rect	214	21	215	22
rect	221	21	222	22
rect	253	21	254	22
rect	262	21	263	22
rect	265	21	266	22
rect	278	21	279	22
rect	11	22	12	23
rect	29	22	30	23
rect	71	22	72	23
rect	95	22	96	23
rect	108	22	109	23
rect	142	22	143	23
rect	167	22	168	23
rect	179	22	180	23
rect	182	22	183	23
rect	191	22	192	23
rect	200	22	201	23
rect	209	22	210	23
rect	214	22	215	23
rect	221	22	222	23
rect	253	22	254	23
rect	256	22	257	23
rect	262	22	263	23
rect	265	22	266	23
rect	278	22	279	23
rect	285	22	286	23
rect	302	22	303	23
rect	71	23	72	24
rect	95	23	96	24
rect	108	23	109	24
rect	167	23	168	24
rect	179	23	180	24
rect	182	23	183	24
rect	191	23	192	24
rect	200	23	201	24
rect	209	23	210	24
rect	221	23	222	24
rect	253	23	254	24
rect	256	23	257	24
rect	265	23	266	24
rect	278	23	279	24
rect	285	23	286	24
rect	302	23	303	24
rect	14	24	15	25
rect	30	24	31	25
rect	50	24	51	25
rect	53	24	54	25
rect	62	24	63	25
rect	71	24	72	25
rect	95	24	96	25
rect	108	24	109	25
rect	125	24	126	25
rect	152	24	153	25
rect	161	24	162	25
rect	167	24	168	25
rect	179	24	180	25
rect	182	24	183	25
rect	191	24	192	25
rect	200	24	201	25
rect	209	24	210	25
rect	218	24	219	25
rect	221	24	222	25
rect	227	24	228	25
rect	244	24	245	25
rect	247	24	248	25
rect	253	24	254	25
rect	256	24	257	25
rect	265	24	266	25
rect	278	24	279	25
rect	285	24	286	25
rect	296	24	297	25
rect	302	24	303	25
rect	14	25	15	26
rect	30	25	31	26
rect	50	25	51	26
rect	53	25	54	26
rect	62	25	63	26
rect	71	25	72	26
rect	95	25	96	26
rect	108	25	109	26
rect	125	25	126	26
rect	152	25	153	26
rect	161	25	162	26
rect	167	25	168	26
rect	179	25	180	26
rect	182	25	183	26
rect	191	25	192	26
rect	200	25	201	26
rect	209	25	210	26
rect	218	25	219	26
rect	221	25	222	26
rect	227	25	228	26
rect	244	25	245	26
rect	247	25	248	26
rect	253	25	254	26
rect	256	25	257	26
rect	265	25	266	26
rect	278	25	279	26
rect	285	25	286	26
rect	296	25	297	26
rect	302	25	303	26
rect	11	26	12	27
rect	14	26	15	27
rect	30	26	31	27
rect	50	26	51	27
rect	53	26	54	27
rect	62	26	63	27
rect	71	26	72	27
rect	95	26	96	27
rect	108	26	109	27
rect	125	26	126	27
rect	152	26	153	27
rect	161	26	162	27
rect	164	26	165	27
rect	167	26	168	27
rect	170	26	171	27
rect	176	26	177	27
rect	179	26	180	27
rect	182	26	183	27
rect	188	26	189	27
rect	191	26	192	27
rect	200	26	201	27
rect	209	26	210	27
rect	218	26	219	27
rect	221	26	222	27
rect	227	26	228	27
rect	244	26	245	27
rect	247	26	248	27
rect	253	26	254	27
rect	256	26	257	27
rect	265	26	266	27
rect	278	26	279	27
rect	285	26	286	27
rect	296	26	297	27
rect	302	26	303	27
rect	305	26	306	27
rect	14	33	15	34
rect	30	33	31	34
rect	47	33	48	34
rect	53	33	54	34
rect	56	33	57	34
rect	62	33	63	34
rect	71	33	72	34
rect	77	33	78	34
rect	108	33	109	34
rect	114	33	115	34
rect	146	33	147	34
rect	149	33	150	34
rect	152	33	153	34
rect	161	33	162	34
rect	164	33	165	34
rect	167	33	168	34
rect	173	33	174	34
rect	176	33	177	34
rect	179	33	180	34
rect	182	33	183	34
rect	191	33	192	34
rect	194	33	195	34
rect	197	33	198	34
rect	200	33	201	34
rect	203	33	204	34
rect	209	33	210	34
rect	218	33	219	34
rect	221	33	222	34
rect	231	33	232	34
rect	244	33	245	34
rect	250	33	251	34
rect	253	33	254	34
rect	256	33	257	34
rect	265	33	266	34
rect	278	33	279	34
rect	302	33	303	34
rect	305	33	306	34
rect	14	34	15	35
rect	30	34	31	35
rect	47	34	48	35
rect	53	34	54	35
rect	56	34	57	35
rect	62	34	63	35
rect	71	34	72	35
rect	77	34	78	35
rect	108	34	109	35
rect	114	34	115	35
rect	146	34	147	35
rect	149	34	150	35
rect	152	34	153	35
rect	161	34	162	35
rect	164	34	165	35
rect	167	34	168	35
rect	173	34	174	35
rect	176	34	177	35
rect	179	34	180	35
rect	182	34	183	35
rect	191	34	192	35
rect	194	34	195	35
rect	197	34	198	35
rect	200	34	201	35
rect	203	34	204	35
rect	209	34	210	35
rect	221	34	222	35
rect	231	34	232	35
rect	244	34	245	35
rect	250	34	251	35
rect	253	34	254	35
rect	256	34	257	35
rect	265	34	266	35
rect	278	34	279	35
rect	302	34	303	35
rect	305	34	306	35
rect	14	35	15	36
rect	30	35	31	36
rect	47	35	48	36
rect	53	35	54	36
rect	56	35	57	36
rect	62	35	63	36
rect	71	35	72	36
rect	77	35	78	36
rect	108	35	109	36
rect	114	35	115	36
rect	146	35	147	36
rect	149	35	150	36
rect	152	35	153	36
rect	161	35	162	36
rect	164	35	165	36
rect	167	35	168	36
rect	173	35	174	36
rect	176	35	177	36
rect	179	35	180	36
rect	182	35	183	36
rect	191	35	192	36
rect	194	35	195	36
rect	197	35	198	36
rect	200	35	201	36
rect	203	35	204	36
rect	209	35	210	36
rect	215	35	216	36
rect	221	35	222	36
rect	231	35	232	36
rect	244	35	245	36
rect	250	35	251	36
rect	253	35	254	36
rect	256	35	257	36
rect	265	35	266	36
rect	278	35	279	36
rect	302	35	303	36
rect	305	35	306	36
rect	14	36	15	37
rect	30	36	31	37
rect	47	36	48	37
rect	53	36	54	37
rect	56	36	57	37
rect	62	36	63	37
rect	71	36	72	37
rect	77	36	78	37
rect	108	36	109	37
rect	114	36	115	37
rect	146	36	147	37
rect	149	36	150	37
rect	152	36	153	37
rect	161	36	162	37
rect	164	36	165	37
rect	167	36	168	37
rect	173	36	174	37
rect	176	36	177	37
rect	179	36	180	37
rect	182	36	183	37
rect	191	36	192	37
rect	194	36	195	37
rect	197	36	198	37
rect	200	36	201	37
rect	209	36	210	37
rect	215	36	216	37
rect	221	36	222	37
rect	231	36	232	37
rect	244	36	245	37
rect	250	36	251	37
rect	253	36	254	37
rect	256	36	257	37
rect	265	36	266	37
rect	278	36	279	37
rect	302	36	303	37
rect	305	36	306	37
rect	14	37	15	38
rect	30	37	31	38
rect	47	37	48	38
rect	53	37	54	38
rect	56	37	57	38
rect	62	37	63	38
rect	71	37	72	38
rect	77	37	78	38
rect	108	37	109	38
rect	114	37	115	38
rect	146	37	147	38
rect	149	37	150	38
rect	152	37	153	38
rect	161	37	162	38
rect	164	37	165	38
rect	167	37	168	38
rect	173	37	174	38
rect	176	37	177	38
rect	179	37	180	38
rect	182	37	183	38
rect	191	37	192	38
rect	194	37	195	38
rect	197	37	198	38
rect	200	37	201	38
rect	209	37	210	38
rect	215	37	216	38
rect	218	37	219	38
rect	221	37	222	38
rect	231	37	232	38
rect	244	37	245	38
rect	250	37	251	38
rect	253	37	254	38
rect	256	37	257	38
rect	265	37	266	38
rect	278	37	279	38
rect	302	37	303	38
rect	305	37	306	38
rect	14	38	15	39
rect	30	38	31	39
rect	47	38	48	39
rect	53	38	54	39
rect	56	38	57	39
rect	62	38	63	39
rect	71	38	72	39
rect	77	38	78	39
rect	108	38	109	39
rect	114	38	115	39
rect	146	38	147	39
rect	149	38	150	39
rect	152	38	153	39
rect	161	38	162	39
rect	164	38	165	39
rect	167	38	168	39
rect	173	38	174	39
rect	176	38	177	39
rect	179	38	180	39
rect	182	38	183	39
rect	191	38	192	39
rect	194	38	195	39
rect	197	38	198	39
rect	209	38	210	39
rect	215	38	216	39
rect	218	38	219	39
rect	221	38	222	39
rect	231	38	232	39
rect	244	38	245	39
rect	250	38	251	39
rect	253	38	254	39
rect	256	38	257	39
rect	265	38	266	39
rect	278	38	279	39
rect	302	38	303	39
rect	305	38	306	39
rect	14	39	15	40
rect	30	39	31	40
rect	47	39	48	40
rect	53	39	54	40
rect	56	39	57	40
rect	62	39	63	40
rect	71	39	72	40
rect	77	39	78	40
rect	108	39	109	40
rect	114	39	115	40
rect	146	39	147	40
rect	149	39	150	40
rect	152	39	153	40
rect	161	39	162	40
rect	164	39	165	40
rect	167	39	168	40
rect	173	39	174	40
rect	176	39	177	40
rect	179	39	180	40
rect	182	39	183	40
rect	191	39	192	40
rect	194	39	195	40
rect	197	39	198	40
rect	203	39	204	40
rect	209	39	210	40
rect	215	39	216	40
rect	218	39	219	40
rect	221	39	222	40
rect	231	39	232	40
rect	244	39	245	40
rect	250	39	251	40
rect	253	39	254	40
rect	256	39	257	40
rect	265	39	266	40
rect	278	39	279	40
rect	302	39	303	40
rect	305	39	306	40
rect	14	40	15	41
rect	30	40	31	41
rect	47	40	48	41
rect	53	40	54	41
rect	56	40	57	41
rect	62	40	63	41
rect	71	40	72	41
rect	77	40	78	41
rect	108	40	109	41
rect	114	40	115	41
rect	146	40	147	41
rect	149	40	150	41
rect	152	40	153	41
rect	161	40	162	41
rect	164	40	165	41
rect	167	40	168	41
rect	173	40	174	41
rect	176	40	177	41
rect	179	40	180	41
rect	182	40	183	41
rect	191	40	192	41
rect	194	40	195	41
rect	203	40	204	41
rect	209	40	210	41
rect	215	40	216	41
rect	218	40	219	41
rect	221	40	222	41
rect	231	40	232	41
rect	244	40	245	41
rect	250	40	251	41
rect	253	40	254	41
rect	256	40	257	41
rect	265	40	266	41
rect	278	40	279	41
rect	302	40	303	41
rect	305	40	306	41
rect	14	41	15	42
rect	30	41	31	42
rect	47	41	48	42
rect	53	41	54	42
rect	56	41	57	42
rect	62	41	63	42
rect	71	41	72	42
rect	77	41	78	42
rect	108	41	109	42
rect	114	41	115	42
rect	146	41	147	42
rect	149	41	150	42
rect	152	41	153	42
rect	161	41	162	42
rect	164	41	165	42
rect	167	41	168	42
rect	173	41	174	42
rect	176	41	177	42
rect	179	41	180	42
rect	182	41	183	42
rect	191	41	192	42
rect	194	41	195	42
rect	203	41	204	42
rect	209	41	210	42
rect	215	41	216	42
rect	218	41	219	42
rect	221	41	222	42
rect	231	41	232	42
rect	244	41	245	42
rect	250	41	251	42
rect	253	41	254	42
rect	256	41	257	42
rect	265	41	266	42
rect	278	41	279	42
rect	302	41	303	42
rect	305	41	306	42
rect	309	41	310	42
rect	14	42	15	43
rect	30	42	31	43
rect	47	42	48	43
rect	53	42	54	43
rect	56	42	57	43
rect	62	42	63	43
rect	71	42	72	43
rect	77	42	78	43
rect	108	42	109	43
rect	114	42	115	43
rect	146	42	147	43
rect	149	42	150	43
rect	152	42	153	43
rect	161	42	162	43
rect	164	42	165	43
rect	167	42	168	43
rect	173	42	174	43
rect	179	42	180	43
rect	182	42	183	43
rect	191	42	192	43
rect	194	42	195	43
rect	203	42	204	43
rect	209	42	210	43
rect	215	42	216	43
rect	218	42	219	43
rect	221	42	222	43
rect	231	42	232	43
rect	244	42	245	43
rect	250	42	251	43
rect	253	42	254	43
rect	256	42	257	43
rect	278	42	279	43
rect	302	42	303	43
rect	305	42	306	43
rect	309	42	310	43
rect	14	43	15	44
rect	30	43	31	44
rect	47	43	48	44
rect	53	43	54	44
rect	56	43	57	44
rect	62	43	63	44
rect	71	43	72	44
rect	77	43	78	44
rect	108	43	109	44
rect	114	43	115	44
rect	146	43	147	44
rect	149	43	150	44
rect	152	43	153	44
rect	161	43	162	44
rect	164	43	165	44
rect	167	43	168	44
rect	173	43	174	44
rect	179	43	180	44
rect	182	43	183	44
rect	191	43	192	44
rect	194	43	195	44
rect	200	43	201	44
rect	203	43	204	44
rect	209	43	210	44
rect	215	43	216	44
rect	218	43	219	44
rect	221	43	222	44
rect	231	43	232	44
rect	244	43	245	44
rect	250	43	251	44
rect	253	43	254	44
rect	256	43	257	44
rect	276	43	277	44
rect	278	43	279	44
rect	302	43	303	44
rect	305	43	306	44
rect	309	43	310	44
rect	14	44	15	45
rect	30	44	31	45
rect	47	44	48	45
rect	53	44	54	45
rect	56	44	57	45
rect	62	44	63	45
rect	71	44	72	45
rect	77	44	78	45
rect	108	44	109	45
rect	114	44	115	45
rect	146	44	147	45
rect	149	44	150	45
rect	152	44	153	45
rect	161	44	162	45
rect	164	44	165	45
rect	167	44	168	45
rect	179	44	180	45
rect	182	44	183	45
rect	191	44	192	45
rect	194	44	195	45
rect	200	44	201	45
rect	203	44	204	45
rect	209	44	210	45
rect	215	44	216	45
rect	218	44	219	45
rect	221	44	222	45
rect	231	44	232	45
rect	244	44	245	45
rect	250	44	251	45
rect	253	44	254	45
rect	256	44	257	45
rect	276	44	277	45
rect	278	44	279	45
rect	302	44	303	45
rect	305	44	306	45
rect	309	44	310	45
rect	14	45	15	46
rect	30	45	31	46
rect	47	45	48	46
rect	53	45	54	46
rect	56	45	57	46
rect	62	45	63	46
rect	71	45	72	46
rect	77	45	78	46
rect	108	45	109	46
rect	114	45	115	46
rect	146	45	147	46
rect	149	45	150	46
rect	152	45	153	46
rect	161	45	162	46
rect	164	45	165	46
rect	167	45	168	46
rect	179	45	180	46
rect	182	45	183	46
rect	191	45	192	46
rect	194	45	195	46
rect	197	45	198	46
rect	200	45	201	46
rect	203	45	204	46
rect	209	45	210	46
rect	215	45	216	46
rect	218	45	219	46
rect	221	45	222	46
rect	231	45	232	46
rect	244	45	245	46
rect	250	45	251	46
rect	253	45	254	46
rect	256	45	257	46
rect	261	45	262	46
rect	273	45	274	46
rect	276	45	277	46
rect	278	45	279	46
rect	302	45	303	46
rect	305	45	306	46
rect	309	45	310	46
rect	14	46	15	47
rect	30	46	31	47
rect	47	46	48	47
rect	53	46	54	47
rect	56	46	57	47
rect	62	46	63	47
rect	71	46	72	47
rect	77	46	78	47
rect	108	46	109	47
rect	114	46	115	47
rect	146	46	147	47
rect	149	46	150	47
rect	152	46	153	47
rect	161	46	162	47
rect	164	46	165	47
rect	179	46	180	47
rect	182	46	183	47
rect	191	46	192	47
rect	194	46	195	47
rect	197	46	198	47
rect	200	46	201	47
rect	203	46	204	47
rect	209	46	210	47
rect	215	46	216	47
rect	218	46	219	47
rect	221	46	222	47
rect	244	46	245	47
rect	250	46	251	47
rect	253	46	254	47
rect	256	46	257	47
rect	261	46	262	47
rect	273	46	274	47
rect	276	46	277	47
rect	278	46	279	47
rect	302	46	303	47
rect	305	46	306	47
rect	309	46	310	47
rect	14	47	15	48
rect	30	47	31	48
rect	47	47	48	48
rect	53	47	54	48
rect	56	47	57	48
rect	62	47	63	48
rect	71	47	72	48
rect	77	47	78	48
rect	108	47	109	48
rect	114	47	115	48
rect	146	47	147	48
rect	149	47	150	48
rect	152	47	153	48
rect	161	47	162	48
rect	164	47	165	48
rect	176	47	177	48
rect	179	47	180	48
rect	182	47	183	48
rect	191	47	192	48
rect	194	47	195	48
rect	197	47	198	48
rect	200	47	201	48
rect	203	47	204	48
rect	209	47	210	48
rect	215	47	216	48
rect	218	47	219	48
rect	221	47	222	48
rect	244	47	245	48
rect	246	47	247	48
rect	250	47	251	48
rect	253	47	254	48
rect	256	47	257	48
rect	258	47	259	48
rect	261	47	262	48
rect	270	47	271	48
rect	273	47	274	48
rect	276	47	277	48
rect	278	47	279	48
rect	302	47	303	48
rect	305	47	306	48
rect	309	47	310	48
rect	14	48	15	49
rect	30	48	31	49
rect	47	48	48	49
rect	53	48	54	49
rect	56	48	57	49
rect	62	48	63	49
rect	71	48	72	49
rect	77	48	78	49
rect	108	48	109	49
rect	114	48	115	49
rect	146	48	147	49
rect	149	48	150	49
rect	152	48	153	49
rect	161	48	162	49
rect	176	48	177	49
rect	179	48	180	49
rect	182	48	183	49
rect	191	48	192	49
rect	194	48	195	49
rect	197	48	198	49
rect	200	48	201	49
rect	203	48	204	49
rect	209	48	210	49
rect	215	48	216	49
rect	218	48	219	49
rect	221	48	222	49
rect	244	48	245	49
rect	246	48	247	49
rect	253	48	254	49
rect	256	48	257	49
rect	258	48	259	49
rect	261	48	262	49
rect	270	48	271	49
rect	273	48	274	49
rect	276	48	277	49
rect	278	48	279	49
rect	302	48	303	49
rect	305	48	306	49
rect	309	48	310	49
rect	14	49	15	50
rect	30	49	31	50
rect	47	49	48	50
rect	53	49	54	50
rect	56	49	57	50
rect	62	49	63	50
rect	71	49	72	50
rect	77	49	78	50
rect	108	49	109	50
rect	114	49	115	50
rect	146	49	147	50
rect	149	49	150	50
rect	152	49	153	50
rect	161	49	162	50
rect	173	49	174	50
rect	176	49	177	50
rect	179	49	180	50
rect	182	49	183	50
rect	191	49	192	50
rect	194	49	195	50
rect	197	49	198	50
rect	200	49	201	50
rect	203	49	204	50
rect	209	49	210	50
rect	215	49	216	50
rect	218	49	219	50
rect	221	49	222	50
rect	227	49	228	50
rect	233	49	234	50
rect	244	49	245	50
rect	246	49	247	50
rect	253	49	254	50
rect	256	49	257	50
rect	258	49	259	50
rect	261	49	262	50
rect	270	49	271	50
rect	273	49	274	50
rect	276	49	277	50
rect	278	49	279	50
rect	300	49	301	50
rect	302	49	303	50
rect	305	49	306	50
rect	309	49	310	50
rect	14	50	15	51
rect	30	50	31	51
rect	47	50	48	51
rect	53	50	54	51
rect	56	50	57	51
rect	62	50	63	51
rect	71	50	72	51
rect	77	50	78	51
rect	108	50	109	51
rect	114	50	115	51
rect	146	50	147	51
rect	149	50	150	51
rect	161	50	162	51
rect	173	50	174	51
rect	176	50	177	51
rect	179	50	180	51
rect	191	50	192	51
rect	194	50	195	51
rect	197	50	198	51
rect	200	50	201	51
rect	203	50	204	51
rect	215	50	216	51
rect	218	50	219	51
rect	227	50	228	51
rect	233	50	234	51
rect	244	50	245	51
rect	246	50	247	51
rect	253	50	254	51
rect	256	50	257	51
rect	258	50	259	51
rect	261	50	262	51
rect	270	50	271	51
rect	273	50	274	51
rect	276	50	277	51
rect	278	50	279	51
rect	300	50	301	51
rect	302	50	303	51
rect	309	50	310	51
rect	14	51	15	52
rect	30	51	31	52
rect	47	51	48	52
rect	53	51	54	52
rect	56	51	57	52
rect	62	51	63	52
rect	71	51	72	52
rect	77	51	78	52
rect	108	51	109	52
rect	114	51	115	52
rect	119	51	120	52
rect	122	51	123	52
rect	146	51	147	52
rect	149	51	150	52
rect	161	51	162	52
rect	167	51	168	52
rect	170	51	171	52
rect	173	51	174	52
rect	176	51	177	52
rect	179	51	180	52
rect	191	51	192	52
rect	194	51	195	52
rect	197	51	198	52
rect	200	51	201	52
rect	203	51	204	52
rect	206	51	207	52
rect	215	51	216	52
rect	218	51	219	52
rect	227	51	228	52
rect	230	51	231	52
rect	233	51	234	52
rect	240	51	241	52
rect	244	51	245	52
rect	246	51	247	52
rect	253	51	254	52
rect	256	51	257	52
rect	258	51	259	52
rect	261	51	262	52
rect	270	51	271	52
rect	273	51	274	52
rect	276	51	277	52
rect	278	51	279	52
rect	288	51	289	52
rect	300	51	301	52
rect	302	51	303	52
rect	309	51	310	52
rect	330	51	331	52
rect	14	52	15	53
rect	30	52	31	53
rect	47	52	48	53
rect	53	52	54	53
rect	71	52	72	53
rect	108	52	109	53
rect	114	52	115	53
rect	119	52	120	53
rect	122	52	123	53
rect	146	52	147	53
rect	149	52	150	53
rect	161	52	162	53
rect	167	52	168	53
rect	170	52	171	53
rect	173	52	174	53
rect	176	52	177	53
rect	179	52	180	53
rect	191	52	192	53
rect	194	52	195	53
rect	197	52	198	53
rect	200	52	201	53
rect	203	52	204	53
rect	206	52	207	53
rect	215	52	216	53
rect	218	52	219	53
rect	227	52	228	53
rect	230	52	231	53
rect	233	52	234	53
rect	240	52	241	53
rect	244	52	245	53
rect	246	52	247	53
rect	253	52	254	53
rect	256	52	257	53
rect	258	52	259	53
rect	261	52	262	53
rect	270	52	271	53
rect	273	52	274	53
rect	276	52	277	53
rect	278	52	279	53
rect	288	52	289	53
rect	300	52	301	53
rect	309	52	310	53
rect	330	52	331	53
rect	14	53	15	54
rect	30	53	31	54
rect	47	53	48	54
rect	53	53	54	54
rect	71	53	72	54
rect	108	53	109	54
rect	114	53	115	54
rect	119	53	120	54
rect	122	53	123	54
rect	146	53	147	54
rect	149	53	150	54
rect	161	53	162	54
rect	167	53	168	54
rect	170	53	171	54
rect	173	53	174	54
rect	176	53	177	54
rect	179	53	180	54
rect	191	53	192	54
rect	194	53	195	54
rect	197	53	198	54
rect	200	53	201	54
rect	203	53	204	54
rect	206	53	207	54
rect	215	53	216	54
rect	218	53	219	54
rect	227	53	228	54
rect	230	53	231	54
rect	233	53	234	54
rect	240	53	241	54
rect	244	53	245	54
rect	246	53	247	54
rect	253	53	254	54
rect	256	53	257	54
rect	258	53	259	54
rect	261	53	262	54
rect	267	53	268	54
rect	270	53	271	54
rect	273	53	274	54
rect	276	53	277	54
rect	278	53	279	54
rect	288	53	289	54
rect	300	53	301	54
rect	309	53	310	54
rect	330	53	331	54
rect	339	53	340	54
rect	14	54	15	55
rect	30	54	31	55
rect	47	54	48	55
rect	119	54	120	55
rect	122	54	123	55
rect	146	54	147	55
rect	161	54	162	55
rect	167	54	168	55
rect	170	54	171	55
rect	173	54	174	55
rect	176	54	177	55
rect	197	54	198	55
rect	200	54	201	55
rect	203	54	204	55
rect	206	54	207	55
rect	215	54	216	55
rect	218	54	219	55
rect	227	54	228	55
rect	230	54	231	55
rect	233	54	234	55
rect	240	54	241	55
rect	244	54	245	55
rect	246	54	247	55
rect	253	54	254	55
rect	256	54	257	55
rect	258	54	259	55
rect	261	54	262	55
rect	267	54	268	55
rect	270	54	271	55
rect	273	54	274	55
rect	276	54	277	55
rect	278	54	279	55
rect	288	54	289	55
rect	300	54	301	55
rect	309	54	310	55
rect	330	54	331	55
rect	339	54	340	55
rect	14	55	15	56
rect	30	55	31	56
rect	47	55	48	56
rect	62	55	63	56
rect	80	55	81	56
rect	110	55	111	56
rect	119	55	120	56
rect	122	55	123	56
rect	128	55	129	56
rect	146	55	147	56
rect	158	55	159	56
rect	161	55	162	56
rect	164	55	165	56
rect	167	55	168	56
rect	170	55	171	56
rect	173	55	174	56
rect	176	55	177	56
rect	188	55	189	56
rect	197	55	198	56
rect	200	55	201	56
rect	203	55	204	56
rect	206	55	207	56
rect	215	55	216	56
rect	218	55	219	56
rect	227	55	228	56
rect	230	55	231	56
rect	233	55	234	56
rect	240	55	241	56
rect	244	55	245	56
rect	246	55	247	56
rect	253	55	254	56
rect	256	55	257	56
rect	258	55	259	56
rect	261	55	262	56
rect	267	55	268	56
rect	270	55	271	56
rect	273	55	274	56
rect	276	55	277	56
rect	278	55	279	56
rect	288	55	289	56
rect	300	55	301	56
rect	309	55	310	56
rect	330	55	331	56
rect	339	55	340	56
rect	357	55	358	56
rect	14	56	15	57
rect	30	56	31	57
rect	47	56	48	57
rect	62	56	63	57
rect	80	56	81	57
rect	110	56	111	57
rect	119	56	120	57
rect	122	56	123	57
rect	128	56	129	57
rect	146	56	147	57
rect	158	56	159	57
rect	161	56	162	57
rect	164	56	165	57
rect	167	56	168	57
rect	170	56	171	57
rect	173	56	174	57
rect	176	56	177	57
rect	188	56	189	57
rect	197	56	198	57
rect	200	56	201	57
rect	203	56	204	57
rect	206	56	207	57
rect	215	56	216	57
rect	218	56	219	57
rect	227	56	228	57
rect	230	56	231	57
rect	233	56	234	57
rect	240	56	241	57
rect	246	56	247	57
rect	258	56	259	57
rect	261	56	262	57
rect	267	56	268	57
rect	270	56	271	57
rect	273	56	274	57
rect	276	56	277	57
rect	288	56	289	57
rect	300	56	301	57
rect	309	56	310	57
rect	330	56	331	57
rect	339	56	340	57
rect	357	56	358	57
rect	14	57	15	58
rect	30	57	31	58
rect	34	57	35	58
rect	47	57	48	58
rect	62	57	63	58
rect	80	57	81	58
rect	110	57	111	58
rect	119	57	120	58
rect	122	57	123	58
rect	128	57	129	58
rect	146	57	147	58
rect	158	57	159	58
rect	161	57	162	58
rect	164	57	165	58
rect	167	57	168	58
rect	170	57	171	58
rect	173	57	174	58
rect	176	57	177	58
rect	179	57	180	58
rect	188	57	189	58
rect	191	57	192	58
rect	197	57	198	58
rect	200	57	201	58
rect	203	57	204	58
rect	206	57	207	58
rect	215	57	216	58
rect	218	57	219	58
rect	227	57	228	58
rect	230	57	231	58
rect	233	57	234	58
rect	240	57	241	58
rect	246	57	247	58
rect	249	57	250	58
rect	258	57	259	58
rect	261	57	262	58
rect	264	57	265	58
rect	267	57	268	58
rect	270	57	271	58
rect	273	57	274	58
rect	276	57	277	58
rect	279	57	280	58
rect	288	57	289	58
rect	297	57	298	58
rect	300	57	301	58
rect	306	57	307	58
rect	309	57	310	58
rect	330	57	331	58
rect	339	57	340	58
rect	357	57	358	58
rect	34	58	35	59
rect	62	58	63	59
rect	80	58	81	59
rect	110	58	111	59
rect	119	58	120	59
rect	122	58	123	59
rect	128	58	129	59
rect	158	58	159	59
rect	161	58	162	59
rect	164	58	165	59
rect	167	58	168	59
rect	170	58	171	59
rect	173	58	174	59
rect	176	58	177	59
rect	179	58	180	59
rect	188	58	189	59
rect	191	58	192	59
rect	197	58	198	59
rect	200	58	201	59
rect	203	58	204	59
rect	206	58	207	59
rect	215	58	216	59
rect	218	58	219	59
rect	227	58	228	59
rect	230	58	231	59
rect	233	58	234	59
rect	240	58	241	59
rect	246	58	247	59
rect	249	58	250	59
rect	258	58	259	59
rect	261	58	262	59
rect	264	58	265	59
rect	267	58	268	59
rect	270	58	271	59
rect	273	58	274	59
rect	276	58	277	59
rect	279	58	280	59
rect	288	58	289	59
rect	297	58	298	59
rect	300	58	301	59
rect	306	58	307	59
rect	309	58	310	59
rect	330	58	331	59
rect	339	58	340	59
rect	357	58	358	59
rect	21	59	22	60
rect	34	59	35	60
rect	37	59	38	60
rect	53	59	54	60
rect	62	59	63	60
rect	71	59	72	60
rect	80	59	81	60
rect	110	59	111	60
rect	119	59	120	60
rect	122	59	123	60
rect	128	59	129	60
rect	141	59	142	60
rect	158	59	159	60
rect	161	59	162	60
rect	164	59	165	60
rect	167	59	168	60
rect	170	59	171	60
rect	173	59	174	60
rect	176	59	177	60
rect	179	59	180	60
rect	188	59	189	60
rect	191	59	192	60
rect	197	59	198	60
rect	200	59	201	60
rect	203	59	204	60
rect	206	59	207	60
rect	215	59	216	60
rect	218	59	219	60
rect	227	59	228	60
rect	230	59	231	60
rect	233	59	234	60
rect	240	59	241	60
rect	246	59	247	60
rect	249	59	250	60
rect	258	59	259	60
rect	261	59	262	60
rect	264	59	265	60
rect	267	59	268	60
rect	270	59	271	60
rect	273	59	274	60
rect	276	59	277	60
rect	279	59	280	60
rect	288	59	289	60
rect	297	59	298	60
rect	300	59	301	60
rect	306	59	307	60
rect	309	59	310	60
rect	318	59	319	60
rect	321	59	322	60
rect	330	59	331	60
rect	333	59	334	60
rect	339	59	340	60
rect	348	59	349	60
rect	354	59	355	60
rect	357	59	358	60
rect	11	66	12	67
rect	21	66	22	67
rect	37	66	38	67
rect	50	66	51	67
rect	53	66	54	67
rect	62	66	63	67
rect	71	66	72	67
rect	77	66	78	67
rect	80	66	81	67
rect	110	66	111	67
rect	119	66	120	67
rect	128	66	129	67
rect	138	66	139	67
rect	148	66	149	67
rect	155	66	156	67
rect	158	66	159	67
rect	161	66	162	67
rect	164	66	165	67
rect	167	66	168	67
rect	170	66	171	67
rect	173	66	174	67
rect	176	66	177	67
rect	179	66	180	67
rect	188	66	189	67
rect	194	66	195	67
rect	197	66	198	67
rect	200	66	201	67
rect	203	66	204	67
rect	206	66	207	67
rect	209	66	210	67
rect	215	66	216	67
rect	218	66	219	67
rect	227	66	228	67
rect	230	66	231	67
rect	246	66	247	67
rect	249	66	250	67
rect	255	66	256	67
rect	258	66	259	67
rect	261	66	262	67
rect	264	66	265	67
rect	267	66	268	67
rect	276	66	277	67
rect	279	66	280	67
rect	288	66	289	67
rect	294	66	295	67
rect	297	66	298	67
rect	300	66	301	67
rect	309	66	310	67
rect	318	66	319	67
rect	321	66	322	67
rect	330	66	331	67
rect	339	66	340	67
rect	348	66	349	67
rect	357	66	358	67
rect	11	67	12	68
rect	21	67	22	68
rect	37	67	38	68
rect	50	67	51	68
rect	53	67	54	68
rect	62	67	63	68
rect	71	67	72	68
rect	77	67	78	68
rect	80	67	81	68
rect	110	67	111	68
rect	119	67	120	68
rect	128	67	129	68
rect	138	67	139	68
rect	148	67	149	68
rect	155	67	156	68
rect	158	67	159	68
rect	161	67	162	68
rect	164	67	165	68
rect	167	67	168	68
rect	170	67	171	68
rect	173	67	174	68
rect	176	67	177	68
rect	179	67	180	68
rect	188	67	189	68
rect	194	67	195	68
rect	197	67	198	68
rect	200	67	201	68
rect	203	67	204	68
rect	206	67	207	68
rect	209	67	210	68
rect	215	67	216	68
rect	218	67	219	68
rect	227	67	228	68
rect	230	67	231	68
rect	246	67	247	68
rect	249	67	250	68
rect	255	67	256	68
rect	258	67	259	68
rect	261	67	262	68
rect	264	67	265	68
rect	267	67	268	68
rect	276	67	277	68
rect	279	67	280	68
rect	288	67	289	68
rect	294	67	295	68
rect	297	67	298	68
rect	300	67	301	68
rect	309	67	310	68
rect	318	67	319	68
rect	321	67	322	68
rect	330	67	331	68
rect	339	67	340	68
rect	348	67	349	68
rect	11	68	12	69
rect	21	68	22	69
rect	37	68	38	69
rect	50	68	51	69
rect	53	68	54	69
rect	62	68	63	69
rect	71	68	72	69
rect	77	68	78	69
rect	80	68	81	69
rect	110	68	111	69
rect	119	68	120	69
rect	128	68	129	69
rect	138	68	139	69
rect	148	68	149	69
rect	155	68	156	69
rect	158	68	159	69
rect	161	68	162	69
rect	164	68	165	69
rect	167	68	168	69
rect	170	68	171	69
rect	173	68	174	69
rect	176	68	177	69
rect	179	68	180	69
rect	188	68	189	69
rect	194	68	195	69
rect	197	68	198	69
rect	200	68	201	69
rect	203	68	204	69
rect	206	68	207	69
rect	209	68	210	69
rect	215	68	216	69
rect	218	68	219	69
rect	227	68	228	69
rect	230	68	231	69
rect	246	68	247	69
rect	249	68	250	69
rect	255	68	256	69
rect	258	68	259	69
rect	261	68	262	69
rect	264	68	265	69
rect	267	68	268	69
rect	276	68	277	69
rect	279	68	280	69
rect	288	68	289	69
rect	294	68	295	69
rect	297	68	298	69
rect	300	68	301	69
rect	309	68	310	69
rect	318	68	319	69
rect	321	68	322	69
rect	330	68	331	69
rect	339	68	340	69
rect	348	68	349	69
rect	396	68	397	69
rect	11	69	12	70
rect	21	69	22	70
rect	37	69	38	70
rect	50	69	51	70
rect	53	69	54	70
rect	62	69	63	70
rect	71	69	72	70
rect	77	69	78	70
rect	80	69	81	70
rect	110	69	111	70
rect	119	69	120	70
rect	128	69	129	70
rect	138	69	139	70
rect	148	69	149	70
rect	155	69	156	70
rect	158	69	159	70
rect	161	69	162	70
rect	164	69	165	70
rect	167	69	168	70
rect	170	69	171	70
rect	173	69	174	70
rect	176	69	177	70
rect	179	69	180	70
rect	188	69	189	70
rect	194	69	195	70
rect	197	69	198	70
rect	200	69	201	70
rect	203	69	204	70
rect	206	69	207	70
rect	209	69	210	70
rect	215	69	216	70
rect	218	69	219	70
rect	227	69	228	70
rect	230	69	231	70
rect	246	69	247	70
rect	249	69	250	70
rect	255	69	256	70
rect	258	69	259	70
rect	261	69	262	70
rect	264	69	265	70
rect	267	69	268	70
rect	276	69	277	70
rect	279	69	280	70
rect	288	69	289	70
rect	294	69	295	70
rect	297	69	298	70
rect	300	69	301	70
rect	309	69	310	70
rect	318	69	319	70
rect	321	69	322	70
rect	330	69	331	70
rect	348	69	349	70
rect	396	69	397	70
rect	11	70	12	71
rect	21	70	22	71
rect	37	70	38	71
rect	50	70	51	71
rect	53	70	54	71
rect	62	70	63	71
rect	71	70	72	71
rect	77	70	78	71
rect	80	70	81	71
rect	110	70	111	71
rect	119	70	120	71
rect	128	70	129	71
rect	138	70	139	71
rect	148	70	149	71
rect	155	70	156	71
rect	158	70	159	71
rect	161	70	162	71
rect	164	70	165	71
rect	167	70	168	71
rect	170	70	171	71
rect	173	70	174	71
rect	176	70	177	71
rect	179	70	180	71
rect	188	70	189	71
rect	194	70	195	71
rect	197	70	198	71
rect	200	70	201	71
rect	203	70	204	71
rect	206	70	207	71
rect	209	70	210	71
rect	215	70	216	71
rect	218	70	219	71
rect	227	70	228	71
rect	230	70	231	71
rect	246	70	247	71
rect	249	70	250	71
rect	255	70	256	71
rect	258	70	259	71
rect	261	70	262	71
rect	264	70	265	71
rect	267	70	268	71
rect	276	70	277	71
rect	279	70	280	71
rect	288	70	289	71
rect	294	70	295	71
rect	297	70	298	71
rect	300	70	301	71
rect	309	70	310	71
rect	318	70	319	71
rect	321	70	322	71
rect	330	70	331	71
rect	348	70	349	71
rect	357	70	358	71
rect	396	70	397	71
rect	11	71	12	72
rect	21	71	22	72
rect	37	71	38	72
rect	50	71	51	72
rect	53	71	54	72
rect	62	71	63	72
rect	71	71	72	72
rect	77	71	78	72
rect	80	71	81	72
rect	110	71	111	72
rect	119	71	120	72
rect	128	71	129	72
rect	138	71	139	72
rect	148	71	149	72
rect	155	71	156	72
rect	158	71	159	72
rect	161	71	162	72
rect	164	71	165	72
rect	167	71	168	72
rect	170	71	171	72
rect	173	71	174	72
rect	176	71	177	72
rect	179	71	180	72
rect	188	71	189	72
rect	194	71	195	72
rect	197	71	198	72
rect	200	71	201	72
rect	203	71	204	72
rect	206	71	207	72
rect	209	71	210	72
rect	215	71	216	72
rect	218	71	219	72
rect	227	71	228	72
rect	230	71	231	72
rect	246	71	247	72
rect	249	71	250	72
rect	255	71	256	72
rect	258	71	259	72
rect	261	71	262	72
rect	264	71	265	72
rect	267	71	268	72
rect	276	71	277	72
rect	279	71	280	72
rect	288	71	289	72
rect	294	71	295	72
rect	297	71	298	72
rect	300	71	301	72
rect	309	71	310	72
rect	318	71	319	72
rect	321	71	322	72
rect	348	71	349	72
rect	357	71	358	72
rect	396	71	397	72
rect	11	72	12	73
rect	21	72	22	73
rect	37	72	38	73
rect	50	72	51	73
rect	53	72	54	73
rect	62	72	63	73
rect	71	72	72	73
rect	77	72	78	73
rect	80	72	81	73
rect	110	72	111	73
rect	119	72	120	73
rect	128	72	129	73
rect	138	72	139	73
rect	148	72	149	73
rect	155	72	156	73
rect	158	72	159	73
rect	161	72	162	73
rect	164	72	165	73
rect	167	72	168	73
rect	170	72	171	73
rect	173	72	174	73
rect	176	72	177	73
rect	179	72	180	73
rect	188	72	189	73
rect	194	72	195	73
rect	197	72	198	73
rect	200	72	201	73
rect	203	72	204	73
rect	206	72	207	73
rect	209	72	210	73
rect	215	72	216	73
rect	218	72	219	73
rect	227	72	228	73
rect	230	72	231	73
rect	246	72	247	73
rect	249	72	250	73
rect	255	72	256	73
rect	258	72	259	73
rect	261	72	262	73
rect	264	72	265	73
rect	267	72	268	73
rect	276	72	277	73
rect	279	72	280	73
rect	288	72	289	73
rect	294	72	295	73
rect	297	72	298	73
rect	300	72	301	73
rect	309	72	310	73
rect	318	72	319	73
rect	321	72	322	73
rect	339	72	340	73
rect	348	72	349	73
rect	357	72	358	73
rect	396	72	397	73
rect	11	73	12	74
rect	21	73	22	74
rect	37	73	38	74
rect	50	73	51	74
rect	53	73	54	74
rect	62	73	63	74
rect	71	73	72	74
rect	77	73	78	74
rect	80	73	81	74
rect	110	73	111	74
rect	119	73	120	74
rect	128	73	129	74
rect	138	73	139	74
rect	148	73	149	74
rect	155	73	156	74
rect	158	73	159	74
rect	161	73	162	74
rect	164	73	165	74
rect	167	73	168	74
rect	170	73	171	74
rect	173	73	174	74
rect	176	73	177	74
rect	179	73	180	74
rect	188	73	189	74
rect	194	73	195	74
rect	197	73	198	74
rect	200	73	201	74
rect	203	73	204	74
rect	206	73	207	74
rect	209	73	210	74
rect	215	73	216	74
rect	218	73	219	74
rect	227	73	228	74
rect	230	73	231	74
rect	246	73	247	74
rect	249	73	250	74
rect	255	73	256	74
rect	258	73	259	74
rect	261	73	262	74
rect	264	73	265	74
rect	267	73	268	74
rect	276	73	277	74
rect	279	73	280	74
rect	288	73	289	74
rect	297	73	298	74
rect	300	73	301	74
rect	309	73	310	74
rect	318	73	319	74
rect	321	73	322	74
rect	339	73	340	74
rect	348	73	349	74
rect	357	73	358	74
rect	396	73	397	74
rect	11	74	12	75
rect	21	74	22	75
rect	37	74	38	75
rect	50	74	51	75
rect	53	74	54	75
rect	62	74	63	75
rect	71	74	72	75
rect	77	74	78	75
rect	80	74	81	75
rect	110	74	111	75
rect	119	74	120	75
rect	128	74	129	75
rect	138	74	139	75
rect	148	74	149	75
rect	155	74	156	75
rect	158	74	159	75
rect	161	74	162	75
rect	164	74	165	75
rect	167	74	168	75
rect	170	74	171	75
rect	173	74	174	75
rect	176	74	177	75
rect	179	74	180	75
rect	188	74	189	75
rect	194	74	195	75
rect	197	74	198	75
rect	200	74	201	75
rect	203	74	204	75
rect	206	74	207	75
rect	209	74	210	75
rect	215	74	216	75
rect	218	74	219	75
rect	227	74	228	75
rect	230	74	231	75
rect	246	74	247	75
rect	249	74	250	75
rect	255	74	256	75
rect	258	74	259	75
rect	261	74	262	75
rect	264	74	265	75
rect	267	74	268	75
rect	276	74	277	75
rect	279	74	280	75
rect	288	74	289	75
rect	297	74	298	75
rect	300	74	301	75
rect	309	74	310	75
rect	318	74	319	75
rect	321	74	322	75
rect	330	74	331	75
rect	339	74	340	75
rect	348	74	349	75
rect	357	74	358	75
rect	396	74	397	75
rect	11	75	12	76
rect	21	75	22	76
rect	37	75	38	76
rect	50	75	51	76
rect	53	75	54	76
rect	62	75	63	76
rect	71	75	72	76
rect	77	75	78	76
rect	80	75	81	76
rect	110	75	111	76
rect	119	75	120	76
rect	128	75	129	76
rect	138	75	139	76
rect	148	75	149	76
rect	155	75	156	76
rect	158	75	159	76
rect	161	75	162	76
rect	164	75	165	76
rect	167	75	168	76
rect	170	75	171	76
rect	173	75	174	76
rect	176	75	177	76
rect	179	75	180	76
rect	188	75	189	76
rect	194	75	195	76
rect	197	75	198	76
rect	200	75	201	76
rect	203	75	204	76
rect	206	75	207	76
rect	209	75	210	76
rect	215	75	216	76
rect	218	75	219	76
rect	227	75	228	76
rect	230	75	231	76
rect	246	75	247	76
rect	249	75	250	76
rect	255	75	256	76
rect	258	75	259	76
rect	261	75	262	76
rect	264	75	265	76
rect	267	75	268	76
rect	276	75	277	76
rect	279	75	280	76
rect	297	75	298	76
rect	300	75	301	76
rect	309	75	310	76
rect	318	75	319	76
rect	321	75	322	76
rect	330	75	331	76
rect	339	75	340	76
rect	348	75	349	76
rect	357	75	358	76
rect	396	75	397	76
rect	11	76	12	77
rect	21	76	22	77
rect	37	76	38	77
rect	50	76	51	77
rect	53	76	54	77
rect	62	76	63	77
rect	71	76	72	77
rect	77	76	78	77
rect	80	76	81	77
rect	110	76	111	77
rect	119	76	120	77
rect	128	76	129	77
rect	138	76	139	77
rect	148	76	149	77
rect	155	76	156	77
rect	158	76	159	77
rect	161	76	162	77
rect	164	76	165	77
rect	167	76	168	77
rect	170	76	171	77
rect	173	76	174	77
rect	176	76	177	77
rect	179	76	180	77
rect	188	76	189	77
rect	194	76	195	77
rect	197	76	198	77
rect	200	76	201	77
rect	203	76	204	77
rect	206	76	207	77
rect	209	76	210	77
rect	215	76	216	77
rect	218	76	219	77
rect	227	76	228	77
rect	230	76	231	77
rect	246	76	247	77
rect	249	76	250	77
rect	255	76	256	77
rect	258	76	259	77
rect	261	76	262	77
rect	264	76	265	77
rect	267	76	268	77
rect	276	76	277	77
rect	279	76	280	77
rect	297	76	298	77
rect	300	76	301	77
rect	309	76	310	77
rect	315	76	316	77
rect	318	76	319	77
rect	321	76	322	77
rect	330	76	331	77
rect	339	76	340	77
rect	348	76	349	77
rect	357	76	358	77
rect	396	76	397	77
rect	11	77	12	78
rect	21	77	22	78
rect	37	77	38	78
rect	50	77	51	78
rect	53	77	54	78
rect	62	77	63	78
rect	71	77	72	78
rect	77	77	78	78
rect	80	77	81	78
rect	110	77	111	78
rect	119	77	120	78
rect	128	77	129	78
rect	138	77	139	78
rect	148	77	149	78
rect	155	77	156	78
rect	158	77	159	78
rect	161	77	162	78
rect	164	77	165	78
rect	167	77	168	78
rect	170	77	171	78
rect	173	77	174	78
rect	176	77	177	78
rect	179	77	180	78
rect	188	77	189	78
rect	194	77	195	78
rect	197	77	198	78
rect	203	77	204	78
rect	206	77	207	78
rect	209	77	210	78
rect	215	77	216	78
rect	218	77	219	78
rect	227	77	228	78
rect	230	77	231	78
rect	246	77	247	78
rect	249	77	250	78
rect	255	77	256	78
rect	258	77	259	78
rect	261	77	262	78
rect	264	77	265	78
rect	267	77	268	78
rect	276	77	277	78
rect	279	77	280	78
rect	297	77	298	78
rect	300	77	301	78
rect	309	77	310	78
rect	315	77	316	78
rect	318	77	319	78
rect	321	77	322	78
rect	330	77	331	78
rect	339	77	340	78
rect	348	77	349	78
rect	357	77	358	78
rect	396	77	397	78
rect	11	78	12	79
rect	21	78	22	79
rect	37	78	38	79
rect	50	78	51	79
rect	53	78	54	79
rect	62	78	63	79
rect	71	78	72	79
rect	77	78	78	79
rect	80	78	81	79
rect	110	78	111	79
rect	119	78	120	79
rect	128	78	129	79
rect	138	78	139	79
rect	148	78	149	79
rect	155	78	156	79
rect	158	78	159	79
rect	161	78	162	79
rect	164	78	165	79
rect	167	78	168	79
rect	170	78	171	79
rect	173	78	174	79
rect	176	78	177	79
rect	179	78	180	79
rect	188	78	189	79
rect	194	78	195	79
rect	197	78	198	79
rect	203	78	204	79
rect	206	78	207	79
rect	209	78	210	79
rect	215	78	216	79
rect	218	78	219	79
rect	227	78	228	79
rect	230	78	231	79
rect	246	78	247	79
rect	249	78	250	79
rect	255	78	256	79
rect	258	78	259	79
rect	261	78	262	79
rect	264	78	265	79
rect	267	78	268	79
rect	276	78	277	79
rect	279	78	280	79
rect	297	78	298	79
rect	300	78	301	79
rect	309	78	310	79
rect	315	78	316	79
rect	318	78	319	79
rect	321	78	322	79
rect	324	78	325	79
rect	330	78	331	79
rect	339	78	340	79
rect	348	78	349	79
rect	357	78	358	79
rect	396	78	397	79
rect	11	79	12	80
rect	21	79	22	80
rect	37	79	38	80
rect	50	79	51	80
rect	53	79	54	80
rect	62	79	63	80
rect	71	79	72	80
rect	77	79	78	80
rect	80	79	81	80
rect	110	79	111	80
rect	119	79	120	80
rect	128	79	129	80
rect	138	79	139	80
rect	148	79	149	80
rect	155	79	156	80
rect	158	79	159	80
rect	161	79	162	80
rect	164	79	165	80
rect	170	79	171	80
rect	173	79	174	80
rect	176	79	177	80
rect	179	79	180	80
rect	188	79	189	80
rect	194	79	195	80
rect	197	79	198	80
rect	203	79	204	80
rect	206	79	207	80
rect	209	79	210	80
rect	215	79	216	80
rect	218	79	219	80
rect	227	79	228	80
rect	230	79	231	80
rect	246	79	247	80
rect	255	79	256	80
rect	258	79	259	80
rect	261	79	262	80
rect	267	79	268	80
rect	276	79	277	80
rect	279	79	280	80
rect	297	79	298	80
rect	300	79	301	80
rect	309	79	310	80
rect	315	79	316	80
rect	318	79	319	80
rect	321	79	322	80
rect	324	79	325	80
rect	330	79	331	80
rect	339	79	340	80
rect	348	79	349	80
rect	357	79	358	80
rect	396	79	397	80
rect	11	80	12	81
rect	21	80	22	81
rect	37	80	38	81
rect	50	80	51	81
rect	53	80	54	81
rect	62	80	63	81
rect	71	80	72	81
rect	77	80	78	81
rect	80	80	81	81
rect	110	80	111	81
rect	119	80	120	81
rect	128	80	129	81
rect	138	80	139	81
rect	148	80	149	81
rect	155	80	156	81
rect	158	80	159	81
rect	161	80	162	81
rect	164	80	165	81
rect	170	80	171	81
rect	173	80	174	81
rect	176	80	177	81
rect	179	80	180	81
rect	188	80	189	81
rect	194	80	195	81
rect	197	80	198	81
rect	200	80	201	81
rect	203	80	204	81
rect	206	80	207	81
rect	209	80	210	81
rect	215	80	216	81
rect	218	80	219	81
rect	227	80	228	81
rect	230	80	231	81
rect	246	80	247	81
rect	252	80	253	81
rect	255	80	256	81
rect	258	80	259	81
rect	261	80	262	81
rect	267	80	268	81
rect	276	80	277	81
rect	279	80	280	81
rect	294	80	295	81
rect	297	80	298	81
rect	300	80	301	81
rect	309	80	310	81
rect	315	80	316	81
rect	318	80	319	81
rect	321	80	322	81
rect	324	80	325	81
rect	330	80	331	81
rect	339	80	340	81
rect	348	80	349	81
rect	357	80	358	81
rect	396	80	397	81
rect	11	81	12	82
rect	21	81	22	82
rect	37	81	38	82
rect	50	81	51	82
rect	53	81	54	82
rect	62	81	63	82
rect	71	81	72	82
rect	77	81	78	82
rect	80	81	81	82
rect	110	81	111	82
rect	119	81	120	82
rect	128	81	129	82
rect	138	81	139	82
rect	155	81	156	82
rect	158	81	159	82
rect	161	81	162	82
rect	164	81	165	82
rect	170	81	171	82
rect	173	81	174	82
rect	176	81	177	82
rect	179	81	180	82
rect	194	81	195	82
rect	197	81	198	82
rect	200	81	201	82
rect	203	81	204	82
rect	206	81	207	82
rect	209	81	210	82
rect	215	81	216	82
rect	218	81	219	82
rect	230	81	231	82
rect	246	81	247	82
rect	252	81	253	82
rect	255	81	256	82
rect	258	81	259	82
rect	267	81	268	82
rect	276	81	277	82
rect	279	81	280	82
rect	294	81	295	82
rect	297	81	298	82
rect	300	81	301	82
rect	309	81	310	82
rect	315	81	316	82
rect	318	81	319	82
rect	321	81	322	82
rect	324	81	325	82
rect	330	81	331	82
rect	339	81	340	82
rect	348	81	349	82
rect	357	81	358	82
rect	396	81	397	82
rect	11	82	12	83
rect	21	82	22	83
rect	37	82	38	83
rect	50	82	51	83
rect	53	82	54	83
rect	62	82	63	83
rect	71	82	72	83
rect	77	82	78	83
rect	80	82	81	83
rect	110	82	111	83
rect	119	82	120	83
rect	128	82	129	83
rect	138	82	139	83
rect	155	82	156	83
rect	158	82	159	83
rect	161	82	162	83
rect	164	82	165	83
rect	170	82	171	83
rect	173	82	174	83
rect	176	82	177	83
rect	179	82	180	83
rect	194	82	195	83
rect	197	82	198	83
rect	200	82	201	83
rect	203	82	204	83
rect	206	82	207	83
rect	209	82	210	83
rect	215	82	216	83
rect	218	82	219	83
rect	230	82	231	83
rect	246	82	247	83
rect	249	82	250	83
rect	252	82	253	83
rect	255	82	256	83
rect	258	82	259	83
rect	267	82	268	83
rect	276	82	277	83
rect	279	82	280	83
rect	291	82	292	83
rect	294	82	295	83
rect	297	82	298	83
rect	300	82	301	83
rect	309	82	310	83
rect	315	82	316	83
rect	318	82	319	83
rect	321	82	322	83
rect	324	82	325	83
rect	330	82	331	83
rect	339	82	340	83
rect	348	82	349	83
rect	357	82	358	83
rect	396	82	397	83
rect	11	83	12	84
rect	21	83	22	84
rect	37	83	38	84
rect	50	83	51	84
rect	53	83	54	84
rect	62	83	63	84
rect	71	83	72	84
rect	77	83	78	84
rect	80	83	81	84
rect	110	83	111	84
rect	119	83	120	84
rect	128	83	129	84
rect	138	83	139	84
rect	155	83	156	84
rect	158	83	159	84
rect	161	83	162	84
rect	170	83	171	84
rect	173	83	174	84
rect	176	83	177	84
rect	179	83	180	84
rect	194	83	195	84
rect	197	83	198	84
rect	200	83	201	84
rect	203	83	204	84
rect	206	83	207	84
rect	209	83	210	84
rect	215	83	216	84
rect	230	83	231	84
rect	246	83	247	84
rect	249	83	250	84
rect	252	83	253	84
rect	255	83	256	84
rect	267	83	268	84
rect	276	83	277	84
rect	279	83	280	84
rect	291	83	292	84
rect	294	83	295	84
rect	297	83	298	84
rect	300	83	301	84
rect	309	83	310	84
rect	315	83	316	84
rect	318	83	319	84
rect	321	83	322	84
rect	324	83	325	84
rect	330	83	331	84
rect	339	83	340	84
rect	348	83	349	84
rect	357	83	358	84
rect	396	83	397	84
rect	11	84	12	85
rect	21	84	22	85
rect	37	84	38	85
rect	50	84	51	85
rect	53	84	54	85
rect	62	84	63	85
rect	71	84	72	85
rect	77	84	78	85
rect	80	84	81	85
rect	110	84	111	85
rect	119	84	120	85
rect	128	84	129	85
rect	138	84	139	85
rect	155	84	156	85
rect	158	84	159	85
rect	161	84	162	85
rect	170	84	171	85
rect	173	84	174	85
rect	176	84	177	85
rect	179	84	180	85
rect	188	84	189	85
rect	194	84	195	85
rect	197	84	198	85
rect	200	84	201	85
rect	203	84	204	85
rect	206	84	207	85
rect	209	84	210	85
rect	215	84	216	85
rect	228	84	229	85
rect	230	84	231	85
rect	246	84	247	85
rect	249	84	250	85
rect	252	84	253	85
rect	255	84	256	85
rect	267	84	268	85
rect	276	84	277	85
rect	279	84	280	85
rect	288	84	289	85
rect	291	84	292	85
rect	294	84	295	85
rect	297	84	298	85
rect	300	84	301	85
rect	309	84	310	85
rect	315	84	316	85
rect	318	84	319	85
rect	321	84	322	85
rect	324	84	325	85
rect	330	84	331	85
rect	339	84	340	85
rect	348	84	349	85
rect	357	84	358	85
rect	396	84	397	85
rect	11	85	12	86
rect	21	85	22	86
rect	37	85	38	86
rect	50	85	51	86
rect	53	85	54	86
rect	62	85	63	86
rect	71	85	72	86
rect	77	85	78	86
rect	80	85	81	86
rect	110	85	111	86
rect	119	85	120	86
rect	128	85	129	86
rect	138	85	139	86
rect	155	85	156	86
rect	158	85	159	86
rect	173	85	174	86
rect	176	85	177	86
rect	179	85	180	86
rect	188	85	189	86
rect	197	85	198	86
rect	200	85	201	86
rect	203	85	204	86
rect	206	85	207	86
rect	209	85	210	86
rect	215	85	216	86
rect	228	85	229	86
rect	230	85	231	86
rect	246	85	247	86
rect	249	85	250	86
rect	252	85	253	86
rect	255	85	256	86
rect	267	85	268	86
rect	276	85	277	86
rect	279	85	280	86
rect	288	85	289	86
rect	291	85	292	86
rect	294	85	295	86
rect	300	85	301	86
rect	309	85	310	86
rect	315	85	316	86
rect	318	85	319	86
rect	321	85	322	86
rect	324	85	325	86
rect	330	85	331	86
rect	339	85	340	86
rect	357	85	358	86
rect	396	85	397	86
rect	11	86	12	87
rect	21	86	22	87
rect	37	86	38	87
rect	50	86	51	87
rect	53	86	54	87
rect	62	86	63	87
rect	71	86	72	87
rect	77	86	78	87
rect	80	86	81	87
rect	110	86	111	87
rect	119	86	120	87
rect	128	86	129	87
rect	138	86	139	87
rect	155	86	156	87
rect	158	86	159	87
rect	164	86	165	87
rect	167	86	168	87
rect	173	86	174	87
rect	176	86	177	87
rect	179	86	180	87
rect	188	86	189	87
rect	197	86	198	87
rect	200	86	201	87
rect	203	86	204	87
rect	206	86	207	87
rect	209	86	210	87
rect	215	86	216	87
rect	228	86	229	87
rect	230	86	231	87
rect	246	86	247	87
rect	249	86	250	87
rect	252	86	253	87
rect	255	86	256	87
rect	267	86	268	87
rect	270	86	271	87
rect	276	86	277	87
rect	279	86	280	87
rect	288	86	289	87
rect	291	86	292	87
rect	294	86	295	87
rect	300	86	301	87
rect	309	86	310	87
rect	315	86	316	87
rect	318	86	319	87
rect	321	86	322	87
rect	324	86	325	87
rect	330	86	331	87
rect	333	86	334	87
rect	339	86	340	87
rect	357	86	358	87
rect	369	86	370	87
rect	396	86	397	87
rect	11	87	12	88
rect	21	87	22	88
rect	37	87	38	88
rect	50	87	51	88
rect	62	87	63	88
rect	80	87	81	88
rect	110	87	111	88
rect	119	87	120	88
rect	128	87	129	88
rect	155	87	156	88
rect	164	87	165	88
rect	167	87	168	88
rect	173	87	174	88
rect	176	87	177	88
rect	179	87	180	88
rect	188	87	189	88
rect	197	87	198	88
rect	200	87	201	88
rect	206	87	207	88
rect	209	87	210	88
rect	215	87	216	88
rect	228	87	229	88
rect	230	87	231	88
rect	246	87	247	88
rect	249	87	250	88
rect	252	87	253	88
rect	267	87	268	88
rect	270	87	271	88
rect	276	87	277	88
rect	279	87	280	88
rect	288	87	289	88
rect	291	87	292	88
rect	294	87	295	88
rect	300	87	301	88
rect	309	87	310	88
rect	315	87	316	88
rect	321	87	322	88
rect	324	87	325	88
rect	330	87	331	88
rect	333	87	334	88
rect	339	87	340	88
rect	357	87	358	88
rect	369	87	370	88
rect	396	87	397	88
rect	11	88	12	89
rect	21	88	22	89
rect	37	88	38	89
rect	50	88	51	89
rect	59	88	60	89
rect	62	88	63	89
rect	68	88	69	89
rect	80	88	81	89
rect	110	88	111	89
rect	112	88	113	89
rect	119	88	120	89
rect	128	88	129	89
rect	148	88	149	89
rect	155	88	156	89
rect	164	88	165	89
rect	167	88	168	89
rect	173	88	174	89
rect	176	88	177	89
rect	179	88	180	89
rect	188	88	189	89
rect	194	88	195	89
rect	197	88	198	89
rect	200	88	201	89
rect	206	88	207	89
rect	209	88	210	89
rect	215	88	216	89
rect	225	88	226	89
rect	228	88	229	89
rect	230	88	231	89
rect	246	88	247	89
rect	249	88	250	89
rect	252	88	253	89
rect	267	88	268	89
rect	270	88	271	89
rect	276	88	277	89
rect	279	88	280	89
rect	288	88	289	89
rect	291	88	292	89
rect	294	88	295	89
rect	300	88	301	89
rect	306	88	307	89
rect	309	88	310	89
rect	315	88	316	89
rect	321	88	322	89
rect	324	88	325	89
rect	330	88	331	89
rect	333	88	334	89
rect	339	88	340	89
rect	348	88	349	89
rect	357	88	358	89
rect	369	88	370	89
rect	396	88	397	89
rect	11	89	12	90
rect	21	89	22	90
rect	59	89	60	90
rect	62	89	63	90
rect	68	89	69	90
rect	80	89	81	90
rect	110	89	111	90
rect	112	89	113	90
rect	119	89	120	90
rect	128	89	129	90
rect	148	89	149	90
rect	155	89	156	90
rect	164	89	165	90
rect	167	89	168	90
rect	173	89	174	90
rect	176	89	177	90
rect	179	89	180	90
rect	188	89	189	90
rect	194	89	195	90
rect	197	89	198	90
rect	200	89	201	90
rect	206	89	207	90
rect	209	89	210	90
rect	225	89	226	90
rect	228	89	229	90
rect	246	89	247	90
rect	249	89	250	90
rect	252	89	253	90
rect	267	89	268	90
rect	270	89	271	90
rect	279	89	280	90
rect	288	89	289	90
rect	291	89	292	90
rect	294	89	295	90
rect	300	89	301	90
rect	306	89	307	90
rect	309	89	310	90
rect	315	89	316	90
rect	324	89	325	90
rect	330	89	331	90
rect	333	89	334	90
rect	339	89	340	90
rect	348	89	349	90
rect	357	89	358	90
rect	369	89	370	90
rect	396	89	397	90
rect	11	90	12	91
rect	21	90	22	91
rect	40	90	41	91
rect	59	90	60	91
rect	62	90	63	91
rect	68	90	69	91
rect	80	90	81	91
rect	110	90	111	91
rect	112	90	113	91
rect	119	90	120	91
rect	128	90	129	91
rect	148	90	149	91
rect	155	90	156	91
rect	164	90	165	91
rect	167	90	168	91
rect	173	90	174	91
rect	176	90	177	91
rect	179	90	180	91
rect	188	90	189	91
rect	194	90	195	91
rect	197	90	198	91
rect	200	90	201	91
rect	203	90	204	91
rect	206	90	207	91
rect	209	90	210	91
rect	219	90	220	91
rect	225	90	226	91
rect	228	90	229	91
rect	246	90	247	91
rect	249	90	250	91
rect	252	90	253	91
rect	264	90	265	91
rect	267	90	268	91
rect	270	90	271	91
rect	279	90	280	91
rect	288	90	289	91
rect	291	90	292	91
rect	294	90	295	91
rect	297	90	298	91
rect	300	90	301	91
rect	306	90	307	91
rect	309	90	310	91
rect	315	90	316	91
rect	318	90	319	91
rect	324	90	325	91
rect	330	90	331	91
rect	333	90	334	91
rect	339	90	340	91
rect	348	90	349	91
rect	357	90	358	91
rect	369	90	370	91
rect	396	90	397	91
rect	11	91	12	92
rect	21	91	22	92
rect	40	91	41	92
rect	59	91	60	92
rect	68	91	69	92
rect	110	91	111	92
rect	112	91	113	92
rect	128	91	129	92
rect	148	91	149	92
rect	155	91	156	92
rect	164	91	165	92
rect	167	91	168	92
rect	173	91	174	92
rect	176	91	177	92
rect	179	91	180	92
rect	188	91	189	92
rect	194	91	195	92
rect	197	91	198	92
rect	200	91	201	92
rect	203	91	204	92
rect	206	91	207	92
rect	209	91	210	92
rect	219	91	220	92
rect	225	91	226	92
rect	228	91	229	92
rect	246	91	247	92
rect	249	91	250	92
rect	252	91	253	92
rect	264	91	265	92
rect	267	91	268	92
rect	270	91	271	92
rect	279	91	280	92
rect	288	91	289	92
rect	291	91	292	92
rect	294	91	295	92
rect	297	91	298	92
rect	300	91	301	92
rect	306	91	307	92
rect	309	91	310	92
rect	315	91	316	92
rect	318	91	319	92
rect	324	91	325	92
rect	330	91	331	92
rect	333	91	334	92
rect	339	91	340	92
rect	348	91	349	92
rect	357	91	358	92
rect	369	91	370	92
rect	396	91	397	92
rect	11	92	12	93
rect	21	92	22	93
rect	34	92	35	93
rect	37	92	38	93
rect	40	92	41	93
rect	50	92	51	93
rect	56	92	57	93
rect	59	92	60	93
rect	68	92	69	93
rect	77	92	78	93
rect	86	92	87	93
rect	110	92	111	93
rect	112	92	113	93
rect	128	92	129	93
rect	130	92	131	93
rect	136	92	137	93
rect	139	92	140	93
rect	142	92	143	93
rect	148	92	149	93
rect	155	92	156	93
rect	164	92	165	93
rect	167	92	168	93
rect	173	92	174	93
rect	176	92	177	93
rect	179	92	180	93
rect	188	92	189	93
rect	194	92	195	93
rect	197	92	198	93
rect	200	92	201	93
rect	203	92	204	93
rect	206	92	207	93
rect	209	92	210	93
rect	219	92	220	93
rect	225	92	226	93
rect	228	92	229	93
rect	246	92	247	93
rect	249	92	250	93
rect	252	92	253	93
rect	264	92	265	93
rect	267	92	268	93
rect	270	92	271	93
rect	279	92	280	93
rect	288	92	289	93
rect	291	92	292	93
rect	294	92	295	93
rect	297	92	298	93
rect	300	92	301	93
rect	306	92	307	93
rect	309	92	310	93
rect	315	92	316	93
rect	318	92	319	93
rect	324	92	325	93
rect	330	92	331	93
rect	333	92	334	93
rect	339	92	340	93
rect	348	92	349	93
rect	357	92	358	93
rect	360	92	361	93
rect	369	92	370	93
rect	396	92	397	93
rect	11	93	12	94
rect	34	93	35	94
rect	37	93	38	94
rect	40	93	41	94
rect	50	93	51	94
rect	56	93	57	94
rect	59	93	60	94
rect	68	93	69	94
rect	77	93	78	94
rect	86	93	87	94
rect	112	93	113	94
rect	130	93	131	94
rect	136	93	137	94
rect	139	93	140	94
rect	142	93	143	94
rect	148	93	149	94
rect	164	93	165	94
rect	167	93	168	94
rect	173	93	174	94
rect	176	93	177	94
rect	179	93	180	94
rect	188	93	189	94
rect	194	93	195	94
rect	200	93	201	94
rect	203	93	204	94
rect	206	93	207	94
rect	209	93	210	94
rect	219	93	220	94
rect	225	93	226	94
rect	228	93	229	94
rect	246	93	247	94
rect	249	93	250	94
rect	252	93	253	94
rect	264	93	265	94
rect	270	93	271	94
rect	288	93	289	94
rect	291	93	292	94
rect	294	93	295	94
rect	297	93	298	94
rect	300	93	301	94
rect	306	93	307	94
rect	315	93	316	94
rect	318	93	319	94
rect	324	93	325	94
rect	330	93	331	94
rect	333	93	334	94
rect	339	93	340	94
rect	348	93	349	94
rect	357	93	358	94
rect	360	93	361	94
rect	369	93	370	94
rect	396	93	397	94
rect	11	94	12	95
rect	28	94	29	95
rect	31	94	32	95
rect	34	94	35	95
rect	37	94	38	95
rect	40	94	41	95
rect	50	94	51	95
rect	56	94	57	95
rect	59	94	60	95
rect	68	94	69	95
rect	77	94	78	95
rect	86	94	87	95
rect	89	94	90	95
rect	112	94	113	95
rect	121	94	122	95
rect	130	94	131	95
rect	136	94	137	95
rect	139	94	140	95
rect	142	94	143	95
rect	148	94	149	95
rect	151	94	152	95
rect	164	94	165	95
rect	167	94	168	95
rect	173	94	174	95
rect	176	94	177	95
rect	179	94	180	95
rect	188	94	189	95
rect	191	94	192	95
rect	194	94	195	95
rect	200	94	201	95
rect	203	94	204	95
rect	206	94	207	95
rect	209	94	210	95
rect	219	94	220	95
rect	222	94	223	95
rect	225	94	226	95
rect	228	94	229	95
rect	231	94	232	95
rect	246	94	247	95
rect	249	94	250	95
rect	252	94	253	95
rect	255	94	256	95
rect	258	94	259	95
rect	261	94	262	95
rect	264	94	265	95
rect	270	94	271	95
rect	273	94	274	95
rect	276	94	277	95
rect	288	94	289	95
rect	291	94	292	95
rect	294	94	295	95
rect	297	94	298	95
rect	300	94	301	95
rect	306	94	307	95
rect	315	94	316	95
rect	318	94	319	95
rect	321	94	322	95
rect	324	94	325	95
rect	330	94	331	95
rect	333	94	334	95
rect	339	94	340	95
rect	348	94	349	95
rect	357	94	358	95
rect	360	94	361	95
rect	369	94	370	95
rect	396	94	397	95
rect	28	95	29	96
rect	31	95	32	96
rect	34	95	35	96
rect	37	95	38	96
rect	40	95	41	96
rect	50	95	51	96
rect	56	95	57	96
rect	59	95	60	96
rect	68	95	69	96
rect	77	95	78	96
rect	86	95	87	96
rect	89	95	90	96
rect	112	95	113	96
rect	121	95	122	96
rect	130	95	131	96
rect	136	95	137	96
rect	139	95	140	96
rect	142	95	143	96
rect	148	95	149	96
rect	151	95	152	96
rect	164	95	165	96
rect	167	95	168	96
rect	173	95	174	96
rect	176	95	177	96
rect	179	95	180	96
rect	188	95	189	96
rect	191	95	192	96
rect	194	95	195	96
rect	200	95	201	96
rect	203	95	204	96
rect	219	95	220	96
rect	222	95	223	96
rect	225	95	226	96
rect	228	95	229	96
rect	231	95	232	96
rect	249	95	250	96
rect	252	95	253	96
rect	255	95	256	96
rect	258	95	259	96
rect	261	95	262	96
rect	264	95	265	96
rect	270	95	271	96
rect	273	95	274	96
rect	276	95	277	96
rect	288	95	289	96
rect	291	95	292	96
rect	294	95	295	96
rect	297	95	298	96
rect	306	95	307	96
rect	315	95	316	96
rect	318	95	319	96
rect	321	95	322	96
rect	324	95	325	96
rect	330	95	331	96
rect	333	95	334	96
rect	339	95	340	96
rect	348	95	349	96
rect	357	95	358	96
rect	360	95	361	96
rect	369	95	370	96
rect	396	95	397	96
rect	28	96	29	97
rect	31	96	32	97
rect	34	96	35	97
rect	37	96	38	97
rect	40	96	41	97
rect	50	96	51	97
rect	56	96	57	97
rect	59	96	60	97
rect	68	96	69	97
rect	77	96	78	97
rect	86	96	87	97
rect	89	96	90	97
rect	112	96	113	97
rect	121	96	122	97
rect	130	96	131	97
rect	136	96	137	97
rect	139	96	140	97
rect	142	96	143	97
rect	148	96	149	97
rect	151	96	152	97
rect	164	96	165	97
rect	167	96	168	97
rect	170	96	171	97
rect	173	96	174	97
rect	176	96	177	97
rect	179	96	180	97
rect	188	96	189	97
rect	191	96	192	97
rect	194	96	195	97
rect	197	96	198	97
rect	200	96	201	97
rect	203	96	204	97
rect	219	96	220	97
rect	222	96	223	97
rect	225	96	226	97
rect	228	96	229	97
rect	231	96	232	97
rect	240	96	241	97
rect	249	96	250	97
rect	252	96	253	97
rect	255	96	256	97
rect	258	96	259	97
rect	261	96	262	97
rect	264	96	265	97
rect	267	96	268	97
rect	270	96	271	97
rect	273	96	274	97
rect	276	96	277	97
rect	279	96	280	97
rect	285	96	286	97
rect	288	96	289	97
rect	291	96	292	97
rect	294	96	295	97
rect	297	96	298	97
rect	306	96	307	97
rect	315	96	316	97
rect	318	96	319	97
rect	321	96	322	97
rect	324	96	325	97
rect	330	96	331	97
rect	333	96	334	97
rect	336	96	337	97
rect	339	96	340	97
rect	348	96	349	97
rect	357	96	358	97
rect	360	96	361	97
rect	369	96	370	97
rect	378	96	379	97
rect	381	96	382	97
rect	384	96	385	97
rect	387	96	388	97
rect	396	96	397	97
rect	11	103	12	104
rect	28	103	29	104
rect	31	103	32	104
rect	34	103	35	104
rect	37	103	38	104
rect	40	103	41	104
rect	56	103	57	104
rect	59	103	60	104
rect	68	103	69	104
rect	77	103	78	104
rect	86	103	87	104
rect	89	103	90	104
rect	112	103	113	104
rect	121	103	122	104
rect	130	103	131	104
rect	139	103	140	104
rect	148	103	149	104
rect	151	103	152	104
rect	167	103	168	104
rect	170	103	171	104
rect	173	103	174	104
rect	176	103	177	104
rect	179	103	180	104
rect	185	103	186	104
rect	188	103	189	104
rect	191	103	192	104
rect	194	103	195	104
rect	197	103	198	104
rect	200	103	201	104
rect	203	103	204	104
rect	213	103	214	104
rect	219	103	220	104
rect	222	103	223	104
rect	225	103	226	104
rect	228	103	229	104
rect	231	103	232	104
rect	237	103	238	104
rect	240	103	241	104
rect	249	103	250	104
rect	252	103	253	104
rect	258	103	259	104
rect	261	103	262	104
rect	264	103	265	104
rect	267	103	268	104
rect	270	103	271	104
rect	273	103	274	104
rect	276	103	277	104
rect	285	103	286	104
rect	288	103	289	104
rect	291	103	292	104
rect	294	103	295	104
rect	297	103	298	104
rect	300	103	301	104
rect	306	103	307	104
rect	315	103	316	104
rect	318	103	319	104
rect	321	103	322	104
rect	327	103	328	104
rect	330	103	331	104
rect	333	103	334	104
rect	336	103	337	104
rect	339	103	340	104
rect	345	103	346	104
rect	348	103	349	104
rect	351	103	352	104
rect	357	103	358	104
rect	360	103	361	104
rect	369	103	370	104
rect	378	103	379	104
rect	387	103	388	104
rect	396	103	397	104
rect	402	103	403	104
rect	11	104	12	105
rect	28	104	29	105
rect	31	104	32	105
rect	34	104	35	105
rect	37	104	38	105
rect	40	104	41	105
rect	56	104	57	105
rect	59	104	60	105
rect	68	104	69	105
rect	77	104	78	105
rect	86	104	87	105
rect	89	104	90	105
rect	112	104	113	105
rect	121	104	122	105
rect	130	104	131	105
rect	139	104	140	105
rect	148	104	149	105
rect	151	104	152	105
rect	167	104	168	105
rect	170	104	171	105
rect	173	104	174	105
rect	176	104	177	105
rect	179	104	180	105
rect	185	104	186	105
rect	188	104	189	105
rect	191	104	192	105
rect	194	104	195	105
rect	197	104	198	105
rect	200	104	201	105
rect	203	104	204	105
rect	222	104	223	105
rect	225	104	226	105
rect	228	104	229	105
rect	231	104	232	105
rect	237	104	238	105
rect	240	104	241	105
rect	249	104	250	105
rect	252	104	253	105
rect	258	104	259	105
rect	261	104	262	105
rect	264	104	265	105
rect	267	104	268	105
rect	270	104	271	105
rect	273	104	274	105
rect	276	104	277	105
rect	285	104	286	105
rect	288	104	289	105
rect	291	104	292	105
rect	294	104	295	105
rect	297	104	298	105
rect	300	104	301	105
rect	306	104	307	105
rect	315	104	316	105
rect	318	104	319	105
rect	321	104	322	105
rect	327	104	328	105
rect	330	104	331	105
rect	333	104	334	105
rect	336	104	337	105
rect	345	104	346	105
rect	348	104	349	105
rect	351	104	352	105
rect	357	104	358	105
rect	360	104	361	105
rect	369	104	370	105
rect	387	104	388	105
rect	396	104	397	105
rect	402	104	403	105
rect	11	105	12	106
rect	28	105	29	106
rect	31	105	32	106
rect	34	105	35	106
rect	37	105	38	106
rect	40	105	41	106
rect	56	105	57	106
rect	59	105	60	106
rect	68	105	69	106
rect	77	105	78	106
rect	86	105	87	106
rect	89	105	90	106
rect	112	105	113	106
rect	121	105	122	106
rect	130	105	131	106
rect	139	105	140	106
rect	148	105	149	106
rect	151	105	152	106
rect	167	105	168	106
rect	170	105	171	106
rect	173	105	174	106
rect	176	105	177	106
rect	179	105	180	106
rect	185	105	186	106
rect	188	105	189	106
rect	191	105	192	106
rect	194	105	195	106
rect	197	105	198	106
rect	200	105	201	106
rect	203	105	204	106
rect	222	105	223	106
rect	225	105	226	106
rect	228	105	229	106
rect	231	105	232	106
rect	237	105	238	106
rect	240	105	241	106
rect	249	105	250	106
rect	252	105	253	106
rect	258	105	259	106
rect	261	105	262	106
rect	264	105	265	106
rect	267	105	268	106
rect	270	105	271	106
rect	273	105	274	106
rect	276	105	277	106
rect	285	105	286	106
rect	288	105	289	106
rect	291	105	292	106
rect	294	105	295	106
rect	297	105	298	106
rect	300	105	301	106
rect	306	105	307	106
rect	315	105	316	106
rect	318	105	319	106
rect	321	105	322	106
rect	327	105	328	106
rect	330	105	331	106
rect	333	105	334	106
rect	336	105	337	106
rect	342	105	343	106
rect	345	105	346	106
rect	348	105	349	106
rect	351	105	352	106
rect	357	105	358	106
rect	360	105	361	106
rect	369	105	370	106
rect	387	105	388	106
rect	396	105	397	106
rect	402	105	403	106
rect	419	105	420	106
rect	11	106	12	107
rect	28	106	29	107
rect	31	106	32	107
rect	34	106	35	107
rect	37	106	38	107
rect	40	106	41	107
rect	56	106	57	107
rect	59	106	60	107
rect	68	106	69	107
rect	77	106	78	107
rect	86	106	87	107
rect	89	106	90	107
rect	112	106	113	107
rect	121	106	122	107
rect	130	106	131	107
rect	139	106	140	107
rect	148	106	149	107
rect	151	106	152	107
rect	167	106	168	107
rect	170	106	171	107
rect	173	106	174	107
rect	176	106	177	107
rect	179	106	180	107
rect	185	106	186	107
rect	188	106	189	107
rect	191	106	192	107
rect	194	106	195	107
rect	197	106	198	107
rect	200	106	201	107
rect	222	106	223	107
rect	225	106	226	107
rect	228	106	229	107
rect	231	106	232	107
rect	237	106	238	107
rect	240	106	241	107
rect	249	106	250	107
rect	252	106	253	107
rect	258	106	259	107
rect	261	106	262	107
rect	264	106	265	107
rect	270	106	271	107
rect	273	106	274	107
rect	276	106	277	107
rect	285	106	286	107
rect	288	106	289	107
rect	291	106	292	107
rect	294	106	295	107
rect	300	106	301	107
rect	306	106	307	107
rect	315	106	316	107
rect	318	106	319	107
rect	321	106	322	107
rect	327	106	328	107
rect	333	106	334	107
rect	336	106	337	107
rect	342	106	343	107
rect	345	106	346	107
rect	348	106	349	107
rect	351	106	352	107
rect	357	106	358	107
rect	360	106	361	107
rect	369	106	370	107
rect	387	106	388	107
rect	396	106	397	107
rect	419	106	420	107
rect	11	107	12	108
rect	28	107	29	108
rect	31	107	32	108
rect	34	107	35	108
rect	37	107	38	108
rect	40	107	41	108
rect	56	107	57	108
rect	59	107	60	108
rect	68	107	69	108
rect	77	107	78	108
rect	86	107	87	108
rect	89	107	90	108
rect	112	107	113	108
rect	121	107	122	108
rect	130	107	131	108
rect	139	107	140	108
rect	148	107	149	108
rect	151	107	152	108
rect	167	107	168	108
rect	170	107	171	108
rect	173	107	174	108
rect	176	107	177	108
rect	179	107	180	108
rect	185	107	186	108
rect	188	107	189	108
rect	191	107	192	108
rect	194	107	195	108
rect	197	107	198	108
rect	200	107	201	108
rect	219	107	220	108
rect	222	107	223	108
rect	225	107	226	108
rect	228	107	229	108
rect	231	107	232	108
rect	237	107	238	108
rect	240	107	241	108
rect	249	107	250	108
rect	252	107	253	108
rect	258	107	259	108
rect	261	107	262	108
rect	264	107	265	108
rect	270	107	271	108
rect	273	107	274	108
rect	276	107	277	108
rect	279	107	280	108
rect	285	107	286	108
rect	288	107	289	108
rect	291	107	292	108
rect	294	107	295	108
rect	300	107	301	108
rect	303	107	304	108
rect	306	107	307	108
rect	315	107	316	108
rect	318	107	319	108
rect	321	107	322	108
rect	327	107	328	108
rect	333	107	334	108
rect	336	107	337	108
rect	342	107	343	108
rect	345	107	346	108
rect	348	107	349	108
rect	351	107	352	108
rect	357	107	358	108
rect	360	107	361	108
rect	369	107	370	108
rect	387	107	388	108
rect	396	107	397	108
rect	419	107	420	108
rect	11	108	12	109
rect	28	108	29	109
rect	31	108	32	109
rect	34	108	35	109
rect	37	108	38	109
rect	40	108	41	109
rect	56	108	57	109
rect	59	108	60	109
rect	68	108	69	109
rect	77	108	78	109
rect	86	108	87	109
rect	89	108	90	109
rect	112	108	113	109
rect	121	108	122	109
rect	130	108	131	109
rect	139	108	140	109
rect	148	108	149	109
rect	151	108	152	109
rect	167	108	168	109
rect	170	108	171	109
rect	173	108	174	109
rect	176	108	177	109
rect	179	108	180	109
rect	188	108	189	109
rect	191	108	192	109
rect	194	108	195	109
rect	197	108	198	109
rect	200	108	201	109
rect	219	108	220	109
rect	222	108	223	109
rect	225	108	226	109
rect	228	108	229	109
rect	231	108	232	109
rect	237	108	238	109
rect	240	108	241	109
rect	249	108	250	109
rect	252	108	253	109
rect	258	108	259	109
rect	264	108	265	109
rect	270	108	271	109
rect	273	108	274	109
rect	276	108	277	109
rect	279	108	280	109
rect	285	108	286	109
rect	288	108	289	109
rect	291	108	292	109
rect	294	108	295	109
rect	303	108	304	109
rect	315	108	316	109
rect	318	108	319	109
rect	321	108	322	109
rect	327	108	328	109
rect	333	108	334	109
rect	342	108	343	109
rect	345	108	346	109
rect	348	108	349	109
rect	351	108	352	109
rect	357	108	358	109
rect	360	108	361	109
rect	369	108	370	109
rect	396	108	397	109
rect	419	108	420	109
rect	11	109	12	110
rect	28	109	29	110
rect	31	109	32	110
rect	34	109	35	110
rect	37	109	38	110
rect	40	109	41	110
rect	56	109	57	110
rect	59	109	60	110
rect	68	109	69	110
rect	77	109	78	110
rect	86	109	87	110
rect	89	109	90	110
rect	112	109	113	110
rect	121	109	122	110
rect	130	109	131	110
rect	139	109	140	110
rect	148	109	149	110
rect	151	109	152	110
rect	167	109	168	110
rect	170	109	171	110
rect	173	109	174	110
rect	176	109	177	110
rect	179	109	180	110
rect	188	109	189	110
rect	191	109	192	110
rect	194	109	195	110
rect	197	109	198	110
rect	200	109	201	110
rect	204	109	205	110
rect	219	109	220	110
rect	222	109	223	110
rect	225	109	226	110
rect	228	109	229	110
rect	231	109	232	110
rect	237	109	238	110
rect	240	109	241	110
rect	249	109	250	110
rect	252	109	253	110
rect	258	109	259	110
rect	264	109	265	110
rect	270	109	271	110
rect	273	109	274	110
rect	276	109	277	110
rect	279	109	280	110
rect	285	109	286	110
rect	288	109	289	110
rect	291	109	292	110
rect	294	109	295	110
rect	297	109	298	110
rect	303	109	304	110
rect	315	109	316	110
rect	318	109	319	110
rect	321	109	322	110
rect	327	109	328	110
rect	333	109	334	110
rect	342	109	343	110
rect	345	109	346	110
rect	348	109	349	110
rect	351	109	352	110
rect	357	109	358	110
rect	360	109	361	110
rect	369	109	370	110
rect	378	109	379	110
rect	396	109	397	110
rect	402	109	403	110
rect	419	109	420	110
rect	11	110	12	111
rect	28	110	29	111
rect	31	110	32	111
rect	34	110	35	111
rect	37	110	38	111
rect	40	110	41	111
rect	56	110	57	111
rect	59	110	60	111
rect	68	110	69	111
rect	77	110	78	111
rect	86	110	87	111
rect	89	110	90	111
rect	112	110	113	111
rect	121	110	122	111
rect	130	110	131	111
rect	139	110	140	111
rect	148	110	149	111
rect	151	110	152	111
rect	167	110	168	111
rect	170	110	171	111
rect	173	110	174	111
rect	176	110	177	111
rect	179	110	180	111
rect	194	110	195	111
rect	197	110	198	111
rect	200	110	201	111
rect	204	110	205	111
rect	219	110	220	111
rect	222	110	223	111
rect	225	110	226	111
rect	228	110	229	111
rect	231	110	232	111
rect	237	110	238	111
rect	240	110	241	111
rect	252	110	253	111
rect	258	110	259	111
rect	270	110	271	111
rect	273	110	274	111
rect	276	110	277	111
rect	279	110	280	111
rect	285	110	286	111
rect	288	110	289	111
rect	291	110	292	111
rect	294	110	295	111
rect	297	110	298	111
rect	303	110	304	111
rect	315	110	316	111
rect	318	110	319	111
rect	327	110	328	111
rect	333	110	334	111
rect	342	110	343	111
rect	345	110	346	111
rect	348	110	349	111
rect	357	110	358	111
rect	360	110	361	111
rect	369	110	370	111
rect	378	110	379	111
rect	396	110	397	111
rect	402	110	403	111
rect	419	110	420	111
rect	11	111	12	112
rect	28	111	29	112
rect	31	111	32	112
rect	34	111	35	112
rect	37	111	38	112
rect	40	111	41	112
rect	56	111	57	112
rect	59	111	60	112
rect	68	111	69	112
rect	77	111	78	112
rect	86	111	87	112
rect	89	111	90	112
rect	112	111	113	112
rect	121	111	122	112
rect	130	111	131	112
rect	139	111	140	112
rect	148	111	149	112
rect	151	111	152	112
rect	167	111	168	112
rect	170	111	171	112
rect	173	111	174	112
rect	176	111	177	112
rect	179	111	180	112
rect	183	111	184	112
rect	194	111	195	112
rect	197	111	198	112
rect	200	111	201	112
rect	204	111	205	112
rect	213	111	214	112
rect	219	111	220	112
rect	222	111	223	112
rect	225	111	226	112
rect	228	111	229	112
rect	231	111	232	112
rect	237	111	238	112
rect	240	111	241	112
rect	252	111	253	112
rect	258	111	259	112
rect	261	111	262	112
rect	270	111	271	112
rect	273	111	274	112
rect	276	111	277	112
rect	279	111	280	112
rect	285	111	286	112
rect	288	111	289	112
rect	291	111	292	112
rect	294	111	295	112
rect	297	111	298	112
rect	303	111	304	112
rect	312	111	313	112
rect	315	111	316	112
rect	318	111	319	112
rect	327	111	328	112
rect	333	111	334	112
rect	339	111	340	112
rect	342	111	343	112
rect	345	111	346	112
rect	348	111	349	112
rect	357	111	358	112
rect	360	111	361	112
rect	369	111	370	112
rect	378	111	379	112
rect	387	111	388	112
rect	396	111	397	112
rect	402	111	403	112
rect	419	111	420	112
rect	11	112	12	113
rect	28	112	29	113
rect	31	112	32	113
rect	34	112	35	113
rect	37	112	38	113
rect	40	112	41	113
rect	56	112	57	113
rect	59	112	60	113
rect	68	112	69	113
rect	77	112	78	113
rect	86	112	87	113
rect	89	112	90	113
rect	112	112	113	113
rect	121	112	122	113
rect	130	112	131	113
rect	139	112	140	113
rect	148	112	149	113
rect	151	112	152	113
rect	167	112	168	113
rect	170	112	171	113
rect	176	112	177	113
rect	179	112	180	113
rect	183	112	184	113
rect	197	112	198	113
rect	200	112	201	113
rect	204	112	205	113
rect	213	112	214	113
rect	219	112	220	113
rect	225	112	226	113
rect	228	112	229	113
rect	231	112	232	113
rect	237	112	238	113
rect	240	112	241	113
rect	258	112	259	113
rect	261	112	262	113
rect	270	112	271	113
rect	273	112	274	113
rect	279	112	280	113
rect	285	112	286	113
rect	288	112	289	113
rect	291	112	292	113
rect	297	112	298	113
rect	303	112	304	113
rect	312	112	313	113
rect	315	112	316	113
rect	318	112	319	113
rect	327	112	328	113
rect	333	112	334	113
rect	339	112	340	113
rect	342	112	343	113
rect	345	112	346	113
rect	348	112	349	113
rect	360	112	361	113
rect	369	112	370	113
rect	378	112	379	113
rect	387	112	388	113
rect	396	112	397	113
rect	402	112	403	113
rect	419	112	420	113
rect	11	113	12	114
rect	28	113	29	114
rect	31	113	32	114
rect	34	113	35	114
rect	37	113	38	114
rect	40	113	41	114
rect	56	113	57	114
rect	59	113	60	114
rect	68	113	69	114
rect	77	113	78	114
rect	86	113	87	114
rect	89	113	90	114
rect	112	113	113	114
rect	121	113	122	114
rect	130	113	131	114
rect	139	113	140	114
rect	148	113	149	114
rect	151	113	152	114
rect	167	113	168	114
rect	170	113	171	114
rect	176	113	177	114
rect	179	113	180	114
rect	183	113	184	114
rect	189	113	190	114
rect	197	113	198	114
rect	200	113	201	114
rect	204	113	205	114
rect	213	113	214	114
rect	216	113	217	114
rect	219	113	220	114
rect	225	113	226	114
rect	228	113	229	114
rect	231	113	232	114
rect	237	113	238	114
rect	240	113	241	114
rect	243	113	244	114
rect	246	113	247	114
rect	258	113	259	114
rect	261	113	262	114
rect	264	113	265	114
rect	270	113	271	114
rect	273	113	274	114
rect	279	113	280	114
rect	285	113	286	114
rect	288	113	289	114
rect	291	113	292	114
rect	297	113	298	114
rect	303	113	304	114
rect	312	113	313	114
rect	315	113	316	114
rect	318	113	319	114
rect	327	113	328	114
rect	333	113	334	114
rect	339	113	340	114
rect	342	113	343	114
rect	345	113	346	114
rect	348	113	349	114
rect	351	113	352	114
rect	360	113	361	114
rect	369	113	370	114
rect	372	113	373	114
rect	378	113	379	114
rect	387	113	388	114
rect	396	113	397	114
rect	402	113	403	114
rect	419	113	420	114
rect	11	114	12	115
rect	28	114	29	115
rect	31	114	32	115
rect	34	114	35	115
rect	37	114	38	115
rect	40	114	41	115
rect	56	114	57	115
rect	59	114	60	115
rect	68	114	69	115
rect	77	114	78	115
rect	86	114	87	115
rect	89	114	90	115
rect	112	114	113	115
rect	121	114	122	115
rect	130	114	131	115
rect	139	114	140	115
rect	148	114	149	115
rect	167	114	168	115
rect	170	114	171	115
rect	176	114	177	115
rect	183	114	184	115
rect	189	114	190	115
rect	197	114	198	115
rect	204	114	205	115
rect	213	114	214	115
rect	216	114	217	115
rect	219	114	220	115
rect	225	114	226	115
rect	231	114	232	115
rect	237	114	238	115
rect	243	114	244	115
rect	246	114	247	115
rect	258	114	259	115
rect	261	114	262	115
rect	264	114	265	115
rect	270	114	271	115
rect	273	114	274	115
rect	279	114	280	115
rect	288	114	289	115
rect	291	114	292	115
rect	297	114	298	115
rect	303	114	304	115
rect	312	114	313	115
rect	315	114	316	115
rect	318	114	319	115
rect	327	114	328	115
rect	333	114	334	115
rect	339	114	340	115
rect	342	114	343	115
rect	348	114	349	115
rect	351	114	352	115
rect	360	114	361	115
rect	372	114	373	115
rect	378	114	379	115
rect	387	114	388	115
rect	396	114	397	115
rect	402	114	403	115
rect	419	114	420	115
rect	11	115	12	116
rect	28	115	29	116
rect	31	115	32	116
rect	34	115	35	116
rect	37	115	38	116
rect	40	115	41	116
rect	56	115	57	116
rect	59	115	60	116
rect	68	115	69	116
rect	77	115	78	116
rect	86	115	87	116
rect	89	115	90	116
rect	112	115	113	116
rect	121	115	122	116
rect	130	115	131	116
rect	139	115	140	116
rect	148	115	149	116
rect	167	115	168	116
rect	170	115	171	116
rect	174	115	175	116
rect	176	115	177	116
rect	183	115	184	116
rect	189	115	190	116
rect	195	115	196	116
rect	197	115	198	116
rect	204	115	205	116
rect	213	115	214	116
rect	216	115	217	116
rect	219	115	220	116
rect	222	115	223	116
rect	225	115	226	116
rect	231	115	232	116
rect	234	115	235	116
rect	237	115	238	116
rect	243	115	244	116
rect	246	115	247	116
rect	258	115	259	116
rect	261	115	262	116
rect	264	115	265	116
rect	270	115	271	116
rect	273	115	274	116
rect	276	115	277	116
rect	279	115	280	116
rect	288	115	289	116
rect	291	115	292	116
rect	297	115	298	116
rect	303	115	304	116
rect	312	115	313	116
rect	315	115	316	116
rect	318	115	319	116
rect	327	115	328	116
rect	333	115	334	116
rect	336	115	337	116
rect	339	115	340	116
rect	342	115	343	116
rect	348	115	349	116
rect	351	115	352	116
rect	360	115	361	116
rect	372	115	373	116
rect	378	115	379	116
rect	387	115	388	116
rect	396	115	397	116
rect	402	115	403	116
rect	419	115	420	116
rect	11	116	12	117
rect	28	116	29	117
rect	31	116	32	117
rect	34	116	35	117
rect	37	116	38	117
rect	40	116	41	117
rect	56	116	57	117
rect	59	116	60	117
rect	68	116	69	117
rect	77	116	78	117
rect	86	116	87	117
rect	121	116	122	117
rect	130	116	131	117
rect	139	116	140	117
rect	167	116	168	117
rect	170	116	171	117
rect	174	116	175	117
rect	183	116	184	117
rect	189	116	190	117
rect	195	116	196	117
rect	204	116	205	117
rect	213	116	214	117
rect	216	116	217	117
rect	219	116	220	117
rect	222	116	223	117
rect	231	116	232	117
rect	234	116	235	117
rect	237	116	238	117
rect	243	116	244	117
rect	246	116	247	117
rect	258	116	259	117
rect	261	116	262	117
rect	264	116	265	117
rect	270	116	271	117
rect	276	116	277	117
rect	279	116	280	117
rect	288	116	289	117
rect	291	116	292	117
rect	297	116	298	117
rect	303	116	304	117
rect	312	116	313	117
rect	318	116	319	117
rect	327	116	328	117
rect	333	116	334	117
rect	336	116	337	117
rect	339	116	340	117
rect	342	116	343	117
rect	348	116	349	117
rect	351	116	352	117
rect	360	116	361	117
rect	372	116	373	117
rect	378	116	379	117
rect	387	116	388	117
rect	396	116	397	117
rect	402	116	403	117
rect	419	116	420	117
rect	11	117	12	118
rect	28	117	29	118
rect	31	117	32	118
rect	34	117	35	118
rect	37	117	38	118
rect	40	117	41	118
rect	56	117	57	118
rect	59	117	60	118
rect	68	117	69	118
rect	77	117	78	118
rect	86	117	87	118
rect	92	117	93	118
rect	118	117	119	118
rect	121	117	122	118
rect	130	117	131	118
rect	139	117	140	118
rect	155	117	156	118
rect	167	117	168	118
rect	170	117	171	118
rect	174	117	175	118
rect	183	117	184	118
rect	189	117	190	118
rect	192	117	193	118
rect	195	117	196	118
rect	204	117	205	118
rect	207	117	208	118
rect	213	117	214	118
rect	216	117	217	118
rect	219	117	220	118
rect	222	117	223	118
rect	231	117	232	118
rect	234	117	235	118
rect	237	117	238	118
rect	243	117	244	118
rect	246	117	247	118
rect	258	117	259	118
rect	261	117	262	118
rect	264	117	265	118
rect	267	117	268	118
rect	270	117	271	118
rect	276	117	277	118
rect	279	117	280	118
rect	285	117	286	118
rect	288	117	289	118
rect	291	117	292	118
rect	294	117	295	118
rect	297	117	298	118
rect	303	117	304	118
rect	309	117	310	118
rect	312	117	313	118
rect	318	117	319	118
rect	327	117	328	118
rect	333	117	334	118
rect	336	117	337	118
rect	339	117	340	118
rect	342	117	343	118
rect	348	117	349	118
rect	351	117	352	118
rect	360	117	361	118
rect	363	117	364	118
rect	372	117	373	118
rect	378	117	379	118
rect	387	117	388	118
rect	396	117	397	118
rect	402	117	403	118
rect	419	117	420	118
rect	11	118	12	119
rect	28	118	29	119
rect	31	118	32	119
rect	34	118	35	119
rect	37	118	38	119
rect	56	118	57	119
rect	68	118	69	119
rect	77	118	78	119
rect	92	118	93	119
rect	118	118	119	119
rect	155	118	156	119
rect	167	118	168	119
rect	174	118	175	119
rect	183	118	184	119
rect	189	118	190	119
rect	192	118	193	119
rect	195	118	196	119
rect	204	118	205	119
rect	207	118	208	119
rect	213	118	214	119
rect	216	118	217	119
rect	219	118	220	119
rect	222	118	223	119
rect	231	118	232	119
rect	234	118	235	119
rect	237	118	238	119
rect	243	118	244	119
rect	246	118	247	119
rect	258	118	259	119
rect	261	118	262	119
rect	264	118	265	119
rect	267	118	268	119
rect	270	118	271	119
rect	276	118	277	119
rect	279	118	280	119
rect	285	118	286	119
rect	288	118	289	119
rect	291	118	292	119
rect	294	118	295	119
rect	297	118	298	119
rect	303	118	304	119
rect	309	118	310	119
rect	312	118	313	119
rect	318	118	319	119
rect	327	118	328	119
rect	333	118	334	119
rect	336	118	337	119
rect	339	118	340	119
rect	342	118	343	119
rect	348	118	349	119
rect	351	118	352	119
rect	360	118	361	119
rect	363	118	364	119
rect	372	118	373	119
rect	378	118	379	119
rect	387	118	388	119
rect	396	118	397	119
rect	402	118	403	119
rect	419	118	420	119
rect	11	119	12	120
rect	28	119	29	120
rect	31	119	32	120
rect	34	119	35	120
rect	37	119	38	120
rect	42	119	43	120
rect	56	119	57	120
rect	68	119	69	120
rect	70	119	71	120
rect	77	119	78	120
rect	89	119	90	120
rect	92	119	93	120
rect	109	119	110	120
rect	115	119	116	120
rect	118	119	119	120
rect	127	119	128	120
rect	136	119	137	120
rect	152	119	153	120
rect	155	119	156	120
rect	167	119	168	120
rect	174	119	175	120
rect	177	119	178	120
rect	183	119	184	120
rect	186	119	187	120
rect	189	119	190	120
rect	192	119	193	120
rect	195	119	196	120
rect	204	119	205	120
rect	207	119	208	120
rect	213	119	214	120
rect	216	119	217	120
rect	219	119	220	120
rect	222	119	223	120
rect	231	119	232	120
rect	234	119	235	120
rect	237	119	238	120
rect	243	119	244	120
rect	246	119	247	120
rect	258	119	259	120
rect	261	119	262	120
rect	264	119	265	120
rect	267	119	268	120
rect	270	119	271	120
rect	276	119	277	120
rect	279	119	280	120
rect	285	119	286	120
rect	288	119	289	120
rect	291	119	292	120
rect	294	119	295	120
rect	297	119	298	120
rect	303	119	304	120
rect	309	119	310	120
rect	312	119	313	120
rect	318	119	319	120
rect	327	119	328	120
rect	333	119	334	120
rect	336	119	337	120
rect	339	119	340	120
rect	342	119	343	120
rect	348	119	349	120
rect	351	119	352	120
rect	357	119	358	120
rect	360	119	361	120
rect	363	119	364	120
rect	372	119	373	120
rect	378	119	379	120
rect	387	119	388	120
rect	396	119	397	120
rect	402	119	403	120
rect	419	119	420	120
rect	11	120	12	121
rect	28	120	29	121
rect	31	120	32	121
rect	34	120	35	121
rect	42	120	43	121
rect	70	120	71	121
rect	89	120	90	121
rect	92	120	93	121
rect	109	120	110	121
rect	115	120	116	121
rect	118	120	119	121
rect	127	120	128	121
rect	136	120	137	121
rect	152	120	153	121
rect	155	120	156	121
rect	167	120	168	121
rect	174	120	175	121
rect	177	120	178	121
rect	183	120	184	121
rect	186	120	187	121
rect	189	120	190	121
rect	192	120	193	121
rect	195	120	196	121
rect	204	120	205	121
rect	207	120	208	121
rect	213	120	214	121
rect	216	120	217	121
rect	219	120	220	121
rect	222	120	223	121
rect	231	120	232	121
rect	234	120	235	121
rect	237	120	238	121
rect	243	120	244	121
rect	246	120	247	121
rect	258	120	259	121
rect	261	120	262	121
rect	264	120	265	121
rect	267	120	268	121
rect	270	120	271	121
rect	276	120	277	121
rect	279	120	280	121
rect	285	120	286	121
rect	288	120	289	121
rect	291	120	292	121
rect	294	120	295	121
rect	297	120	298	121
rect	303	120	304	121
rect	309	120	310	121
rect	312	120	313	121
rect	318	120	319	121
rect	327	120	328	121
rect	336	120	337	121
rect	339	120	340	121
rect	342	120	343	121
rect	348	120	349	121
rect	351	120	352	121
rect	357	120	358	121
rect	360	120	361	121
rect	363	120	364	121
rect	372	120	373	121
rect	378	120	379	121
rect	387	120	388	121
rect	396	120	397	121
rect	402	120	403	121
rect	419	120	420	121
rect	11	121	12	122
rect	28	121	29	122
rect	31	121	32	122
rect	34	121	35	122
rect	39	121	40	122
rect	42	121	43	122
rect	58	121	59	122
rect	61	121	62	122
rect	70	121	71	122
rect	86	121	87	122
rect	89	121	90	122
rect	92	121	93	122
rect	95	121	96	122
rect	109	121	110	122
rect	115	121	116	122
rect	118	121	119	122
rect	127	121	128	122
rect	136	121	137	122
rect	152	121	153	122
rect	155	121	156	122
rect	167	121	168	122
rect	174	121	175	122
rect	177	121	178	122
rect	183	121	184	122
rect	186	121	187	122
rect	189	121	190	122
rect	192	121	193	122
rect	195	121	196	122
rect	204	121	205	122
rect	207	121	208	122
rect	213	121	214	122
rect	216	121	217	122
rect	219	121	220	122
rect	222	121	223	122
rect	231	121	232	122
rect	234	121	235	122
rect	237	121	238	122
rect	243	121	244	122
rect	246	121	247	122
rect	258	121	259	122
rect	261	121	262	122
rect	264	121	265	122
rect	267	121	268	122
rect	270	121	271	122
rect	276	121	277	122
rect	279	121	280	122
rect	285	121	286	122
rect	288	121	289	122
rect	291	121	292	122
rect	294	121	295	122
rect	297	121	298	122
rect	303	121	304	122
rect	309	121	310	122
rect	312	121	313	122
rect	318	121	319	122
rect	321	121	322	122
rect	327	121	328	122
rect	336	121	337	122
rect	339	121	340	122
rect	342	121	343	122
rect	348	121	349	122
rect	351	121	352	122
rect	357	121	358	122
rect	360	121	361	122
rect	363	121	364	122
rect	366	121	367	122
rect	372	121	373	122
rect	378	121	379	122
rect	387	121	388	122
rect	396	121	397	122
rect	402	121	403	122
rect	419	121	420	122
rect	11	122	12	123
rect	28	122	29	123
rect	34	122	35	123
rect	39	122	40	123
rect	42	122	43	123
rect	58	122	59	123
rect	61	122	62	123
rect	70	122	71	123
rect	86	122	87	123
rect	89	122	90	123
rect	92	122	93	123
rect	95	122	96	123
rect	109	122	110	123
rect	115	122	116	123
rect	118	122	119	123
rect	127	122	128	123
rect	136	122	137	123
rect	152	122	153	123
rect	155	122	156	123
rect	174	122	175	123
rect	177	122	178	123
rect	183	122	184	123
rect	186	122	187	123
rect	189	122	190	123
rect	192	122	193	123
rect	195	122	196	123
rect	204	122	205	123
rect	207	122	208	123
rect	213	122	214	123
rect	216	122	217	123
rect	219	122	220	123
rect	222	122	223	123
rect	234	122	235	123
rect	243	122	244	123
rect	246	122	247	123
rect	258	122	259	123
rect	261	122	262	123
rect	264	122	265	123
rect	267	122	268	123
rect	270	122	271	123
rect	276	122	277	123
rect	279	122	280	123
rect	285	122	286	123
rect	288	122	289	123
rect	291	122	292	123
rect	294	122	295	123
rect	297	122	298	123
rect	303	122	304	123
rect	309	122	310	123
rect	312	122	313	123
rect	321	122	322	123
rect	327	122	328	123
rect	336	122	337	123
rect	339	122	340	123
rect	342	122	343	123
rect	348	122	349	123
rect	351	122	352	123
rect	357	122	358	123
rect	363	122	364	123
rect	366	122	367	123
rect	372	122	373	123
rect	378	122	379	123
rect	387	122	388	123
rect	396	122	397	123
rect	402	122	403	123
rect	419	122	420	123
rect	11	123	12	124
rect	28	123	29	124
rect	34	123	35	124
rect	39	123	40	124
rect	42	123	43	124
rect	58	123	59	124
rect	61	123	62	124
rect	70	123	71	124
rect	86	123	87	124
rect	89	123	90	124
rect	92	123	93	124
rect	95	123	96	124
rect	109	123	110	124
rect	115	123	116	124
rect	118	123	119	124
rect	127	123	128	124
rect	136	123	137	124
rect	152	123	153	124
rect	155	123	156	124
rect	158	123	159	124
rect	174	123	175	124
rect	177	123	178	124
rect	183	123	184	124
rect	186	123	187	124
rect	189	123	190	124
rect	192	123	193	124
rect	195	123	196	124
rect	204	123	205	124
rect	207	123	208	124
rect	210	123	211	124
rect	213	123	214	124
rect	216	123	217	124
rect	219	123	220	124
rect	222	123	223	124
rect	225	123	226	124
rect	234	123	235	124
rect	243	123	244	124
rect	246	123	247	124
rect	258	123	259	124
rect	261	123	262	124
rect	264	123	265	124
rect	267	123	268	124
rect	270	123	271	124
rect	276	123	277	124
rect	279	123	280	124
rect	285	123	286	124
rect	288	123	289	124
rect	291	123	292	124
rect	294	123	295	124
rect	297	123	298	124
rect	303	123	304	124
rect	309	123	310	124
rect	312	123	313	124
rect	315	123	316	124
rect	321	123	322	124
rect	327	123	328	124
rect	333	123	334	124
rect	336	123	337	124
rect	339	123	340	124
rect	342	123	343	124
rect	348	123	349	124
rect	351	123	352	124
rect	357	123	358	124
rect	363	123	364	124
rect	366	123	367	124
rect	369	123	370	124
rect	372	123	373	124
rect	378	123	379	124
rect	387	123	388	124
rect	396	123	397	124
rect	402	123	403	124
rect	419	123	420	124
rect	11	124	12	125
rect	39	124	40	125
rect	42	124	43	125
rect	58	124	59	125
rect	61	124	62	125
rect	70	124	71	125
rect	86	124	87	125
rect	89	124	90	125
rect	92	124	93	125
rect	95	124	96	125
rect	109	124	110	125
rect	115	124	116	125
rect	118	124	119	125
rect	127	124	128	125
rect	136	124	137	125
rect	152	124	153	125
rect	155	124	156	125
rect	158	124	159	125
rect	174	124	175	125
rect	177	124	178	125
rect	183	124	184	125
rect	186	124	187	125
rect	189	124	190	125
rect	192	124	193	125
rect	195	124	196	125
rect	204	124	205	125
rect	207	124	208	125
rect	210	124	211	125
rect	213	124	214	125
rect	216	124	217	125
rect	219	124	220	125
rect	222	124	223	125
rect	225	124	226	125
rect	234	124	235	125
rect	243	124	244	125
rect	246	124	247	125
rect	258	124	259	125
rect	261	124	262	125
rect	264	124	265	125
rect	267	124	268	125
rect	276	124	277	125
rect	279	124	280	125
rect	285	124	286	125
rect	288	124	289	125
rect	294	124	295	125
rect	297	124	298	125
rect	303	124	304	125
rect	309	124	310	125
rect	312	124	313	125
rect	315	124	316	125
rect	321	124	322	125
rect	327	124	328	125
rect	333	124	334	125
rect	336	124	337	125
rect	339	124	340	125
rect	342	124	343	125
rect	348	124	349	125
rect	351	124	352	125
rect	357	124	358	125
rect	363	124	364	125
rect	366	124	367	125
rect	369	124	370	125
rect	372	124	373	125
rect	378	124	379	125
rect	387	124	388	125
rect	402	124	403	125
rect	419	124	420	125
rect	11	125	12	126
rect	18	125	19	126
rect	21	125	22	126
rect	30	125	31	126
rect	39	125	40	126
rect	42	125	43	126
rect	58	125	59	126
rect	61	125	62	126
rect	70	125	71	126
rect	86	125	87	126
rect	89	125	90	126
rect	92	125	93	126
rect	95	125	96	126
rect	109	125	110	126
rect	115	125	116	126
rect	118	125	119	126
rect	127	125	128	126
rect	136	125	137	126
rect	152	125	153	126
rect	155	125	156	126
rect	158	125	159	126
rect	174	125	175	126
rect	177	125	178	126
rect	183	125	184	126
rect	186	125	187	126
rect	189	125	190	126
rect	192	125	193	126
rect	195	125	196	126
rect	204	125	205	126
rect	207	125	208	126
rect	210	125	211	126
rect	213	125	214	126
rect	216	125	217	126
rect	219	125	220	126
rect	222	125	223	126
rect	225	125	226	126
rect	234	125	235	126
rect	243	125	244	126
rect	246	125	247	126
rect	249	125	250	126
rect	258	125	259	126
rect	261	125	262	126
rect	264	125	265	126
rect	267	125	268	126
rect	276	125	277	126
rect	279	125	280	126
rect	282	125	283	126
rect	285	125	286	126
rect	288	125	289	126
rect	294	125	295	126
rect	297	125	298	126
rect	303	125	304	126
rect	309	125	310	126
rect	312	125	313	126
rect	315	125	316	126
rect	318	125	319	126
rect	321	125	322	126
rect	327	125	328	126
rect	333	125	334	126
rect	336	125	337	126
rect	339	125	340	126
rect	342	125	343	126
rect	348	125	349	126
rect	351	125	352	126
rect	354	125	355	126
rect	357	125	358	126
rect	360	125	361	126
rect	363	125	364	126
rect	366	125	367	126
rect	369	125	370	126
rect	372	125	373	126
rect	378	125	379	126
rect	387	125	388	126
rect	402	125	403	126
rect	416	125	417	126
rect	419	125	420	126
rect	18	126	19	127
rect	21	126	22	127
rect	30	126	31	127
rect	39	126	40	127
rect	42	126	43	127
rect	58	126	59	127
rect	61	126	62	127
rect	70	126	71	127
rect	86	126	87	127
rect	89	126	90	127
rect	92	126	93	127
rect	95	126	96	127
rect	109	126	110	127
rect	115	126	116	127
rect	118	126	119	127
rect	127	126	128	127
rect	136	126	137	127
rect	152	126	153	127
rect	155	126	156	127
rect	158	126	159	127
rect	174	126	175	127
rect	177	126	178	127
rect	183	126	184	127
rect	186	126	187	127
rect	189	126	190	127
rect	192	126	193	127
rect	195	126	196	127
rect	204	126	205	127
rect	207	126	208	127
rect	210	126	211	127
rect	213	126	214	127
rect	216	126	217	127
rect	219	126	220	127
rect	222	126	223	127
rect	225	126	226	127
rect	234	126	235	127
rect	243	126	244	127
rect	246	126	247	127
rect	249	126	250	127
rect	261	126	262	127
rect	264	126	265	127
rect	267	126	268	127
rect	276	126	277	127
rect	279	126	280	127
rect	282	126	283	127
rect	285	126	286	127
rect	294	126	295	127
rect	297	126	298	127
rect	303	126	304	127
rect	309	126	310	127
rect	312	126	313	127
rect	315	126	316	127
rect	318	126	319	127
rect	321	126	322	127
rect	333	126	334	127
rect	336	126	337	127
rect	339	126	340	127
rect	342	126	343	127
rect	351	126	352	127
rect	354	126	355	127
rect	357	126	358	127
rect	360	126	361	127
rect	363	126	364	127
rect	366	126	367	127
rect	369	126	370	127
rect	372	126	373	127
rect	378	126	379	127
rect	387	126	388	127
rect	402	126	403	127
rect	416	126	417	127
rect	419	126	420	127
rect	18	127	19	128
rect	21	127	22	128
rect	30	127	31	128
rect	39	127	40	128
rect	42	127	43	128
rect	58	127	59	128
rect	61	127	62	128
rect	70	127	71	128
rect	86	127	87	128
rect	89	127	90	128
rect	92	127	93	128
rect	95	127	96	128
rect	109	127	110	128
rect	115	127	116	128
rect	118	127	119	128
rect	127	127	128	128
rect	136	127	137	128
rect	152	127	153	128
rect	155	127	156	128
rect	158	127	159	128
rect	174	127	175	128
rect	177	127	178	128
rect	183	127	184	128
rect	186	127	187	128
rect	189	127	190	128
rect	192	127	193	128
rect	195	127	196	128
rect	204	127	205	128
rect	207	127	208	128
rect	210	127	211	128
rect	213	127	214	128
rect	216	127	217	128
rect	219	127	220	128
rect	222	127	223	128
rect	225	127	226	128
rect	234	127	235	128
rect	243	127	244	128
rect	246	127	247	128
rect	249	127	250	128
rect	252	127	253	128
rect	261	127	262	128
rect	264	127	265	128
rect	267	127	268	128
rect	273	127	274	128
rect	276	127	277	128
rect	279	127	280	128
rect	282	127	283	128
rect	285	127	286	128
rect	294	127	295	128
rect	297	127	298	128
rect	300	127	301	128
rect	303	127	304	128
rect	309	127	310	128
rect	312	127	313	128
rect	315	127	316	128
rect	318	127	319	128
rect	321	127	322	128
rect	330	127	331	128
rect	333	127	334	128
rect	336	127	337	128
rect	339	127	340	128
rect	342	127	343	128
rect	351	127	352	128
rect	354	127	355	128
rect	357	127	358	128
rect	360	127	361	128
rect	363	127	364	128
rect	366	127	367	128
rect	369	127	370	128
rect	372	127	373	128
rect	378	127	379	128
rect	387	127	388	128
rect	396	127	397	128
rect	402	127	403	128
rect	416	127	417	128
rect	419	127	420	128
rect	21	134	22	135
rect	30	134	31	135
rect	36	134	37	135
rect	39	134	40	135
rect	42	134	43	135
rect	55	134	56	135
rect	58	134	59	135
rect	61	134	62	135
rect	70	134	71	135
rect	86	134	87	135
rect	89	134	90	135
rect	92	134	93	135
rect	112	134	113	135
rect	115	134	116	135
rect	118	134	119	135
rect	127	134	128	135
rect	130	134	131	135
rect	136	134	137	135
rect	152	134	153	135
rect	155	134	156	135
rect	158	134	159	135
rect	174	134	175	135
rect	177	134	178	135
rect	186	134	187	135
rect	189	134	190	135
rect	192	134	193	135
rect	195	134	196	135
rect	204	134	205	135
rect	207	134	208	135
rect	210	134	211	135
rect	213	134	214	135
rect	216	134	217	135
rect	219	134	220	135
rect	222	134	223	135
rect	225	134	226	135
rect	228	134	229	135
rect	234	134	235	135
rect	237	134	238	135
rect	243	134	244	135
rect	246	134	247	135
rect	249	134	250	135
rect	252	134	253	135
rect	261	134	262	135
rect	264	134	265	135
rect	267	134	268	135
rect	273	134	274	135
rect	276	134	277	135
rect	279	134	280	135
rect	282	134	283	135
rect	285	134	286	135
rect	294	134	295	135
rect	297	134	298	135
rect	300	134	301	135
rect	303	134	304	135
rect	312	134	313	135
rect	315	134	316	135
rect	318	134	319	135
rect	321	134	322	135
rect	324	134	325	135
rect	330	134	331	135
rect	333	134	334	135
rect	336	134	337	135
rect	339	134	340	135
rect	342	134	343	135
rect	351	134	352	135
rect	354	134	355	135
rect	357	134	358	135
rect	363	134	364	135
rect	366	134	367	135
rect	369	134	370	135
rect	375	134	376	135
rect	378	134	379	135
rect	387	134	388	135
rect	396	134	397	135
rect	402	134	403	135
rect	419	134	420	135
rect	21	135	22	136
rect	30	135	31	136
rect	36	135	37	136
rect	39	135	40	136
rect	42	135	43	136
rect	55	135	56	136
rect	58	135	59	136
rect	61	135	62	136
rect	70	135	71	136
rect	86	135	87	136
rect	89	135	90	136
rect	92	135	93	136
rect	112	135	113	136
rect	115	135	116	136
rect	118	135	119	136
rect	127	135	128	136
rect	130	135	131	136
rect	136	135	137	136
rect	152	135	153	136
rect	155	135	156	136
rect	158	135	159	136
rect	174	135	175	136
rect	177	135	178	136
rect	186	135	187	136
rect	189	135	190	136
rect	192	135	193	136
rect	195	135	196	136
rect	204	135	205	136
rect	207	135	208	136
rect	210	135	211	136
rect	213	135	214	136
rect	219	135	220	136
rect	222	135	223	136
rect	225	135	226	136
rect	228	135	229	136
rect	234	135	235	136
rect	237	135	238	136
rect	243	135	244	136
rect	246	135	247	136
rect	249	135	250	136
rect	252	135	253	136
rect	261	135	262	136
rect	264	135	265	136
rect	267	135	268	136
rect	273	135	274	136
rect	276	135	277	136
rect	279	135	280	136
rect	282	135	283	136
rect	285	135	286	136
rect	294	135	295	136
rect	297	135	298	136
rect	300	135	301	136
rect	303	135	304	136
rect	312	135	313	136
rect	315	135	316	136
rect	318	135	319	136
rect	321	135	322	136
rect	324	135	325	136
rect	330	135	331	136
rect	333	135	334	136
rect	336	135	337	136
rect	339	135	340	136
rect	342	135	343	136
rect	351	135	352	136
rect	354	135	355	136
rect	357	135	358	136
rect	363	135	364	136
rect	366	135	367	136
rect	369	135	370	136
rect	375	135	376	136
rect	378	135	379	136
rect	387	135	388	136
rect	396	135	397	136
rect	402	135	403	136
rect	419	135	420	136
rect	21	136	22	137
rect	30	136	31	137
rect	36	136	37	137
rect	39	136	40	137
rect	42	136	43	137
rect	55	136	56	137
rect	58	136	59	137
rect	61	136	62	137
rect	70	136	71	137
rect	86	136	87	137
rect	89	136	90	137
rect	92	136	93	137
rect	112	136	113	137
rect	115	136	116	137
rect	118	136	119	137
rect	127	136	128	137
rect	130	136	131	137
rect	136	136	137	137
rect	152	136	153	137
rect	155	136	156	137
rect	158	136	159	137
rect	174	136	175	137
rect	177	136	178	137
rect	186	136	187	137
rect	189	136	190	137
rect	192	136	193	137
rect	195	136	196	137
rect	204	136	205	137
rect	207	136	208	137
rect	210	136	211	137
rect	213	136	214	137
rect	219	136	220	137
rect	222	136	223	137
rect	225	136	226	137
rect	228	136	229	137
rect	231	136	232	137
rect	234	136	235	137
rect	237	136	238	137
rect	243	136	244	137
rect	246	136	247	137
rect	249	136	250	137
rect	252	136	253	137
rect	261	136	262	137
rect	264	136	265	137
rect	267	136	268	137
rect	273	136	274	137
rect	276	136	277	137
rect	279	136	280	137
rect	282	136	283	137
rect	285	136	286	137
rect	294	136	295	137
rect	297	136	298	137
rect	300	136	301	137
rect	303	136	304	137
rect	312	136	313	137
rect	315	136	316	137
rect	318	136	319	137
rect	321	136	322	137
rect	324	136	325	137
rect	330	136	331	137
rect	333	136	334	137
rect	336	136	337	137
rect	339	136	340	137
rect	342	136	343	137
rect	351	136	352	137
rect	354	136	355	137
rect	357	136	358	137
rect	363	136	364	137
rect	366	136	367	137
rect	369	136	370	137
rect	375	136	376	137
rect	378	136	379	137
rect	387	136	388	137
rect	396	136	397	137
rect	402	136	403	137
rect	419	136	420	137
rect	21	137	22	138
rect	30	137	31	138
rect	36	137	37	138
rect	39	137	40	138
rect	42	137	43	138
rect	55	137	56	138
rect	58	137	59	138
rect	61	137	62	138
rect	70	137	71	138
rect	86	137	87	138
rect	89	137	90	138
rect	92	137	93	138
rect	112	137	113	138
rect	115	137	116	138
rect	118	137	119	138
rect	127	137	128	138
rect	130	137	131	138
rect	136	137	137	138
rect	152	137	153	138
rect	155	137	156	138
rect	158	137	159	138
rect	174	137	175	138
rect	177	137	178	138
rect	186	137	187	138
rect	189	137	190	138
rect	192	137	193	138
rect	195	137	196	138
rect	204	137	205	138
rect	207	137	208	138
rect	213	137	214	138
rect	219	137	220	138
rect	222	137	223	138
rect	228	137	229	138
rect	231	137	232	138
rect	234	137	235	138
rect	243	137	244	138
rect	246	137	247	138
rect	249	137	250	138
rect	252	137	253	138
rect	264	137	265	138
rect	267	137	268	138
rect	273	137	274	138
rect	276	137	277	138
rect	279	137	280	138
rect	282	137	283	138
rect	285	137	286	138
rect	294	137	295	138
rect	297	137	298	138
rect	300	137	301	138
rect	303	137	304	138
rect	312	137	313	138
rect	318	137	319	138
rect	321	137	322	138
rect	324	137	325	138
rect	330	137	331	138
rect	333	137	334	138
rect	336	137	337	138
rect	339	137	340	138
rect	342	137	343	138
rect	351	137	352	138
rect	354	137	355	138
rect	357	137	358	138
rect	363	137	364	138
rect	366	137	367	138
rect	369	137	370	138
rect	375	137	376	138
rect	378	137	379	138
rect	387	137	388	138
rect	396	137	397	138
rect	402	137	403	138
rect	419	137	420	138
rect	21	138	22	139
rect	30	138	31	139
rect	36	138	37	139
rect	39	138	40	139
rect	42	138	43	139
rect	55	138	56	139
rect	58	138	59	139
rect	61	138	62	139
rect	70	138	71	139
rect	86	138	87	139
rect	89	138	90	139
rect	92	138	93	139
rect	112	138	113	139
rect	115	138	116	139
rect	118	138	119	139
rect	127	138	128	139
rect	130	138	131	139
rect	136	138	137	139
rect	152	138	153	139
rect	155	138	156	139
rect	158	138	159	139
rect	174	138	175	139
rect	177	138	178	139
rect	186	138	187	139
rect	189	138	190	139
rect	192	138	193	139
rect	195	138	196	139
rect	201	138	202	139
rect	204	138	205	139
rect	207	138	208	139
rect	213	138	214	139
rect	216	138	217	139
rect	219	138	220	139
rect	222	138	223	139
rect	228	138	229	139
rect	231	138	232	139
rect	234	138	235	139
rect	243	138	244	139
rect	246	138	247	139
rect	249	138	250	139
rect	252	138	253	139
rect	264	138	265	139
rect	267	138	268	139
rect	273	138	274	139
rect	276	138	277	139
rect	279	138	280	139
rect	282	138	283	139
rect	285	138	286	139
rect	294	138	295	139
rect	297	138	298	139
rect	300	138	301	139
rect	303	138	304	139
rect	306	138	307	139
rect	312	138	313	139
rect	318	138	319	139
rect	321	138	322	139
rect	324	138	325	139
rect	330	138	331	139
rect	333	138	334	139
rect	336	138	337	139
rect	339	138	340	139
rect	342	138	343	139
rect	351	138	352	139
rect	354	138	355	139
rect	357	138	358	139
rect	363	138	364	139
rect	366	138	367	139
rect	369	138	370	139
rect	375	138	376	139
rect	378	138	379	139
rect	387	138	388	139
rect	396	138	397	139
rect	402	138	403	139
rect	419	138	420	139
rect	21	139	22	140
rect	30	139	31	140
rect	36	139	37	140
rect	39	139	40	140
rect	42	139	43	140
rect	55	139	56	140
rect	58	139	59	140
rect	61	139	62	140
rect	70	139	71	140
rect	86	139	87	140
rect	89	139	90	140
rect	92	139	93	140
rect	112	139	113	140
rect	115	139	116	140
rect	118	139	119	140
rect	127	139	128	140
rect	130	139	131	140
rect	136	139	137	140
rect	152	139	153	140
rect	155	139	156	140
rect	158	139	159	140
rect	174	139	175	140
rect	177	139	178	140
rect	186	139	187	140
rect	189	139	190	140
rect	192	139	193	140
rect	195	139	196	140
rect	201	139	202	140
rect	204	139	205	140
rect	207	139	208	140
rect	213	139	214	140
rect	216	139	217	140
rect	219	139	220	140
rect	222	139	223	140
rect	228	139	229	140
rect	231	139	232	140
rect	234	139	235	140
rect	243	139	244	140
rect	246	139	247	140
rect	249	139	250	140
rect	252	139	253	140
rect	264	139	265	140
rect	273	139	274	140
rect	279	139	280	140
rect	282	139	283	140
rect	285	139	286	140
rect	294	139	295	140
rect	300	139	301	140
rect	303	139	304	140
rect	306	139	307	140
rect	312	139	313	140
rect	318	139	319	140
rect	321	139	322	140
rect	324	139	325	140
rect	330	139	331	140
rect	333	139	334	140
rect	336	139	337	140
rect	339	139	340	140
rect	342	139	343	140
rect	351	139	352	140
rect	354	139	355	140
rect	357	139	358	140
rect	363	139	364	140
rect	366	139	367	140
rect	369	139	370	140
rect	375	139	376	140
rect	378	139	379	140
rect	387	139	388	140
rect	396	139	397	140
rect	402	139	403	140
rect	419	139	420	140
rect	21	140	22	141
rect	30	140	31	141
rect	36	140	37	141
rect	39	140	40	141
rect	42	140	43	141
rect	55	140	56	141
rect	58	140	59	141
rect	61	140	62	141
rect	70	140	71	141
rect	86	140	87	141
rect	89	140	90	141
rect	92	140	93	141
rect	112	140	113	141
rect	115	140	116	141
rect	118	140	119	141
rect	127	140	128	141
rect	130	140	131	141
rect	136	140	137	141
rect	149	140	150	141
rect	152	140	153	141
rect	155	140	156	141
rect	158	140	159	141
rect	174	140	175	141
rect	177	140	178	141
rect	186	140	187	141
rect	189	140	190	141
rect	192	140	193	141
rect	195	140	196	141
rect	201	140	202	141
rect	204	140	205	141
rect	207	140	208	141
rect	213	140	214	141
rect	216	140	217	141
rect	219	140	220	141
rect	222	140	223	141
rect	228	140	229	141
rect	231	140	232	141
rect	234	140	235	141
rect	243	140	244	141
rect	246	140	247	141
rect	249	140	250	141
rect	252	140	253	141
rect	264	140	265	141
rect	273	140	274	141
rect	279	140	280	141
rect	282	140	283	141
rect	285	140	286	141
rect	288	140	289	141
rect	294	140	295	141
rect	300	140	301	141
rect	303	140	304	141
rect	306	140	307	141
rect	312	140	313	141
rect	315	140	316	141
rect	318	140	319	141
rect	321	140	322	141
rect	324	140	325	141
rect	330	140	331	141
rect	333	140	334	141
rect	336	140	337	141
rect	339	140	340	141
rect	342	140	343	141
rect	351	140	352	141
rect	354	140	355	141
rect	357	140	358	141
rect	363	140	364	141
rect	366	140	367	141
rect	369	140	370	141
rect	375	140	376	141
rect	378	140	379	141
rect	387	140	388	141
rect	396	140	397	141
rect	402	140	403	141
rect	419	140	420	141
rect	21	141	22	142
rect	30	141	31	142
rect	36	141	37	142
rect	39	141	40	142
rect	42	141	43	142
rect	55	141	56	142
rect	58	141	59	142
rect	61	141	62	142
rect	70	141	71	142
rect	86	141	87	142
rect	89	141	90	142
rect	92	141	93	142
rect	112	141	113	142
rect	115	141	116	142
rect	118	141	119	142
rect	127	141	128	142
rect	130	141	131	142
rect	136	141	137	142
rect	149	141	150	142
rect	152	141	153	142
rect	155	141	156	142
rect	158	141	159	142
rect	174	141	175	142
rect	177	141	178	142
rect	186	141	187	142
rect	189	141	190	142
rect	192	141	193	142
rect	195	141	196	142
rect	201	141	202	142
rect	204	141	205	142
rect	213	141	214	142
rect	216	141	217	142
rect	219	141	220	142
rect	222	141	223	142
rect	231	141	232	142
rect	243	141	244	142
rect	246	141	247	142
rect	249	141	250	142
rect	252	141	253	142
rect	264	141	265	142
rect	282	141	283	142
rect	285	141	286	142
rect	288	141	289	142
rect	294	141	295	142
rect	303	141	304	142
rect	306	141	307	142
rect	312	141	313	142
rect	315	141	316	142
rect	321	141	322	142
rect	324	141	325	142
rect	330	141	331	142
rect	333	141	334	142
rect	336	141	337	142
rect	339	141	340	142
rect	342	141	343	142
rect	351	141	352	142
rect	354	141	355	142
rect	357	141	358	142
rect	363	141	364	142
rect	366	141	367	142
rect	369	141	370	142
rect	375	141	376	142
rect	378	141	379	142
rect	387	141	388	142
rect	396	141	397	142
rect	402	141	403	142
rect	419	141	420	142
rect	21	142	22	143
rect	30	142	31	143
rect	36	142	37	143
rect	39	142	40	143
rect	42	142	43	143
rect	55	142	56	143
rect	58	142	59	143
rect	61	142	62	143
rect	70	142	71	143
rect	86	142	87	143
rect	89	142	90	143
rect	92	142	93	143
rect	112	142	113	143
rect	115	142	116	143
rect	118	142	119	143
rect	127	142	128	143
rect	130	142	131	143
rect	136	142	137	143
rect	149	142	150	143
rect	152	142	153	143
rect	155	142	156	143
rect	158	142	159	143
rect	174	142	175	143
rect	177	142	178	143
rect	183	142	184	143
rect	186	142	187	143
rect	189	142	190	143
rect	192	142	193	143
rect	195	142	196	143
rect	201	142	202	143
rect	204	142	205	143
rect	213	142	214	143
rect	216	142	217	143
rect	219	142	220	143
rect	222	142	223	143
rect	225	142	226	143
rect	231	142	232	143
rect	243	142	244	143
rect	246	142	247	143
rect	249	142	250	143
rect	252	142	253	143
rect	255	142	256	143
rect	264	142	265	143
rect	267	142	268	143
rect	276	142	277	143
rect	282	142	283	143
rect	285	142	286	143
rect	288	142	289	143
rect	291	142	292	143
rect	294	142	295	143
rect	303	142	304	143
rect	306	142	307	143
rect	312	142	313	143
rect	315	142	316	143
rect	321	142	322	143
rect	324	142	325	143
rect	327	142	328	143
rect	330	142	331	143
rect	333	142	334	143
rect	336	142	337	143
rect	339	142	340	143
rect	342	142	343	143
rect	351	142	352	143
rect	354	142	355	143
rect	357	142	358	143
rect	363	142	364	143
rect	366	142	367	143
rect	369	142	370	143
rect	375	142	376	143
rect	378	142	379	143
rect	387	142	388	143
rect	396	142	397	143
rect	402	142	403	143
rect	419	142	420	143
rect	21	143	22	144
rect	30	143	31	144
rect	36	143	37	144
rect	39	143	40	144
rect	42	143	43	144
rect	55	143	56	144
rect	58	143	59	144
rect	61	143	62	144
rect	70	143	71	144
rect	86	143	87	144
rect	89	143	90	144
rect	92	143	93	144
rect	112	143	113	144
rect	115	143	116	144
rect	118	143	119	144
rect	127	143	128	144
rect	130	143	131	144
rect	136	143	137	144
rect	149	143	150	144
rect	152	143	153	144
rect	155	143	156	144
rect	158	143	159	144
rect	174	143	175	144
rect	177	143	178	144
rect	183	143	184	144
rect	186	143	187	144
rect	192	143	193	144
rect	195	143	196	144
rect	201	143	202	144
rect	204	143	205	144
rect	213	143	214	144
rect	216	143	217	144
rect	219	143	220	144
rect	225	143	226	144
rect	231	143	232	144
rect	246	143	247	144
rect	249	143	250	144
rect	252	143	253	144
rect	255	143	256	144
rect	267	143	268	144
rect	276	143	277	144
rect	282	143	283	144
rect	288	143	289	144
rect	291	143	292	144
rect	294	143	295	144
rect	303	143	304	144
rect	306	143	307	144
rect	315	143	316	144
rect	321	143	322	144
rect	327	143	328	144
rect	330	143	331	144
rect	333	143	334	144
rect	336	143	337	144
rect	339	143	340	144
rect	342	143	343	144
rect	354	143	355	144
rect	357	143	358	144
rect	363	143	364	144
rect	366	143	367	144
rect	375	143	376	144
rect	378	143	379	144
rect	387	143	388	144
rect	396	143	397	144
rect	402	143	403	144
rect	419	143	420	144
rect	21	144	22	145
rect	30	144	31	145
rect	36	144	37	145
rect	39	144	40	145
rect	42	144	43	145
rect	55	144	56	145
rect	58	144	59	145
rect	61	144	62	145
rect	70	144	71	145
rect	86	144	87	145
rect	89	144	90	145
rect	92	144	93	145
rect	112	144	113	145
rect	115	144	116	145
rect	118	144	119	145
rect	127	144	128	145
rect	130	144	131	145
rect	136	144	137	145
rect	149	144	150	145
rect	152	144	153	145
rect	155	144	156	145
rect	158	144	159	145
rect	174	144	175	145
rect	177	144	178	145
rect	183	144	184	145
rect	186	144	187	145
rect	192	144	193	145
rect	195	144	196	145
rect	201	144	202	145
rect	204	144	205	145
rect	207	144	208	145
rect	213	144	214	145
rect	216	144	217	145
rect	219	144	220	145
rect	225	144	226	145
rect	231	144	232	145
rect	234	144	235	145
rect	246	144	247	145
rect	249	144	250	145
rect	252	144	253	145
rect	255	144	256	145
rect	261	144	262	145
rect	267	144	268	145
rect	276	144	277	145
rect	279	144	280	145
rect	282	144	283	145
rect	288	144	289	145
rect	291	144	292	145
rect	294	144	295	145
rect	297	144	298	145
rect	303	144	304	145
rect	306	144	307	145
rect	315	144	316	145
rect	321	144	322	145
rect	327	144	328	145
rect	330	144	331	145
rect	333	144	334	145
rect	336	144	337	145
rect	339	144	340	145
rect	342	144	343	145
rect	352	144	353	145
rect	354	144	355	145
rect	357	144	358	145
rect	363	144	364	145
rect	366	144	367	145
rect	375	144	376	145
rect	378	144	379	145
rect	382	144	383	145
rect	387	144	388	145
rect	396	144	397	145
rect	402	144	403	145
rect	419	144	420	145
rect	21	145	22	146
rect	30	145	31	146
rect	36	145	37	146
rect	39	145	40	146
rect	42	145	43	146
rect	55	145	56	146
rect	58	145	59	146
rect	61	145	62	146
rect	70	145	71	146
rect	86	145	87	146
rect	89	145	90	146
rect	112	145	113	146
rect	115	145	116	146
rect	118	145	119	146
rect	127	145	128	146
rect	130	145	131	146
rect	136	145	137	146
rect	149	145	150	146
rect	152	145	153	146
rect	155	145	156	146
rect	174	145	175	146
rect	177	145	178	146
rect	183	145	184	146
rect	186	145	187	146
rect	192	145	193	146
rect	195	145	196	146
rect	201	145	202	146
rect	204	145	205	146
rect	207	145	208	146
rect	213	145	214	146
rect	216	145	217	146
rect	219	145	220	146
rect	225	145	226	146
rect	231	145	232	146
rect	234	145	235	146
rect	246	145	247	146
rect	249	145	250	146
rect	252	145	253	146
rect	255	145	256	146
rect	261	145	262	146
rect	267	145	268	146
rect	276	145	277	146
rect	279	145	280	146
rect	282	145	283	146
rect	288	145	289	146
rect	291	145	292	146
rect	294	145	295	146
rect	297	145	298	146
rect	303	145	304	146
rect	306	145	307	146
rect	315	145	316	146
rect	321	145	322	146
rect	327	145	328	146
rect	330	145	331	146
rect	333	145	334	146
rect	336	145	337	146
rect	339	145	340	146
rect	342	145	343	146
rect	352	145	353	146
rect	354	145	355	146
rect	357	145	358	146
rect	363	145	364	146
rect	366	145	367	146
rect	375	145	376	146
rect	378	145	379	146
rect	382	145	383	146
rect	387	145	388	146
rect	396	145	397	146
rect	402	145	403	146
rect	419	145	420	146
rect	21	146	22	147
rect	30	146	31	147
rect	36	146	37	147
rect	39	146	40	147
rect	42	146	43	147
rect	55	146	56	147
rect	58	146	59	147
rect	61	146	62	147
rect	70	146	71	147
rect	86	146	87	147
rect	89	146	90	147
rect	98	146	99	147
rect	112	146	113	147
rect	115	146	116	147
rect	118	146	119	147
rect	127	146	128	147
rect	130	146	131	147
rect	136	146	137	147
rect	149	146	150	147
rect	152	146	153	147
rect	155	146	156	147
rect	167	146	168	147
rect	174	146	175	147
rect	177	146	178	147
rect	180	146	181	147
rect	183	146	184	147
rect	186	146	187	147
rect	192	146	193	147
rect	195	146	196	147
rect	201	146	202	147
rect	204	146	205	147
rect	207	146	208	147
rect	213	146	214	147
rect	216	146	217	147
rect	219	146	220	147
rect	225	146	226	147
rect	231	146	232	147
rect	234	146	235	147
rect	246	146	247	147
rect	249	146	250	147
rect	252	146	253	147
rect	255	146	256	147
rect	261	146	262	147
rect	267	146	268	147
rect	276	146	277	147
rect	279	146	280	147
rect	282	146	283	147
rect	288	146	289	147
rect	291	146	292	147
rect	294	146	295	147
rect	297	146	298	147
rect	303	146	304	147
rect	306	146	307	147
rect	315	146	316	147
rect	321	146	322	147
rect	327	146	328	147
rect	330	146	331	147
rect	333	146	334	147
rect	336	146	337	147
rect	339	146	340	147
rect	342	146	343	147
rect	352	146	353	147
rect	354	146	355	147
rect	357	146	358	147
rect	363	146	364	147
rect	366	146	367	147
rect	375	146	376	147
rect	378	146	379	147
rect	382	146	383	147
rect	387	146	388	147
rect	396	146	397	147
rect	402	146	403	147
rect	410	146	411	147
rect	419	146	420	147
rect	21	147	22	148
rect	30	147	31	148
rect	36	147	37	148
rect	39	147	40	148
rect	42	147	43	148
rect	55	147	56	148
rect	58	147	59	148
rect	61	147	62	148
rect	70	147	71	148
rect	86	147	87	148
rect	98	147	99	148
rect	112	147	113	148
rect	115	147	116	148
rect	118	147	119	148
rect	127	147	128	148
rect	130	147	131	148
rect	149	147	150	148
rect	152	147	153	148
rect	155	147	156	148
rect	167	147	168	148
rect	174	147	175	148
rect	177	147	178	148
rect	180	147	181	148
rect	183	147	184	148
rect	186	147	187	148
rect	192	147	193	148
rect	195	147	196	148
rect	201	147	202	148
rect	204	147	205	148
rect	207	147	208	148
rect	213	147	214	148
rect	216	147	217	148
rect	219	147	220	148
rect	225	147	226	148
rect	231	147	232	148
rect	234	147	235	148
rect	246	147	247	148
rect	249	147	250	148
rect	252	147	253	148
rect	255	147	256	148
rect	261	147	262	148
rect	267	147	268	148
rect	276	147	277	148
rect	279	147	280	148
rect	282	147	283	148
rect	288	147	289	148
rect	291	147	292	148
rect	294	147	295	148
rect	297	147	298	148
rect	303	147	304	148
rect	306	147	307	148
rect	315	147	316	148
rect	321	147	322	148
rect	327	147	328	148
rect	333	147	334	148
rect	336	147	337	148
rect	339	147	340	148
rect	342	147	343	148
rect	352	147	353	148
rect	354	147	355	148
rect	363	147	364	148
rect	375	147	376	148
rect	378	147	379	148
rect	382	147	383	148
rect	387	147	388	148
rect	396	147	397	148
rect	402	147	403	148
rect	410	147	411	148
rect	419	147	420	148
rect	21	148	22	149
rect	30	148	31	149
rect	36	148	37	149
rect	39	148	40	149
rect	42	148	43	149
rect	55	148	56	149
rect	58	148	59	149
rect	61	148	62	149
rect	70	148	71	149
rect	86	148	87	149
rect	95	148	96	149
rect	98	148	99	149
rect	112	148	113	149
rect	115	148	116	149
rect	118	148	119	149
rect	127	148	128	149
rect	130	148	131	149
rect	140	148	141	149
rect	149	148	150	149
rect	152	148	153	149
rect	155	148	156	149
rect	158	148	159	149
rect	167	148	168	149
rect	174	148	175	149
rect	177	148	178	149
rect	180	148	181	149
rect	183	148	184	149
rect	186	148	187	149
rect	192	148	193	149
rect	195	148	196	149
rect	201	148	202	149
rect	204	148	205	149
rect	207	148	208	149
rect	213	148	214	149
rect	216	148	217	149
rect	219	148	220	149
rect	225	148	226	149
rect	231	148	232	149
rect	234	148	235	149
rect	246	148	247	149
rect	249	148	250	149
rect	252	148	253	149
rect	255	148	256	149
rect	261	148	262	149
rect	267	148	268	149
rect	276	148	277	149
rect	279	148	280	149
rect	282	148	283	149
rect	288	148	289	149
rect	291	148	292	149
rect	294	148	295	149
rect	297	148	298	149
rect	300	148	301	149
rect	303	148	304	149
rect	306	148	307	149
rect	312	148	313	149
rect	315	148	316	149
rect	321	148	322	149
rect	327	148	328	149
rect	333	148	334	149
rect	336	148	337	149
rect	339	148	340	149
rect	342	148	343	149
rect	346	148	347	149
rect	352	148	353	149
rect	354	148	355	149
rect	363	148	364	149
rect	373	148	374	149
rect	375	148	376	149
rect	378	148	379	149
rect	382	148	383	149
rect	387	148	388	149
rect	396	148	397	149
rect	402	148	403	149
rect	410	148	411	149
rect	419	148	420	149
rect	21	149	22	150
rect	30	149	31	150
rect	36	149	37	150
rect	39	149	40	150
rect	55	149	56	150
rect	58	149	59	150
rect	61	149	62	150
rect	70	149	71	150
rect	95	149	96	150
rect	98	149	99	150
rect	112	149	113	150
rect	115	149	116	150
rect	130	149	131	150
rect	140	149	141	150
rect	149	149	150	150
rect	152	149	153	150
rect	158	149	159	150
rect	167	149	168	150
rect	174	149	175	150
rect	180	149	181	150
rect	183	149	184	150
rect	186	149	187	150
rect	195	149	196	150
rect	201	149	202	150
rect	204	149	205	150
rect	207	149	208	150
rect	216	149	217	150
rect	219	149	220	150
rect	225	149	226	150
rect	231	149	232	150
rect	234	149	235	150
rect	249	149	250	150
rect	255	149	256	150
rect	261	149	262	150
rect	267	149	268	150
rect	276	149	277	150
rect	279	149	280	150
rect	282	149	283	150
rect	288	149	289	150
rect	291	149	292	150
rect	297	149	298	150
rect	300	149	301	150
rect	303	149	304	150
rect	306	149	307	150
rect	312	149	313	150
rect	315	149	316	150
rect	321	149	322	150
rect	327	149	328	150
rect	336	149	337	150
rect	339	149	340	150
rect	346	149	347	150
rect	352	149	353	150
rect	363	149	364	150
rect	373	149	374	150
rect	375	149	376	150
rect	378	149	379	150
rect	382	149	383	150
rect	387	149	388	150
rect	396	149	397	150
rect	402	149	403	150
rect	410	149	411	150
rect	419	149	420	150
rect	21	150	22	151
rect	30	150	31	151
rect	36	150	37	151
rect	39	150	40	151
rect	47	150	48	151
rect	55	150	56	151
rect	58	150	59	151
rect	61	150	62	151
rect	70	150	71	151
rect	95	150	96	151
rect	98	150	99	151
rect	107	150	108	151
rect	112	150	113	151
rect	115	150	116	151
rect	119	150	120	151
rect	130	150	131	151
rect	137	150	138	151
rect	140	150	141	151
rect	149	150	150	151
rect	152	150	153	151
rect	158	150	159	151
rect	164	150	165	151
rect	167	150	168	151
rect	174	150	175	151
rect	180	150	181	151
rect	183	150	184	151
rect	186	150	187	151
rect	189	150	190	151
rect	195	150	196	151
rect	201	150	202	151
rect	204	150	205	151
rect	207	150	208	151
rect	210	150	211	151
rect	216	150	217	151
rect	219	150	220	151
rect	225	150	226	151
rect	228	150	229	151
rect	231	150	232	151
rect	234	150	235	151
rect	237	150	238	151
rect	249	150	250	151
rect	255	150	256	151
rect	261	150	262	151
rect	264	150	265	151
rect	267	150	268	151
rect	273	150	274	151
rect	276	150	277	151
rect	279	150	280	151
rect	282	150	283	151
rect	288	150	289	151
rect	291	150	292	151
rect	297	150	298	151
rect	300	150	301	151
rect	303	150	304	151
rect	306	150	307	151
rect	309	150	310	151
rect	312	150	313	151
rect	315	150	316	151
rect	321	150	322	151
rect	327	150	328	151
rect	336	150	337	151
rect	339	150	340	151
rect	346	150	347	151
rect	349	150	350	151
rect	352	150	353	151
rect	363	150	364	151
rect	370	150	371	151
rect	373	150	374	151
rect	375	150	376	151
rect	378	150	379	151
rect	382	150	383	151
rect	387	150	388	151
rect	396	150	397	151
rect	402	150	403	151
rect	410	150	411	151
rect	419	150	420	151
rect	21	151	22	152
rect	30	151	31	152
rect	39	151	40	152
rect	47	151	48	152
rect	55	151	56	152
rect	58	151	59	152
rect	61	151	62	152
rect	70	151	71	152
rect	95	151	96	152
rect	98	151	99	152
rect	107	151	108	152
rect	119	151	120	152
rect	137	151	138	152
rect	140	151	141	152
rect	149	151	150	152
rect	158	151	159	152
rect	164	151	165	152
rect	167	151	168	152
rect	180	151	181	152
rect	183	151	184	152
rect	186	151	187	152
rect	189	151	190	152
rect	201	151	202	152
rect	204	151	205	152
rect	207	151	208	152
rect	210	151	211	152
rect	216	151	217	152
rect	225	151	226	152
rect	228	151	229	152
rect	231	151	232	152
rect	234	151	235	152
rect	237	151	238	152
rect	255	151	256	152
rect	261	151	262	152
rect	264	151	265	152
rect	267	151	268	152
rect	273	151	274	152
rect	276	151	277	152
rect	279	151	280	152
rect	288	151	289	152
rect	291	151	292	152
rect	297	151	298	152
rect	300	151	301	152
rect	306	151	307	152
rect	309	151	310	152
rect	312	151	313	152
rect	315	151	316	152
rect	327	151	328	152
rect	336	151	337	152
rect	346	151	347	152
rect	349	151	350	152
rect	352	151	353	152
rect	363	151	364	152
rect	370	151	371	152
rect	373	151	374	152
rect	375	151	376	152
rect	378	151	379	152
rect	382	151	383	152
rect	387	151	388	152
rect	396	151	397	152
rect	402	151	403	152
rect	410	151	411	152
rect	419	151	420	152
rect	21	152	22	153
rect	30	152	31	153
rect	39	152	40	153
rect	47	152	48	153
rect	55	152	56	153
rect	58	152	59	153
rect	61	152	62	153
rect	70	152	71	153
rect	95	152	96	153
rect	98	152	99	153
rect	107	152	108	153
rect	116	152	117	153
rect	119	152	120	153
rect	128	152	129	153
rect	137	152	138	153
rect	140	152	141	153
rect	149	152	150	153
rect	158	152	159	153
rect	161	152	162	153
rect	164	152	165	153
rect	167	152	168	153
rect	180	152	181	153
rect	183	152	184	153
rect	186	152	187	153
rect	189	152	190	153
rect	192	152	193	153
rect	201	152	202	153
rect	204	152	205	153
rect	207	152	208	153
rect	210	152	211	153
rect	213	152	214	153
rect	216	152	217	153
rect	225	152	226	153
rect	228	152	229	153
rect	231	152	232	153
rect	234	152	235	153
rect	237	152	238	153
rect	246	152	247	153
rect	255	152	256	153
rect	258	152	259	153
rect	261	152	262	153
rect	264	152	265	153
rect	267	152	268	153
rect	273	152	274	153
rect	276	152	277	153
rect	279	152	280	153
rect	288	152	289	153
rect	291	152	292	153
rect	294	152	295	153
rect	297	152	298	153
rect	300	152	301	153
rect	306	152	307	153
rect	309	152	310	153
rect	312	152	313	153
rect	315	152	316	153
rect	318	152	319	153
rect	327	152	328	153
rect	330	152	331	153
rect	336	152	337	153
rect	346	152	347	153
rect	349	152	350	153
rect	352	152	353	153
rect	363	152	364	153
rect	367	152	368	153
rect	370	152	371	153
rect	373	152	374	153
rect	375	152	376	153
rect	378	152	379	153
rect	382	152	383	153
rect	387	152	388	153
rect	396	152	397	153
rect	402	152	403	153
rect	410	152	411	153
rect	419	152	420	153
rect	30	153	31	154
rect	39	153	40	154
rect	47	153	48	154
rect	61	153	62	154
rect	70	153	71	154
rect	95	153	96	154
rect	98	153	99	154
rect	107	153	108	154
rect	116	153	117	154
rect	119	153	120	154
rect	128	153	129	154
rect	137	153	138	154
rect	140	153	141	154
rect	149	153	150	154
rect	158	153	159	154
rect	161	153	162	154
rect	164	153	165	154
rect	167	153	168	154
rect	180	153	181	154
rect	183	153	184	154
rect	186	153	187	154
rect	189	153	190	154
rect	192	153	193	154
rect	201	153	202	154
rect	204	153	205	154
rect	207	153	208	154
rect	210	153	211	154
rect	213	153	214	154
rect	216	153	217	154
rect	225	153	226	154
rect	228	153	229	154
rect	231	153	232	154
rect	234	153	235	154
rect	237	153	238	154
rect	246	153	247	154
rect	255	153	256	154
rect	258	153	259	154
rect	261	153	262	154
rect	264	153	265	154
rect	267	153	268	154
rect	273	153	274	154
rect	276	153	277	154
rect	279	153	280	154
rect	288	153	289	154
rect	291	153	292	154
rect	294	153	295	154
rect	297	153	298	154
rect	300	153	301	154
rect	306	153	307	154
rect	309	153	310	154
rect	312	153	313	154
rect	315	153	316	154
rect	318	153	319	154
rect	327	153	328	154
rect	330	153	331	154
rect	336	153	337	154
rect	346	153	347	154
rect	349	153	350	154
rect	352	153	353	154
rect	363	153	364	154
rect	367	153	368	154
rect	370	153	371	154
rect	373	153	374	154
rect	375	153	376	154
rect	378	153	379	154
rect	382	153	383	154
rect	410	153	411	154
rect	419	153	420	154
rect	30	154	31	155
rect	39	154	40	155
rect	47	154	48	155
rect	61	154	62	155
rect	65	154	66	155
rect	70	154	71	155
rect	75	154	76	155
rect	95	154	96	155
rect	98	154	99	155
rect	107	154	108	155
rect	116	154	117	155
rect	119	154	120	155
rect	128	154	129	155
rect	137	154	138	155
rect	140	154	141	155
rect	149	154	150	155
rect	158	154	159	155
rect	161	154	162	155
rect	164	154	165	155
rect	167	154	168	155
rect	180	154	181	155
rect	183	154	184	155
rect	186	154	187	155
rect	189	154	190	155
rect	192	154	193	155
rect	201	154	202	155
rect	204	154	205	155
rect	207	154	208	155
rect	210	154	211	155
rect	213	154	214	155
rect	216	154	217	155
rect	225	154	226	155
rect	228	154	229	155
rect	231	154	232	155
rect	234	154	235	155
rect	237	154	238	155
rect	246	154	247	155
rect	255	154	256	155
rect	258	154	259	155
rect	261	154	262	155
rect	264	154	265	155
rect	267	154	268	155
rect	273	154	274	155
rect	276	154	277	155
rect	279	154	280	155
rect	288	154	289	155
rect	291	154	292	155
rect	294	154	295	155
rect	297	154	298	155
rect	300	154	301	155
rect	306	154	307	155
rect	309	154	310	155
rect	312	154	313	155
rect	315	154	316	155
rect	318	154	319	155
rect	327	154	328	155
rect	330	154	331	155
rect	336	154	337	155
rect	346	154	347	155
rect	349	154	350	155
rect	352	154	353	155
rect	358	154	359	155
rect	363	154	364	155
rect	367	154	368	155
rect	370	154	371	155
rect	373	154	374	155
rect	375	154	376	155
rect	378	154	379	155
rect	382	154	383	155
rect	391	154	392	155
rect	410	154	411	155
rect	419	154	420	155
rect	47	155	48	156
rect	65	155	66	156
rect	75	155	76	156
rect	95	155	96	156
rect	98	155	99	156
rect	107	155	108	156
rect	116	155	117	156
rect	119	155	120	156
rect	128	155	129	156
rect	137	155	138	156
rect	140	155	141	156
rect	149	155	150	156
rect	158	155	159	156
rect	161	155	162	156
rect	164	155	165	156
rect	167	155	168	156
rect	180	155	181	156
rect	183	155	184	156
rect	186	155	187	156
rect	189	155	190	156
rect	192	155	193	156
rect	201	155	202	156
rect	204	155	205	156
rect	207	155	208	156
rect	210	155	211	156
rect	213	155	214	156
rect	216	155	217	156
rect	225	155	226	156
rect	228	155	229	156
rect	231	155	232	156
rect	234	155	235	156
rect	237	155	238	156
rect	246	155	247	156
rect	255	155	256	156
rect	258	155	259	156
rect	261	155	262	156
rect	264	155	265	156
rect	267	155	268	156
rect	273	155	274	156
rect	276	155	277	156
rect	279	155	280	156
rect	288	155	289	156
rect	291	155	292	156
rect	294	155	295	156
rect	297	155	298	156
rect	300	155	301	156
rect	306	155	307	156
rect	309	155	310	156
rect	312	155	313	156
rect	315	155	316	156
rect	318	155	319	156
rect	327	155	328	156
rect	330	155	331	156
rect	346	155	347	156
rect	349	155	350	156
rect	352	155	353	156
rect	358	155	359	156
rect	367	155	368	156
rect	370	155	371	156
rect	373	155	374	156
rect	382	155	383	156
rect	391	155	392	156
rect	410	155	411	156
rect	35	156	36	157
rect	44	156	45	157
rect	47	156	48	157
rect	56	156	57	157
rect	65	156	66	157
rect	75	156	76	157
rect	95	156	96	157
rect	98	156	99	157
rect	107	156	108	157
rect	116	156	117	157
rect	119	156	120	157
rect	128	156	129	157
rect	137	156	138	157
rect	140	156	141	157
rect	149	156	150	157
rect	158	156	159	157
rect	161	156	162	157
rect	164	156	165	157
rect	167	156	168	157
rect	180	156	181	157
rect	183	156	184	157
rect	186	156	187	157
rect	189	156	190	157
rect	192	156	193	157
rect	201	156	202	157
rect	204	156	205	157
rect	207	156	208	157
rect	210	156	211	157
rect	213	156	214	157
rect	216	156	217	157
rect	225	156	226	157
rect	228	156	229	157
rect	231	156	232	157
rect	234	156	235	157
rect	237	156	238	157
rect	246	156	247	157
rect	255	156	256	157
rect	258	156	259	157
rect	261	156	262	157
rect	264	156	265	157
rect	267	156	268	157
rect	273	156	274	157
rect	276	156	277	157
rect	279	156	280	157
rect	288	156	289	157
rect	291	156	292	157
rect	294	156	295	157
rect	297	156	298	157
rect	300	156	301	157
rect	306	156	307	157
rect	309	156	310	157
rect	312	156	313	157
rect	315	156	316	157
rect	318	156	319	157
rect	324	156	325	157
rect	327	156	328	157
rect	330	156	331	157
rect	346	156	347	157
rect	349	156	350	157
rect	352	156	353	157
rect	355	156	356	157
rect	358	156	359	157
rect	367	156	368	157
rect	370	156	371	157
rect	373	156	374	157
rect	382	156	383	157
rect	391	156	392	157
rect	394	156	395	157
rect	410	156	411	157
rect	413	156	414	157
rect	8	163	9	164
rect	29	163	30	164
rect	35	163	36	164
rect	44	163	45	164
rect	47	163	48	164
rect	50	163	51	164
rect	56	163	57	164
rect	65	163	66	164
rect	95	163	96	164
rect	98	163	99	164
rect	107	163	108	164
rect	116	163	117	164
rect	119	163	120	164
rect	128	163	129	164
rect	137	163	138	164
rect	140	163	141	164
rect	149	163	150	164
rect	158	163	159	164
rect	161	163	162	164
rect	164	163	165	164
rect	167	163	168	164
rect	173	163	174	164
rect	177	163	178	164
rect	183	163	184	164
rect	186	163	187	164
rect	189	163	190	164
rect	192	163	193	164
rect	201	163	202	164
rect	204	163	205	164
rect	207	163	208	164
rect	210	163	211	164
rect	213	163	214	164
rect	216	163	217	164
rect	219	163	220	164
rect	225	163	226	164
rect	228	163	229	164
rect	231	163	232	164
rect	234	163	235	164
rect	237	163	238	164
rect	240	163	241	164
rect	246	163	247	164
rect	255	163	256	164
rect	258	163	259	164
rect	261	163	262	164
rect	264	163	265	164
rect	273	163	274	164
rect	276	163	277	164
rect	279	163	280	164
rect	288	163	289	164
rect	291	163	292	164
rect	294	163	295	164
rect	297	163	298	164
rect	303	163	304	164
rect	306	163	307	164
rect	309	163	310	164
rect	312	163	313	164
rect	315	163	316	164
rect	318	163	319	164
rect	321	163	322	164
rect	327	163	328	164
rect	330	163	331	164
rect	346	163	347	164
rect	349	163	350	164
rect	358	163	359	164
rect	367	163	368	164
rect	370	163	371	164
rect	373	163	374	164
rect	382	163	383	164
rect	388	163	389	164
rect	391	163	392	164
rect	394	163	395	164
rect	410	163	411	164
rect	413	163	414	164
rect	8	164	9	165
rect	29	164	30	165
rect	35	164	36	165
rect	44	164	45	165
rect	47	164	48	165
rect	50	164	51	165
rect	56	164	57	165
rect	65	164	66	165
rect	95	164	96	165
rect	98	164	99	165
rect	107	164	108	165
rect	116	164	117	165
rect	119	164	120	165
rect	128	164	129	165
rect	137	164	138	165
rect	140	164	141	165
rect	149	164	150	165
rect	158	164	159	165
rect	161	164	162	165
rect	164	164	165	165
rect	167	164	168	165
rect	173	164	174	165
rect	177	164	178	165
rect	183	164	184	165
rect	186	164	187	165
rect	189	164	190	165
rect	192	164	193	165
rect	201	164	202	165
rect	204	164	205	165
rect	207	164	208	165
rect	210	164	211	165
rect	213	164	214	165
rect	216	164	217	165
rect	219	164	220	165
rect	225	164	226	165
rect	228	164	229	165
rect	231	164	232	165
rect	234	164	235	165
rect	237	164	238	165
rect	240	164	241	165
rect	246	164	247	165
rect	255	164	256	165
rect	258	164	259	165
rect	261	164	262	165
rect	264	164	265	165
rect	279	164	280	165
rect	288	164	289	165
rect	291	164	292	165
rect	294	164	295	165
rect	297	164	298	165
rect	303	164	304	165
rect	306	164	307	165
rect	309	164	310	165
rect	312	164	313	165
rect	315	164	316	165
rect	318	164	319	165
rect	321	164	322	165
rect	327	164	328	165
rect	346	164	347	165
rect	349	164	350	165
rect	358	164	359	165
rect	367	164	368	165
rect	370	164	371	165
rect	373	164	374	165
rect	382	164	383	165
rect	388	164	389	165
rect	391	164	392	165
rect	394	164	395	165
rect	410	164	411	165
rect	413	164	414	165
rect	8	165	9	166
rect	29	165	30	166
rect	35	165	36	166
rect	44	165	45	166
rect	47	165	48	166
rect	50	165	51	166
rect	56	165	57	166
rect	65	165	66	166
rect	95	165	96	166
rect	98	165	99	166
rect	107	165	108	166
rect	116	165	117	166
rect	119	165	120	166
rect	128	165	129	166
rect	137	165	138	166
rect	140	165	141	166
rect	149	165	150	166
rect	158	165	159	166
rect	161	165	162	166
rect	164	165	165	166
rect	167	165	168	166
rect	173	165	174	166
rect	177	165	178	166
rect	183	165	184	166
rect	186	165	187	166
rect	189	165	190	166
rect	192	165	193	166
rect	201	165	202	166
rect	204	165	205	166
rect	207	165	208	166
rect	210	165	211	166
rect	213	165	214	166
rect	216	165	217	166
rect	219	165	220	166
rect	225	165	226	166
rect	228	165	229	166
rect	231	165	232	166
rect	234	165	235	166
rect	237	165	238	166
rect	240	165	241	166
rect	246	165	247	166
rect	248	165	249	166
rect	255	165	256	166
rect	258	165	259	166
rect	261	165	262	166
rect	264	165	265	166
rect	279	165	280	166
rect	281	165	282	166
rect	288	165	289	166
rect	291	165	292	166
rect	294	165	295	166
rect	297	165	298	166
rect	303	165	304	166
rect	306	165	307	166
rect	309	165	310	166
rect	312	165	313	166
rect	315	165	316	166
rect	318	165	319	166
rect	321	165	322	166
rect	327	165	328	166
rect	332	165	333	166
rect	346	165	347	166
rect	349	165	350	166
rect	358	165	359	166
rect	367	165	368	166
rect	370	165	371	166
rect	373	165	374	166
rect	382	165	383	166
rect	388	165	389	166
rect	391	165	392	166
rect	394	165	395	166
rect	410	165	411	166
rect	413	165	414	166
rect	8	166	9	167
rect	29	166	30	167
rect	35	166	36	167
rect	44	166	45	167
rect	47	166	48	167
rect	50	166	51	167
rect	56	166	57	167
rect	65	166	66	167
rect	95	166	96	167
rect	98	166	99	167
rect	107	166	108	167
rect	116	166	117	167
rect	119	166	120	167
rect	128	166	129	167
rect	137	166	138	167
rect	140	166	141	167
rect	149	166	150	167
rect	158	166	159	167
rect	161	166	162	167
rect	164	166	165	167
rect	167	166	168	167
rect	173	166	174	167
rect	177	166	178	167
rect	183	166	184	167
rect	186	166	187	167
rect	189	166	190	167
rect	192	166	193	167
rect	201	166	202	167
rect	204	166	205	167
rect	207	166	208	167
rect	210	166	211	167
rect	213	166	214	167
rect	216	166	217	167
rect	219	166	220	167
rect	225	166	226	167
rect	228	166	229	167
rect	231	166	232	167
rect	234	166	235	167
rect	237	166	238	167
rect	240	166	241	167
rect	248	166	249	167
rect	255	166	256	167
rect	258	166	259	167
rect	261	166	262	167
rect	264	166	265	167
rect	279	166	280	167
rect	281	166	282	167
rect	288	166	289	167
rect	291	166	292	167
rect	294	166	295	167
rect	297	166	298	167
rect	303	166	304	167
rect	306	166	307	167
rect	312	166	313	167
rect	315	166	316	167
rect	321	166	322	167
rect	327	166	328	167
rect	332	166	333	167
rect	346	166	347	167
rect	349	166	350	167
rect	358	166	359	167
rect	367	166	368	167
rect	370	166	371	167
rect	373	166	374	167
rect	382	166	383	167
rect	388	166	389	167
rect	391	166	392	167
rect	394	166	395	167
rect	410	166	411	167
rect	413	166	414	167
rect	8	167	9	168
rect	29	167	30	168
rect	35	167	36	168
rect	44	167	45	168
rect	47	167	48	168
rect	50	167	51	168
rect	56	167	57	168
rect	65	167	66	168
rect	95	167	96	168
rect	98	167	99	168
rect	107	167	108	168
rect	116	167	117	168
rect	119	167	120	168
rect	128	167	129	168
rect	137	167	138	168
rect	140	167	141	168
rect	149	167	150	168
rect	158	167	159	168
rect	161	167	162	168
rect	164	167	165	168
rect	167	167	168	168
rect	173	167	174	168
rect	177	167	178	168
rect	183	167	184	168
rect	186	167	187	168
rect	189	167	190	168
rect	192	167	193	168
rect	201	167	202	168
rect	204	167	205	168
rect	207	167	208	168
rect	210	167	211	168
rect	213	167	214	168
rect	216	167	217	168
rect	219	167	220	168
rect	225	167	226	168
rect	228	167	229	168
rect	231	167	232	168
rect	234	167	235	168
rect	237	167	238	168
rect	240	167	241	168
rect	242	167	243	168
rect	248	167	249	168
rect	255	167	256	168
rect	258	167	259	168
rect	261	167	262	168
rect	264	167	265	168
rect	275	167	276	168
rect	279	167	280	168
rect	281	167	282	168
rect	288	167	289	168
rect	291	167	292	168
rect	294	167	295	168
rect	297	167	298	168
rect	303	167	304	168
rect	306	167	307	168
rect	312	167	313	168
rect	315	167	316	168
rect	321	167	322	168
rect	327	167	328	168
rect	329	167	330	168
rect	332	167	333	168
rect	346	167	347	168
rect	349	167	350	168
rect	358	167	359	168
rect	367	167	368	168
rect	370	167	371	168
rect	373	167	374	168
rect	382	167	383	168
rect	388	167	389	168
rect	391	167	392	168
rect	394	167	395	168
rect	410	167	411	168
rect	413	167	414	168
rect	8	168	9	169
rect	29	168	30	169
rect	35	168	36	169
rect	44	168	45	169
rect	47	168	48	169
rect	50	168	51	169
rect	56	168	57	169
rect	65	168	66	169
rect	95	168	96	169
rect	98	168	99	169
rect	107	168	108	169
rect	116	168	117	169
rect	119	168	120	169
rect	128	168	129	169
rect	137	168	138	169
rect	140	168	141	169
rect	149	168	150	169
rect	158	168	159	169
rect	161	168	162	169
rect	164	168	165	169
rect	167	168	168	169
rect	173	168	174	169
rect	177	168	178	169
rect	183	168	184	169
rect	186	168	187	169
rect	189	168	190	169
rect	192	168	193	169
rect	201	168	202	169
rect	204	168	205	169
rect	207	168	208	169
rect	210	168	211	169
rect	213	168	214	169
rect	216	168	217	169
rect	219	168	220	169
rect	225	168	226	169
rect	228	168	229	169
rect	231	168	232	169
rect	234	168	235	169
rect	237	168	238	169
rect	240	168	241	169
rect	242	168	243	169
rect	248	168	249	169
rect	258	168	259	169
rect	261	168	262	169
rect	264	168	265	169
rect	275	168	276	169
rect	281	168	282	169
rect	288	168	289	169
rect	291	168	292	169
rect	294	168	295	169
rect	297	168	298	169
rect	303	168	304	169
rect	312	168	313	169
rect	315	168	316	169
rect	327	168	328	169
rect	329	168	330	169
rect	332	168	333	169
rect	346	168	347	169
rect	349	168	350	169
rect	358	168	359	169
rect	367	168	368	169
rect	370	168	371	169
rect	373	168	374	169
rect	382	168	383	169
rect	388	168	389	169
rect	391	168	392	169
rect	394	168	395	169
rect	410	168	411	169
rect	413	168	414	169
rect	8	169	9	170
rect	29	169	30	170
rect	35	169	36	170
rect	44	169	45	170
rect	47	169	48	170
rect	50	169	51	170
rect	56	169	57	170
rect	65	169	66	170
rect	95	169	96	170
rect	98	169	99	170
rect	107	169	108	170
rect	116	169	117	170
rect	119	169	120	170
rect	128	169	129	170
rect	137	169	138	170
rect	140	169	141	170
rect	149	169	150	170
rect	158	169	159	170
rect	161	169	162	170
rect	164	169	165	170
rect	167	169	168	170
rect	173	169	174	170
rect	177	169	178	170
rect	183	169	184	170
rect	186	169	187	170
rect	189	169	190	170
rect	192	169	193	170
rect	201	169	202	170
rect	204	169	205	170
rect	207	169	208	170
rect	210	169	211	170
rect	213	169	214	170
rect	216	169	217	170
rect	219	169	220	170
rect	225	169	226	170
rect	228	169	229	170
rect	231	169	232	170
rect	234	169	235	170
rect	237	169	238	170
rect	240	169	241	170
rect	242	169	243	170
rect	245	169	246	170
rect	248	169	249	170
rect	258	169	259	170
rect	261	169	262	170
rect	264	169	265	170
rect	269	169	270	170
rect	275	169	276	170
rect	281	169	282	170
rect	288	169	289	170
rect	291	169	292	170
rect	294	169	295	170
rect	297	169	298	170
rect	303	169	304	170
rect	312	169	313	170
rect	315	169	316	170
rect	327	169	328	170
rect	329	169	330	170
rect	332	169	333	170
rect	346	169	347	170
rect	349	169	350	170
rect	358	169	359	170
rect	367	169	368	170
rect	370	169	371	170
rect	373	169	374	170
rect	382	169	383	170
rect	388	169	389	170
rect	391	169	392	170
rect	394	169	395	170
rect	410	169	411	170
rect	413	169	414	170
rect	8	170	9	171
rect	29	170	30	171
rect	35	170	36	171
rect	44	170	45	171
rect	47	170	48	171
rect	50	170	51	171
rect	56	170	57	171
rect	65	170	66	171
rect	95	170	96	171
rect	98	170	99	171
rect	107	170	108	171
rect	116	170	117	171
rect	119	170	120	171
rect	128	170	129	171
rect	137	170	138	171
rect	140	170	141	171
rect	149	170	150	171
rect	158	170	159	171
rect	161	170	162	171
rect	164	170	165	171
rect	167	170	168	171
rect	173	170	174	171
rect	177	170	178	171
rect	183	170	184	171
rect	186	170	187	171
rect	189	170	190	171
rect	192	170	193	171
rect	201	170	202	171
rect	204	170	205	171
rect	207	170	208	171
rect	210	170	211	171
rect	213	170	214	171
rect	216	170	217	171
rect	219	170	220	171
rect	225	170	226	171
rect	228	170	229	171
rect	234	170	235	171
rect	237	170	238	171
rect	240	170	241	171
rect	242	170	243	171
rect	245	170	246	171
rect	248	170	249	171
rect	258	170	259	171
rect	261	170	262	171
rect	269	170	270	171
rect	275	170	276	171
rect	281	170	282	171
rect	288	170	289	171
rect	291	170	292	171
rect	294	170	295	171
rect	303	170	304	171
rect	312	170	313	171
rect	327	170	328	171
rect	329	170	330	171
rect	332	170	333	171
rect	346	170	347	171
rect	349	170	350	171
rect	358	170	359	171
rect	367	170	368	171
rect	370	170	371	171
rect	373	170	374	171
rect	382	170	383	171
rect	388	170	389	171
rect	391	170	392	171
rect	394	170	395	171
rect	410	170	411	171
rect	413	170	414	171
rect	8	171	9	172
rect	29	171	30	172
rect	35	171	36	172
rect	44	171	45	172
rect	47	171	48	172
rect	50	171	51	172
rect	56	171	57	172
rect	65	171	66	172
rect	95	171	96	172
rect	98	171	99	172
rect	107	171	108	172
rect	116	171	117	172
rect	119	171	120	172
rect	128	171	129	172
rect	137	171	138	172
rect	140	171	141	172
rect	149	171	150	172
rect	158	171	159	172
rect	161	171	162	172
rect	164	171	165	172
rect	167	171	168	172
rect	173	171	174	172
rect	177	171	178	172
rect	183	171	184	172
rect	186	171	187	172
rect	189	171	190	172
rect	192	171	193	172
rect	201	171	202	172
rect	204	171	205	172
rect	207	171	208	172
rect	210	171	211	172
rect	213	171	214	172
rect	216	171	217	172
rect	219	171	220	172
rect	225	171	226	172
rect	228	171	229	172
rect	234	171	235	172
rect	237	171	238	172
rect	240	171	241	172
rect	242	171	243	172
rect	245	171	246	172
rect	248	171	249	172
rect	251	171	252	172
rect	258	171	259	172
rect	261	171	262	172
rect	269	171	270	172
rect	275	171	276	172
rect	278	171	279	172
rect	281	171	282	172
rect	288	171	289	172
rect	291	171	292	172
rect	294	171	295	172
rect	303	171	304	172
rect	305	171	306	172
rect	312	171	313	172
rect	317	171	318	172
rect	327	171	328	172
rect	329	171	330	172
rect	332	171	333	172
rect	346	171	347	172
rect	349	171	350	172
rect	358	171	359	172
rect	367	171	368	172
rect	370	171	371	172
rect	373	171	374	172
rect	382	171	383	172
rect	388	171	389	172
rect	391	171	392	172
rect	394	171	395	172
rect	410	171	411	172
rect	413	171	414	172
rect	8	172	9	173
rect	29	172	30	173
rect	35	172	36	173
rect	44	172	45	173
rect	47	172	48	173
rect	50	172	51	173
rect	56	172	57	173
rect	65	172	66	173
rect	95	172	96	173
rect	98	172	99	173
rect	107	172	108	173
rect	116	172	117	173
rect	119	172	120	173
rect	128	172	129	173
rect	137	172	138	173
rect	140	172	141	173
rect	149	172	150	173
rect	158	172	159	173
rect	161	172	162	173
rect	164	172	165	173
rect	167	172	168	173
rect	173	172	174	173
rect	177	172	178	173
rect	183	172	184	173
rect	186	172	187	173
rect	189	172	190	173
rect	192	172	193	173
rect	201	172	202	173
rect	204	172	205	173
rect	210	172	211	173
rect	213	172	214	173
rect	216	172	217	173
rect	219	172	220	173
rect	225	172	226	173
rect	228	172	229	173
rect	237	172	238	173
rect	240	172	241	173
rect	242	172	243	173
rect	245	172	246	173
rect	248	172	249	173
rect	251	172	252	173
rect	261	172	262	173
rect	269	172	270	173
rect	275	172	276	173
rect	278	172	279	173
rect	281	172	282	173
rect	288	172	289	173
rect	291	172	292	173
rect	294	172	295	173
rect	303	172	304	173
rect	305	172	306	173
rect	312	172	313	173
rect	317	172	318	173
rect	327	172	328	173
rect	329	172	330	173
rect	332	172	333	173
rect	346	172	347	173
rect	349	172	350	173
rect	358	172	359	173
rect	367	172	368	173
rect	370	172	371	173
rect	382	172	383	173
rect	388	172	389	173
rect	391	172	392	173
rect	394	172	395	173
rect	410	172	411	173
rect	413	172	414	173
rect	8	173	9	174
rect	29	173	30	174
rect	35	173	36	174
rect	44	173	45	174
rect	47	173	48	174
rect	50	173	51	174
rect	56	173	57	174
rect	65	173	66	174
rect	95	173	96	174
rect	98	173	99	174
rect	107	173	108	174
rect	116	173	117	174
rect	119	173	120	174
rect	128	173	129	174
rect	137	173	138	174
rect	140	173	141	174
rect	149	173	150	174
rect	158	173	159	174
rect	161	173	162	174
rect	164	173	165	174
rect	167	173	168	174
rect	173	173	174	174
rect	177	173	178	174
rect	183	173	184	174
rect	186	173	187	174
rect	189	173	190	174
rect	192	173	193	174
rect	201	173	202	174
rect	204	173	205	174
rect	210	173	211	174
rect	213	173	214	174
rect	216	173	217	174
rect	219	173	220	174
rect	225	173	226	174
rect	228	173	229	174
rect	230	173	231	174
rect	237	173	238	174
rect	240	173	241	174
rect	242	173	243	174
rect	245	173	246	174
rect	248	173	249	174
rect	251	173	252	174
rect	254	173	255	174
rect	261	173	262	174
rect	266	173	267	174
rect	269	173	270	174
rect	272	173	273	174
rect	275	173	276	174
rect	278	173	279	174
rect	281	173	282	174
rect	288	173	289	174
rect	291	173	292	174
rect	294	173	295	174
rect	303	173	304	174
rect	305	173	306	174
rect	312	173	313	174
rect	317	173	318	174
rect	327	173	328	174
rect	329	173	330	174
rect	332	173	333	174
rect	346	173	347	174
rect	349	173	350	174
rect	358	173	359	174
rect	367	173	368	174
rect	370	173	371	174
rect	382	173	383	174
rect	388	173	389	174
rect	391	173	392	174
rect	394	173	395	174
rect	410	173	411	174
rect	413	173	414	174
rect	8	174	9	175
rect	29	174	30	175
rect	35	174	36	175
rect	44	174	45	175
rect	47	174	48	175
rect	56	174	57	175
rect	65	174	66	175
rect	95	174	96	175
rect	98	174	99	175
rect	107	174	108	175
rect	116	174	117	175
rect	119	174	120	175
rect	128	174	129	175
rect	137	174	138	175
rect	140	174	141	175
rect	149	174	150	175
rect	158	174	159	175
rect	161	174	162	175
rect	164	174	165	175
rect	167	174	168	175
rect	173	174	174	175
rect	177	174	178	175
rect	183	174	184	175
rect	186	174	187	175
rect	189	174	190	175
rect	192	174	193	175
rect	201	174	202	175
rect	204	174	205	175
rect	210	174	211	175
rect	213	174	214	175
rect	216	174	217	175
rect	219	174	220	175
rect	225	174	226	175
rect	228	174	229	175
rect	230	174	231	175
rect	237	174	238	175
rect	240	174	241	175
rect	242	174	243	175
rect	245	174	246	175
rect	248	174	249	175
rect	251	174	252	175
rect	254	174	255	175
rect	261	174	262	175
rect	266	174	267	175
rect	269	174	270	175
rect	272	174	273	175
rect	275	174	276	175
rect	278	174	279	175
rect	281	174	282	175
rect	288	174	289	175
rect	303	174	304	175
rect	305	174	306	175
rect	312	174	313	175
rect	317	174	318	175
rect	327	174	328	175
rect	329	174	330	175
rect	332	174	333	175
rect	346	174	347	175
rect	349	174	350	175
rect	358	174	359	175
rect	367	174	368	175
rect	370	174	371	175
rect	382	174	383	175
rect	388	174	389	175
rect	391	174	392	175
rect	394	174	395	175
rect	410	174	411	175
rect	413	174	414	175
rect	8	175	9	176
rect	29	175	30	176
rect	35	175	36	176
rect	44	175	45	176
rect	47	175	48	176
rect	56	175	57	176
rect	65	175	66	176
rect	95	175	96	176
rect	98	175	99	176
rect	107	175	108	176
rect	116	175	117	176
rect	119	175	120	176
rect	128	175	129	176
rect	137	175	138	176
rect	140	175	141	176
rect	149	175	150	176
rect	158	175	159	176
rect	161	175	162	176
rect	164	175	165	176
rect	167	175	168	176
rect	173	175	174	176
rect	177	175	178	176
rect	183	175	184	176
rect	186	175	187	176
rect	189	175	190	176
rect	192	175	193	176
rect	201	175	202	176
rect	204	175	205	176
rect	210	175	211	176
rect	213	175	214	176
rect	216	175	217	176
rect	219	175	220	176
rect	225	175	226	176
rect	228	175	229	176
rect	230	175	231	176
rect	237	175	238	176
rect	240	175	241	176
rect	242	175	243	176
rect	245	175	246	176
rect	248	175	249	176
rect	251	175	252	176
rect	254	175	255	176
rect	261	175	262	176
rect	266	175	267	176
rect	269	175	270	176
rect	272	175	273	176
rect	275	175	276	176
rect	278	175	279	176
rect	281	175	282	176
rect	288	175	289	176
rect	303	175	304	176
rect	305	175	306	176
rect	312	175	313	176
rect	314	175	315	176
rect	317	175	318	176
rect	327	175	328	176
rect	329	175	330	176
rect	332	175	333	176
rect	346	175	347	176
rect	349	175	350	176
rect	358	175	359	176
rect	367	175	368	176
rect	370	175	371	176
rect	382	175	383	176
rect	388	175	389	176
rect	391	175	392	176
rect	394	175	395	176
rect	410	175	411	176
rect	413	175	414	176
rect	8	176	9	177
rect	29	176	30	177
rect	35	176	36	177
rect	44	176	45	177
rect	47	176	48	177
rect	56	176	57	177
rect	65	176	66	177
rect	95	176	96	177
rect	98	176	99	177
rect	107	176	108	177
rect	116	176	117	177
rect	119	176	120	177
rect	128	176	129	177
rect	137	176	138	177
rect	140	176	141	177
rect	158	176	159	177
rect	161	176	162	177
rect	164	176	165	177
rect	167	176	168	177
rect	173	176	174	177
rect	177	176	178	177
rect	183	176	184	177
rect	186	176	187	177
rect	189	176	190	177
rect	201	176	202	177
rect	204	176	205	177
rect	210	176	211	177
rect	213	176	214	177
rect	216	176	217	177
rect	225	176	226	177
rect	228	176	229	177
rect	230	176	231	177
rect	237	176	238	177
rect	240	176	241	177
rect	242	176	243	177
rect	245	176	246	177
rect	248	176	249	177
rect	251	176	252	177
rect	254	176	255	177
rect	261	176	262	177
rect	266	176	267	177
rect	269	176	270	177
rect	272	176	273	177
rect	275	176	276	177
rect	278	176	279	177
rect	281	176	282	177
rect	288	176	289	177
rect	303	176	304	177
rect	305	176	306	177
rect	314	176	315	177
rect	317	176	318	177
rect	327	176	328	177
rect	329	176	330	177
rect	332	176	333	177
rect	346	176	347	177
rect	349	176	350	177
rect	358	176	359	177
rect	370	176	371	177
rect	382	176	383	177
rect	388	176	389	177
rect	391	176	392	177
rect	394	176	395	177
rect	410	176	411	177
rect	413	176	414	177
rect	8	177	9	178
rect	29	177	30	178
rect	35	177	36	178
rect	44	177	45	178
rect	47	177	48	178
rect	56	177	57	178
rect	65	177	66	178
rect	95	177	96	178
rect	98	177	99	178
rect	107	177	108	178
rect	116	177	117	178
rect	119	177	120	178
rect	128	177	129	178
rect	137	177	138	178
rect	140	177	141	178
rect	152	177	153	178
rect	158	177	159	178
rect	161	177	162	178
rect	164	177	165	178
rect	167	177	168	178
rect	173	177	174	178
rect	177	177	178	178
rect	183	177	184	178
rect	186	177	187	178
rect	189	177	190	178
rect	201	177	202	178
rect	204	177	205	178
rect	208	177	209	178
rect	210	177	211	178
rect	213	177	214	178
rect	216	177	217	178
rect	225	177	226	178
rect	228	177	229	178
rect	230	177	231	178
rect	237	177	238	178
rect	240	177	241	178
rect	242	177	243	178
rect	245	177	246	178
rect	248	177	249	178
rect	251	177	252	178
rect	254	177	255	178
rect	261	177	262	178
rect	266	177	267	178
rect	269	177	270	178
rect	272	177	273	178
rect	275	177	276	178
rect	278	177	279	178
rect	281	177	282	178
rect	288	177	289	178
rect	290	177	291	178
rect	293	177	294	178
rect	303	177	304	178
rect	305	177	306	178
rect	314	177	315	178
rect	317	177	318	178
rect	327	177	328	178
rect	329	177	330	178
rect	332	177	333	178
rect	346	177	347	178
rect	349	177	350	178
rect	353	177	354	178
rect	358	177	359	178
rect	370	177	371	178
rect	382	177	383	178
rect	388	177	389	178
rect	391	177	392	178
rect	394	177	395	178
rect	410	177	411	178
rect	413	177	414	178
rect	8	178	9	179
rect	29	178	30	179
rect	35	178	36	179
rect	44	178	45	179
rect	47	178	48	179
rect	56	178	57	179
rect	65	178	66	179
rect	95	178	96	179
rect	98	178	99	179
rect	107	178	108	179
rect	116	178	117	179
rect	119	178	120	179
rect	128	178	129	179
rect	140	178	141	179
rect	152	178	153	179
rect	158	178	159	179
rect	161	178	162	179
rect	164	178	165	179
rect	167	178	168	179
rect	173	178	174	179
rect	186	178	187	179
rect	189	178	190	179
rect	208	178	209	179
rect	210	178	211	179
rect	216	178	217	179
rect	225	178	226	179
rect	228	178	229	179
rect	230	178	231	179
rect	240	178	241	179
rect	242	178	243	179
rect	245	178	246	179
rect	248	178	249	179
rect	251	178	252	179
rect	254	178	255	179
rect	261	178	262	179
rect	266	178	267	179
rect	269	178	270	179
rect	272	178	273	179
rect	275	178	276	179
rect	278	178	279	179
rect	281	178	282	179
rect	288	178	289	179
rect	290	178	291	179
rect	293	178	294	179
rect	303	178	304	179
rect	305	178	306	179
rect	314	178	315	179
rect	317	178	318	179
rect	329	178	330	179
rect	332	178	333	179
rect	346	178	347	179
rect	353	178	354	179
rect	370	178	371	179
rect	388	178	389	179
rect	391	178	392	179
rect	394	178	395	179
rect	410	178	411	179
rect	413	178	414	179
rect	8	179	9	180
rect	29	179	30	180
rect	35	179	36	180
rect	44	179	45	180
rect	47	179	48	180
rect	56	179	57	180
rect	65	179	66	180
rect	95	179	96	180
rect	98	179	99	180
rect	107	179	108	180
rect	116	179	117	180
rect	119	179	120	180
rect	128	179	129	180
rect	140	179	141	180
rect	149	179	150	180
rect	152	179	153	180
rect	158	179	159	180
rect	161	179	162	180
rect	164	179	165	180
rect	167	179	168	180
rect	173	179	174	180
rect	186	179	187	180
rect	189	179	190	180
rect	192	179	193	180
rect	205	179	206	180
rect	208	179	209	180
rect	210	179	211	180
rect	216	179	217	180
rect	225	179	226	180
rect	228	179	229	180
rect	230	179	231	180
rect	233	179	234	180
rect	240	179	241	180
rect	242	179	243	180
rect	245	179	246	180
rect	248	179	249	180
rect	251	179	252	180
rect	254	179	255	180
rect	257	179	258	180
rect	261	179	262	180
rect	263	179	264	180
rect	266	179	267	180
rect	269	179	270	180
rect	272	179	273	180
rect	275	179	276	180
rect	278	179	279	180
rect	281	179	282	180
rect	288	179	289	180
rect	290	179	291	180
rect	293	179	294	180
rect	303	179	304	180
rect	305	179	306	180
rect	314	179	315	180
rect	317	179	318	180
rect	329	179	330	180
rect	332	179	333	180
rect	344	179	345	180
rect	346	179	347	180
rect	353	179	354	180
rect	359	179	360	180
rect	368	179	369	180
rect	370	179	371	180
rect	388	179	389	180
rect	391	179	392	180
rect	394	179	395	180
rect	410	179	411	180
rect	413	179	414	180
rect	8	180	9	181
rect	29	180	30	181
rect	35	180	36	181
rect	47	180	48	181
rect	56	180	57	181
rect	65	180	66	181
rect	95	180	96	181
rect	98	180	99	181
rect	107	180	108	181
rect	116	180	117	181
rect	119	180	120	181
rect	140	180	141	181
rect	149	180	150	181
rect	152	180	153	181
rect	158	180	159	181
rect	161	180	162	181
rect	164	180	165	181
rect	186	180	187	181
rect	189	180	190	181
rect	192	180	193	181
rect	205	180	206	181
rect	208	180	209	181
rect	210	180	211	181
rect	216	180	217	181
rect	225	180	226	181
rect	228	180	229	181
rect	230	180	231	181
rect	233	180	234	181
rect	240	180	241	181
rect	242	180	243	181
rect	245	180	246	181
rect	248	180	249	181
rect	251	180	252	181
rect	254	180	255	181
rect	257	180	258	181
rect	261	180	262	181
rect	263	180	264	181
rect	266	180	267	181
rect	269	180	270	181
rect	272	180	273	181
rect	275	180	276	181
rect	278	180	279	181
rect	281	180	282	181
rect	290	180	291	181
rect	293	180	294	181
rect	303	180	304	181
rect	305	180	306	181
rect	314	180	315	181
rect	317	180	318	181
rect	329	180	330	181
rect	332	180	333	181
rect	344	180	345	181
rect	353	180	354	181
rect	359	180	360	181
rect	368	180	369	181
rect	388	180	389	181
rect	391	180	392	181
rect	410	180	411	181
rect	413	180	414	181
rect	8	181	9	182
rect	29	181	30	182
rect	35	181	36	182
rect	42	181	43	182
rect	47	181	48	182
rect	56	181	57	182
rect	65	181	66	182
rect	95	181	96	182
rect	98	181	99	182
rect	107	181	108	182
rect	116	181	117	182
rect	119	181	120	182
rect	137	181	138	182
rect	140	181	141	182
rect	149	181	150	182
rect	152	181	153	182
rect	158	181	159	182
rect	161	181	162	182
rect	164	181	165	182
rect	168	181	169	182
rect	186	181	187	182
rect	189	181	190	182
rect	192	181	193	182
rect	205	181	206	182
rect	208	181	209	182
rect	210	181	211	182
rect	216	181	217	182
rect	225	181	226	182
rect	228	181	229	182
rect	230	181	231	182
rect	233	181	234	182
rect	240	181	241	182
rect	242	181	243	182
rect	245	181	246	182
rect	248	181	249	182
rect	251	181	252	182
rect	254	181	255	182
rect	257	181	258	182
rect	261	181	262	182
rect	263	181	264	182
rect	266	181	267	182
rect	269	181	270	182
rect	272	181	273	182
rect	275	181	276	182
rect	278	181	279	182
rect	281	181	282	182
rect	284	181	285	182
rect	290	181	291	182
rect	293	181	294	182
rect	296	181	297	182
rect	303	181	304	182
rect	305	181	306	182
rect	314	181	315	182
rect	317	181	318	182
rect	329	181	330	182
rect	332	181	333	182
rect	341	181	342	182
rect	344	181	345	182
rect	353	181	354	182
rect	356	181	357	182
rect	359	181	360	182
rect	368	181	369	182
rect	388	181	389	182
rect	391	181	392	182
rect	397	181	398	182
rect	410	181	411	182
rect	413	181	414	182
rect	8	182	9	183
rect	29	182	30	183
rect	42	182	43	183
rect	47	182	48	183
rect	56	182	57	183
rect	65	182	66	183
rect	95	182	96	183
rect	107	182	108	183
rect	116	182	117	183
rect	137	182	138	183
rect	140	182	141	183
rect	149	182	150	183
rect	152	182	153	183
rect	158	182	159	183
rect	161	182	162	183
rect	168	182	169	183
rect	192	182	193	183
rect	205	182	206	183
rect	208	182	209	183
rect	230	182	231	183
rect	233	182	234	183
rect	242	182	243	183
rect	245	182	246	183
rect	248	182	249	183
rect	251	182	252	183
rect	254	182	255	183
rect	257	182	258	183
rect	263	182	264	183
rect	266	182	267	183
rect	269	182	270	183
rect	272	182	273	183
rect	275	182	276	183
rect	278	182	279	183
rect	281	182	282	183
rect	284	182	285	183
rect	290	182	291	183
rect	293	182	294	183
rect	296	182	297	183
rect	303	182	304	183
rect	305	182	306	183
rect	314	182	315	183
rect	317	182	318	183
rect	329	182	330	183
rect	332	182	333	183
rect	341	182	342	183
rect	344	182	345	183
rect	353	182	354	183
rect	356	182	357	183
rect	359	182	360	183
rect	368	182	369	183
rect	397	182	398	183
rect	410	182	411	183
rect	8	183	9	184
rect	29	183	30	184
rect	42	183	43	184
rect	45	183	46	184
rect	47	183	48	184
rect	56	183	57	184
rect	65	183	66	184
rect	95	183	96	184
rect	100	183	101	184
rect	107	183	108	184
rect	116	183	117	184
rect	128	183	129	184
rect	137	183	138	184
rect	140	183	141	184
rect	149	183	150	184
rect	152	183	153	184
rect	158	183	159	184
rect	161	183	162	184
rect	168	183	169	184
rect	174	183	175	184
rect	183	183	184	184
rect	192	183	193	184
rect	202	183	203	184
rect	205	183	206	184
rect	208	183	209	184
rect	211	183	212	184
rect	214	183	215	184
rect	220	183	221	184
rect	230	183	231	184
rect	233	183	234	184
rect	242	183	243	184
rect	245	183	246	184
rect	248	183	249	184
rect	251	183	252	184
rect	254	183	255	184
rect	257	183	258	184
rect	263	183	264	184
rect	266	183	267	184
rect	269	183	270	184
rect	272	183	273	184
rect	275	183	276	184
rect	278	183	279	184
rect	281	183	282	184
rect	284	183	285	184
rect	290	183	291	184
rect	293	183	294	184
rect	296	183	297	184
rect	303	183	304	184
rect	305	183	306	184
rect	314	183	315	184
rect	317	183	318	184
rect	329	183	330	184
rect	332	183	333	184
rect	341	183	342	184
rect	344	183	345	184
rect	353	183	354	184
rect	356	183	357	184
rect	359	183	360	184
rect	368	183	369	184
rect	371	183	372	184
rect	394	183	395	184
rect	397	183	398	184
rect	410	183	411	184
rect	42	184	43	185
rect	45	184	46	185
rect	100	184	101	185
rect	116	184	117	185
rect	128	184	129	185
rect	137	184	138	185
rect	140	184	141	185
rect	149	184	150	185
rect	152	184	153	185
rect	158	184	159	185
rect	168	184	169	185
rect	174	184	175	185
rect	183	184	184	185
rect	192	184	193	185
rect	202	184	203	185
rect	205	184	206	185
rect	208	184	209	185
rect	211	184	212	185
rect	214	184	215	185
rect	220	184	221	185
rect	230	184	231	185
rect	233	184	234	185
rect	242	184	243	185
rect	245	184	246	185
rect	248	184	249	185
rect	251	184	252	185
rect	254	184	255	185
rect	257	184	258	185
rect	263	184	264	185
rect	266	184	267	185
rect	269	184	270	185
rect	272	184	273	185
rect	275	184	276	185
rect	278	184	279	185
rect	281	184	282	185
rect	284	184	285	185
rect	290	184	291	185
rect	293	184	294	185
rect	296	184	297	185
rect	305	184	306	185
rect	314	184	315	185
rect	317	184	318	185
rect	329	184	330	185
rect	332	184	333	185
rect	341	184	342	185
rect	344	184	345	185
rect	353	184	354	185
rect	356	184	357	185
rect	359	184	360	185
rect	368	184	369	185
rect	371	184	372	185
rect	394	184	395	185
rect	397	184	398	185
rect	14	185	15	186
rect	30	185	31	186
rect	36	185	37	186
rect	39	185	40	186
rect	42	185	43	186
rect	45	185	46	186
rect	48	185	49	186
rect	51	185	52	186
rect	67	185	68	186
rect	97	185	98	186
rect	100	185	101	186
rect	116	185	117	186
rect	119	185	120	186
rect	128	185	129	186
rect	137	185	138	186
rect	140	185	141	186
rect	149	185	150	186
rect	152	185	153	186
rect	158	185	159	186
rect	168	185	169	186
rect	171	185	172	186
rect	174	185	175	186
rect	183	185	184	186
rect	186	185	187	186
rect	192	185	193	186
rect	202	185	203	186
rect	205	185	206	186
rect	208	185	209	186
rect	211	185	212	186
rect	214	185	215	186
rect	220	185	221	186
rect	230	185	231	186
rect	233	185	234	186
rect	242	185	243	186
rect	245	185	246	186
rect	248	185	249	186
rect	251	185	252	186
rect	254	185	255	186
rect	257	185	258	186
rect	263	185	264	186
rect	266	185	267	186
rect	269	185	270	186
rect	272	185	273	186
rect	275	185	276	186
rect	278	185	279	186
rect	281	185	282	186
rect	284	185	285	186
rect	290	185	291	186
rect	293	185	294	186
rect	296	185	297	186
rect	305	185	306	186
rect	314	185	315	186
rect	317	185	318	186
rect	326	185	327	186
rect	329	185	330	186
rect	332	185	333	186
rect	341	185	342	186
rect	344	185	345	186
rect	353	185	354	186
rect	356	185	357	186
rect	359	185	360	186
rect	368	185	369	186
rect	371	185	372	186
rect	388	185	389	186
rect	391	185	392	186
rect	394	185	395	186
rect	397	185	398	186
rect	8	192	9	193
rect	14	192	15	193
rect	24	192	25	193
rect	27	192	28	193
rect	30	192	31	193
rect	39	192	40	193
rect	42	192	43	193
rect	45	192	46	193
rect	48	192	49	193
rect	51	192	52	193
rect	61	192	62	193
rect	67	192	68	193
rect	97	192	98	193
rect	100	192	101	193
rect	116	192	117	193
rect	119	192	120	193
rect	128	192	129	193
rect	137	192	138	193
rect	140	192	141	193
rect	149	192	150	193
rect	152	192	153	193
rect	168	192	169	193
rect	171	192	172	193
rect	174	192	175	193
rect	180	192	181	193
rect	183	192	184	193
rect	186	192	187	193
rect	202	192	203	193
rect	205	192	206	193
rect	208	192	209	193
rect	211	192	212	193
rect	214	192	215	193
rect	227	192	228	193
rect	230	192	231	193
rect	233	192	234	193
rect	242	192	243	193
rect	245	192	246	193
rect	248	192	249	193
rect	251	192	252	193
rect	254	192	255	193
rect	257	192	258	193
rect	260	192	261	193
rect	266	192	267	193
rect	269	192	270	193
rect	278	192	279	193
rect	281	192	282	193
rect	290	192	291	193
rect	293	192	294	193
rect	296	192	297	193
rect	305	192	306	193
rect	314	192	315	193
rect	317	192	318	193
rect	320	192	321	193
rect	326	192	327	193
rect	329	192	330	193
rect	332	192	333	193
rect	338	192	339	193
rect	341	192	342	193
rect	344	192	345	193
rect	353	192	354	193
rect	356	192	357	193
rect	359	192	360	193
rect	368	192	369	193
rect	385	192	386	193
rect	388	192	389	193
rect	391	192	392	193
rect	394	192	395	193
rect	397	192	398	193
rect	8	193	9	194
rect	14	193	15	194
rect	24	193	25	194
rect	27	193	28	194
rect	30	193	31	194
rect	39	193	40	194
rect	42	193	43	194
rect	45	193	46	194
rect	48	193	49	194
rect	51	193	52	194
rect	61	193	62	194
rect	67	193	68	194
rect	97	193	98	194
rect	100	193	101	194
rect	116	193	117	194
rect	119	193	120	194
rect	128	193	129	194
rect	137	193	138	194
rect	140	193	141	194
rect	149	193	150	194
rect	152	193	153	194
rect	168	193	169	194
rect	171	193	172	194
rect	174	193	175	194
rect	180	193	181	194
rect	183	193	184	194
rect	186	193	187	194
rect	202	193	203	194
rect	205	193	206	194
rect	208	193	209	194
rect	211	193	212	194
rect	214	193	215	194
rect	227	193	228	194
rect	230	193	231	194
rect	233	193	234	194
rect	242	193	243	194
rect	245	193	246	194
rect	248	193	249	194
rect	251	193	252	194
rect	254	193	255	194
rect	257	193	258	194
rect	260	193	261	194
rect	266	193	267	194
rect	269	193	270	194
rect	278	193	279	194
rect	281	193	282	194
rect	290	193	291	194
rect	293	193	294	194
rect	296	193	297	194
rect	305	193	306	194
rect	314	193	315	194
rect	317	193	318	194
rect	320	193	321	194
rect	326	193	327	194
rect	329	193	330	194
rect	338	193	339	194
rect	341	193	342	194
rect	344	193	345	194
rect	353	193	354	194
rect	356	193	357	194
rect	359	193	360	194
rect	368	193	369	194
rect	385	193	386	194
rect	388	193	389	194
rect	391	193	392	194
rect	394	193	395	194
rect	397	193	398	194
rect	8	194	9	195
rect	14	194	15	195
rect	24	194	25	195
rect	27	194	28	195
rect	30	194	31	195
rect	39	194	40	195
rect	42	194	43	195
rect	45	194	46	195
rect	48	194	49	195
rect	51	194	52	195
rect	61	194	62	195
rect	67	194	68	195
rect	97	194	98	195
rect	100	194	101	195
rect	116	194	117	195
rect	119	194	120	195
rect	128	194	129	195
rect	137	194	138	195
rect	140	194	141	195
rect	149	194	150	195
rect	152	194	153	195
rect	168	194	169	195
rect	171	194	172	195
rect	174	194	175	195
rect	180	194	181	195
rect	183	194	184	195
rect	186	194	187	195
rect	202	194	203	195
rect	205	194	206	195
rect	208	194	209	195
rect	211	194	212	195
rect	214	194	215	195
rect	227	194	228	195
rect	230	194	231	195
rect	233	194	234	195
rect	242	194	243	195
rect	245	194	246	195
rect	248	194	249	195
rect	251	194	252	195
rect	254	194	255	195
rect	257	194	258	195
rect	260	194	261	195
rect	266	194	267	195
rect	269	194	270	195
rect	278	194	279	195
rect	281	194	282	195
rect	290	194	291	195
rect	293	194	294	195
rect	296	194	297	195
rect	305	194	306	195
rect	312	194	313	195
rect	314	194	315	195
rect	317	194	318	195
rect	320	194	321	195
rect	326	194	327	195
rect	329	194	330	195
rect	338	194	339	195
rect	341	194	342	195
rect	344	194	345	195
rect	353	194	354	195
rect	356	194	357	195
rect	359	194	360	195
rect	368	194	369	195
rect	385	194	386	195
rect	388	194	389	195
rect	391	194	392	195
rect	394	194	395	195
rect	397	194	398	195
rect	8	195	9	196
rect	14	195	15	196
rect	24	195	25	196
rect	27	195	28	196
rect	30	195	31	196
rect	39	195	40	196
rect	42	195	43	196
rect	45	195	46	196
rect	48	195	49	196
rect	51	195	52	196
rect	61	195	62	196
rect	67	195	68	196
rect	97	195	98	196
rect	100	195	101	196
rect	116	195	117	196
rect	119	195	120	196
rect	128	195	129	196
rect	137	195	138	196
rect	140	195	141	196
rect	149	195	150	196
rect	152	195	153	196
rect	168	195	169	196
rect	171	195	172	196
rect	174	195	175	196
rect	180	195	181	196
rect	183	195	184	196
rect	186	195	187	196
rect	202	195	203	196
rect	205	195	206	196
rect	208	195	209	196
rect	211	195	212	196
rect	214	195	215	196
rect	227	195	228	196
rect	230	195	231	196
rect	233	195	234	196
rect	242	195	243	196
rect	245	195	246	196
rect	248	195	249	196
rect	251	195	252	196
rect	254	195	255	196
rect	257	195	258	196
rect	260	195	261	196
rect	266	195	267	196
rect	269	195	270	196
rect	278	195	279	196
rect	281	195	282	196
rect	290	195	291	196
rect	293	195	294	196
rect	296	195	297	196
rect	305	195	306	196
rect	312	195	313	196
rect	314	195	315	196
rect	317	195	318	196
rect	320	195	321	196
rect	329	195	330	196
rect	338	195	339	196
rect	341	195	342	196
rect	344	195	345	196
rect	353	195	354	196
rect	356	195	357	196
rect	359	195	360	196
rect	368	195	369	196
rect	385	195	386	196
rect	388	195	389	196
rect	391	195	392	196
rect	394	195	395	196
rect	397	195	398	196
rect	8	196	9	197
rect	14	196	15	197
rect	24	196	25	197
rect	27	196	28	197
rect	30	196	31	197
rect	39	196	40	197
rect	42	196	43	197
rect	45	196	46	197
rect	48	196	49	197
rect	51	196	52	197
rect	61	196	62	197
rect	67	196	68	197
rect	97	196	98	197
rect	100	196	101	197
rect	116	196	117	197
rect	119	196	120	197
rect	128	196	129	197
rect	137	196	138	197
rect	140	196	141	197
rect	149	196	150	197
rect	152	196	153	197
rect	168	196	169	197
rect	171	196	172	197
rect	174	196	175	197
rect	180	196	181	197
rect	183	196	184	197
rect	186	196	187	197
rect	202	196	203	197
rect	205	196	206	197
rect	208	196	209	197
rect	211	196	212	197
rect	214	196	215	197
rect	227	196	228	197
rect	230	196	231	197
rect	233	196	234	197
rect	242	196	243	197
rect	245	196	246	197
rect	248	196	249	197
rect	251	196	252	197
rect	254	196	255	197
rect	257	196	258	197
rect	260	196	261	197
rect	266	196	267	197
rect	269	196	270	197
rect	278	196	279	197
rect	281	196	282	197
rect	290	196	291	197
rect	293	196	294	197
rect	296	196	297	197
rect	305	196	306	197
rect	310	196	311	197
rect	312	196	313	197
rect	314	196	315	197
rect	317	196	318	197
rect	320	196	321	197
rect	329	196	330	197
rect	338	196	339	197
rect	341	196	342	197
rect	344	196	345	197
rect	353	196	354	197
rect	356	196	357	197
rect	359	196	360	197
rect	368	196	369	197
rect	385	196	386	197
rect	388	196	389	197
rect	391	196	392	197
rect	394	196	395	197
rect	397	196	398	197
rect	8	197	9	198
rect	14	197	15	198
rect	24	197	25	198
rect	27	197	28	198
rect	30	197	31	198
rect	39	197	40	198
rect	42	197	43	198
rect	45	197	46	198
rect	48	197	49	198
rect	51	197	52	198
rect	61	197	62	198
rect	67	197	68	198
rect	97	197	98	198
rect	100	197	101	198
rect	116	197	117	198
rect	119	197	120	198
rect	128	197	129	198
rect	137	197	138	198
rect	140	197	141	198
rect	149	197	150	198
rect	152	197	153	198
rect	168	197	169	198
rect	171	197	172	198
rect	174	197	175	198
rect	180	197	181	198
rect	183	197	184	198
rect	186	197	187	198
rect	202	197	203	198
rect	208	197	209	198
rect	211	197	212	198
rect	214	197	215	198
rect	230	197	231	198
rect	233	197	234	198
rect	242	197	243	198
rect	245	197	246	198
rect	248	197	249	198
rect	251	197	252	198
rect	254	197	255	198
rect	257	197	258	198
rect	260	197	261	198
rect	266	197	267	198
rect	269	197	270	198
rect	278	197	279	198
rect	281	197	282	198
rect	290	197	291	198
rect	293	197	294	198
rect	296	197	297	198
rect	305	197	306	198
rect	310	197	311	198
rect	312	197	313	198
rect	314	197	315	198
rect	320	197	321	198
rect	329	197	330	198
rect	338	197	339	198
rect	341	197	342	198
rect	344	197	345	198
rect	353	197	354	198
rect	356	197	357	198
rect	359	197	360	198
rect	368	197	369	198
rect	385	197	386	198
rect	388	197	389	198
rect	391	197	392	198
rect	394	197	395	198
rect	397	197	398	198
rect	8	198	9	199
rect	14	198	15	199
rect	24	198	25	199
rect	27	198	28	199
rect	30	198	31	199
rect	39	198	40	199
rect	42	198	43	199
rect	45	198	46	199
rect	48	198	49	199
rect	51	198	52	199
rect	61	198	62	199
rect	67	198	68	199
rect	97	198	98	199
rect	100	198	101	199
rect	116	198	117	199
rect	119	198	120	199
rect	128	198	129	199
rect	137	198	138	199
rect	140	198	141	199
rect	149	198	150	199
rect	152	198	153	199
rect	168	198	169	199
rect	171	198	172	199
rect	174	198	175	199
rect	180	198	181	199
rect	183	198	184	199
rect	186	198	187	199
rect	202	198	203	199
rect	208	198	209	199
rect	211	198	212	199
rect	214	198	215	199
rect	230	198	231	199
rect	233	198	234	199
rect	242	198	243	199
rect	245	198	246	199
rect	248	198	249	199
rect	251	198	252	199
rect	254	198	255	199
rect	257	198	258	199
rect	260	198	261	199
rect	266	198	267	199
rect	269	198	270	199
rect	278	198	279	199
rect	281	198	282	199
rect	290	198	291	199
rect	293	198	294	199
rect	296	198	297	199
rect	305	198	306	199
rect	310	198	311	199
rect	312	198	313	199
rect	314	198	315	199
rect	320	198	321	199
rect	325	198	326	199
rect	329	198	330	199
rect	338	198	339	199
rect	341	198	342	199
rect	344	198	345	199
rect	353	198	354	199
rect	356	198	357	199
rect	359	198	360	199
rect	368	198	369	199
rect	385	198	386	199
rect	388	198	389	199
rect	391	198	392	199
rect	394	198	395	199
rect	397	198	398	199
rect	8	199	9	200
rect	14	199	15	200
rect	24	199	25	200
rect	27	199	28	200
rect	30	199	31	200
rect	39	199	40	200
rect	42	199	43	200
rect	45	199	46	200
rect	48	199	49	200
rect	51	199	52	200
rect	61	199	62	200
rect	67	199	68	200
rect	97	199	98	200
rect	100	199	101	200
rect	116	199	117	200
rect	119	199	120	200
rect	128	199	129	200
rect	137	199	138	200
rect	140	199	141	200
rect	149	199	150	200
rect	152	199	153	200
rect	168	199	169	200
rect	171	199	172	200
rect	174	199	175	200
rect	180	199	181	200
rect	183	199	184	200
rect	186	199	187	200
rect	202	199	203	200
rect	208	199	209	200
rect	211	199	212	200
rect	230	199	231	200
rect	233	199	234	200
rect	242	199	243	200
rect	245	199	246	200
rect	248	199	249	200
rect	251	199	252	200
rect	254	199	255	200
rect	257	199	258	200
rect	260	199	261	200
rect	266	199	267	200
rect	269	199	270	200
rect	278	199	279	200
rect	281	199	282	200
rect	290	199	291	200
rect	293	199	294	200
rect	296	199	297	200
rect	305	199	306	200
rect	310	199	311	200
rect	312	199	313	200
rect	314	199	315	200
rect	325	199	326	200
rect	329	199	330	200
rect	338	199	339	200
rect	341	199	342	200
rect	344	199	345	200
rect	353	199	354	200
rect	356	199	357	200
rect	359	199	360	200
rect	368	199	369	200
rect	385	199	386	200
rect	388	199	389	200
rect	391	199	392	200
rect	394	199	395	200
rect	397	199	398	200
rect	8	200	9	201
rect	14	200	15	201
rect	24	200	25	201
rect	27	200	28	201
rect	30	200	31	201
rect	39	200	40	201
rect	42	200	43	201
rect	45	200	46	201
rect	48	200	49	201
rect	51	200	52	201
rect	61	200	62	201
rect	67	200	68	201
rect	97	200	98	201
rect	100	200	101	201
rect	116	200	117	201
rect	119	200	120	201
rect	128	200	129	201
rect	137	200	138	201
rect	140	200	141	201
rect	149	200	150	201
rect	152	200	153	201
rect	168	200	169	201
rect	171	200	172	201
rect	174	200	175	201
rect	180	200	181	201
rect	183	200	184	201
rect	186	200	187	201
rect	202	200	203	201
rect	206	200	207	201
rect	208	200	209	201
rect	211	200	212	201
rect	230	200	231	201
rect	233	200	234	201
rect	242	200	243	201
rect	245	200	246	201
rect	248	200	249	201
rect	251	200	252	201
rect	254	200	255	201
rect	257	200	258	201
rect	260	200	261	201
rect	266	200	267	201
rect	269	200	270	201
rect	278	200	279	201
rect	281	200	282	201
rect	290	200	291	201
rect	293	200	294	201
rect	296	200	297	201
rect	305	200	306	201
rect	310	200	311	201
rect	312	200	313	201
rect	314	200	315	201
rect	316	200	317	201
rect	325	200	326	201
rect	329	200	330	201
rect	338	200	339	201
rect	341	200	342	201
rect	344	200	345	201
rect	353	200	354	201
rect	356	200	357	201
rect	359	200	360	201
rect	368	200	369	201
rect	385	200	386	201
rect	388	200	389	201
rect	391	200	392	201
rect	394	200	395	201
rect	397	200	398	201
rect	8	201	9	202
rect	14	201	15	202
rect	24	201	25	202
rect	27	201	28	202
rect	30	201	31	202
rect	39	201	40	202
rect	42	201	43	202
rect	45	201	46	202
rect	48	201	49	202
rect	51	201	52	202
rect	61	201	62	202
rect	67	201	68	202
rect	97	201	98	202
rect	100	201	101	202
rect	116	201	117	202
rect	119	201	120	202
rect	128	201	129	202
rect	137	201	138	202
rect	140	201	141	202
rect	149	201	150	202
rect	152	201	153	202
rect	168	201	169	202
rect	171	201	172	202
rect	174	201	175	202
rect	180	201	181	202
rect	183	201	184	202
rect	186	201	187	202
rect	202	201	203	202
rect	206	201	207	202
rect	208	201	209	202
rect	230	201	231	202
rect	233	201	234	202
rect	245	201	246	202
rect	248	201	249	202
rect	251	201	252	202
rect	254	201	255	202
rect	257	201	258	202
rect	266	201	267	202
rect	269	201	270	202
rect	278	201	279	202
rect	281	201	282	202
rect	290	201	291	202
rect	293	201	294	202
rect	296	201	297	202
rect	305	201	306	202
rect	310	201	311	202
rect	312	201	313	202
rect	314	201	315	202
rect	316	201	317	202
rect	325	201	326	202
rect	329	201	330	202
rect	338	201	339	202
rect	341	201	342	202
rect	353	201	354	202
rect	356	201	357	202
rect	359	201	360	202
rect	368	201	369	202
rect	385	201	386	202
rect	388	201	389	202
rect	391	201	392	202
rect	394	201	395	202
rect	397	201	398	202
rect	8	202	9	203
rect	14	202	15	203
rect	24	202	25	203
rect	27	202	28	203
rect	30	202	31	203
rect	39	202	40	203
rect	42	202	43	203
rect	45	202	46	203
rect	48	202	49	203
rect	51	202	52	203
rect	61	202	62	203
rect	67	202	68	203
rect	97	202	98	203
rect	100	202	101	203
rect	116	202	117	203
rect	119	202	120	203
rect	128	202	129	203
rect	137	202	138	203
rect	140	202	141	203
rect	149	202	150	203
rect	152	202	153	203
rect	168	202	169	203
rect	171	202	172	203
rect	174	202	175	203
rect	180	202	181	203
rect	183	202	184	203
rect	186	202	187	203
rect	202	202	203	203
rect	206	202	207	203
rect	208	202	209	203
rect	215	202	216	203
rect	230	202	231	203
rect	233	202	234	203
rect	245	202	246	203
rect	248	202	249	203
rect	251	202	252	203
rect	254	202	255	203
rect	257	202	258	203
rect	266	202	267	203
rect	269	202	270	203
rect	278	202	279	203
rect	281	202	282	203
rect	290	202	291	203
rect	293	202	294	203
rect	296	202	297	203
rect	305	202	306	203
rect	310	202	311	203
rect	312	202	313	203
rect	314	202	315	203
rect	316	202	317	203
rect	319	202	320	203
rect	325	202	326	203
rect	329	202	330	203
rect	338	202	339	203
rect	341	202	342	203
rect	353	202	354	203
rect	356	202	357	203
rect	359	202	360	203
rect	368	202	369	203
rect	385	202	386	203
rect	388	202	389	203
rect	391	202	392	203
rect	394	202	395	203
rect	397	202	398	203
rect	8	203	9	204
rect	14	203	15	204
rect	24	203	25	204
rect	27	203	28	204
rect	30	203	31	204
rect	39	203	40	204
rect	42	203	43	204
rect	45	203	46	204
rect	51	203	52	204
rect	61	203	62	204
rect	67	203	68	204
rect	97	203	98	204
rect	100	203	101	204
rect	116	203	117	204
rect	119	203	120	204
rect	128	203	129	204
rect	137	203	138	204
rect	140	203	141	204
rect	149	203	150	204
rect	152	203	153	204
rect	168	203	169	204
rect	171	203	172	204
rect	174	203	175	204
rect	180	203	181	204
rect	183	203	184	204
rect	186	203	187	204
rect	202	203	203	204
rect	206	203	207	204
rect	208	203	209	204
rect	215	203	216	204
rect	230	203	231	204
rect	233	203	234	204
rect	245	203	246	204
rect	251	203	252	204
rect	254	203	255	204
rect	257	203	258	204
rect	266	203	267	204
rect	269	203	270	204
rect	278	203	279	204
rect	281	203	282	204
rect	290	203	291	204
rect	293	203	294	204
rect	296	203	297	204
rect	305	203	306	204
rect	310	203	311	204
rect	312	203	313	204
rect	314	203	315	204
rect	316	203	317	204
rect	319	203	320	204
rect	325	203	326	204
rect	338	203	339	204
rect	341	203	342	204
rect	353	203	354	204
rect	356	203	357	204
rect	359	203	360	204
rect	385	203	386	204
rect	388	203	389	204
rect	391	203	392	204
rect	394	203	395	204
rect	397	203	398	204
rect	8	204	9	205
rect	14	204	15	205
rect	24	204	25	205
rect	27	204	28	205
rect	30	204	31	205
rect	39	204	40	205
rect	42	204	43	205
rect	45	204	46	205
rect	51	204	52	205
rect	56	204	57	205
rect	61	204	62	205
rect	67	204	68	205
rect	97	204	98	205
rect	100	204	101	205
rect	116	204	117	205
rect	119	204	120	205
rect	128	204	129	205
rect	137	204	138	205
rect	140	204	141	205
rect	149	204	150	205
rect	152	204	153	205
rect	168	204	169	205
rect	171	204	172	205
rect	174	204	175	205
rect	180	204	181	205
rect	183	204	184	205
rect	186	204	187	205
rect	202	204	203	205
rect	206	204	207	205
rect	208	204	209	205
rect	212	204	213	205
rect	215	204	216	205
rect	230	204	231	205
rect	233	204	234	205
rect	245	204	246	205
rect	251	204	252	205
rect	254	204	255	205
rect	257	204	258	205
rect	266	204	267	205
rect	269	204	270	205
rect	278	204	279	205
rect	281	204	282	205
rect	290	204	291	205
rect	293	204	294	205
rect	296	204	297	205
rect	305	204	306	205
rect	310	204	311	205
rect	312	204	313	205
rect	314	204	315	205
rect	316	204	317	205
rect	319	204	320	205
rect	325	204	326	205
rect	331	204	332	205
rect	338	204	339	205
rect	341	204	342	205
rect	343	204	344	205
rect	353	204	354	205
rect	356	204	357	205
rect	359	204	360	205
rect	385	204	386	205
rect	388	204	389	205
rect	391	204	392	205
rect	394	204	395	205
rect	397	204	398	205
rect	8	205	9	206
rect	14	205	15	206
rect	24	205	25	206
rect	27	205	28	206
rect	30	205	31	206
rect	39	205	40	206
rect	42	205	43	206
rect	51	205	52	206
rect	56	205	57	206
rect	61	205	62	206
rect	67	205	68	206
rect	97	205	98	206
rect	100	205	101	206
rect	116	205	117	206
rect	119	205	120	206
rect	128	205	129	206
rect	137	205	138	206
rect	140	205	141	206
rect	152	205	153	206
rect	168	205	169	206
rect	171	205	172	206
rect	174	205	175	206
rect	180	205	181	206
rect	183	205	184	206
rect	186	205	187	206
rect	202	205	203	206
rect	206	205	207	206
rect	208	205	209	206
rect	212	205	213	206
rect	215	205	216	206
rect	230	205	231	206
rect	233	205	234	206
rect	245	205	246	206
rect	251	205	252	206
rect	254	205	255	206
rect	278	205	279	206
rect	290	205	291	206
rect	293	205	294	206
rect	296	205	297	206
rect	305	205	306	206
rect	310	205	311	206
rect	312	205	313	206
rect	314	205	315	206
rect	316	205	317	206
rect	319	205	320	206
rect	325	205	326	206
rect	331	205	332	206
rect	338	205	339	206
rect	343	205	344	206
rect	353	205	354	206
rect	356	205	357	206
rect	359	205	360	206
rect	385	205	386	206
rect	388	205	389	206
rect	391	205	392	206
rect	394	205	395	206
rect	397	205	398	206
rect	8	206	9	207
rect	14	206	15	207
rect	24	206	25	207
rect	27	206	28	207
rect	30	206	31	207
rect	39	206	40	207
rect	42	206	43	207
rect	51	206	52	207
rect	53	206	54	207
rect	56	206	57	207
rect	61	206	62	207
rect	67	206	68	207
rect	97	206	98	207
rect	100	206	101	207
rect	116	206	117	207
rect	119	206	120	207
rect	128	206	129	207
rect	137	206	138	207
rect	140	206	141	207
rect	152	206	153	207
rect	159	206	160	207
rect	168	206	169	207
rect	171	206	172	207
rect	174	206	175	207
rect	180	206	181	207
rect	183	206	184	207
rect	186	206	187	207
rect	202	206	203	207
rect	206	206	207	207
rect	208	206	209	207
rect	212	206	213	207
rect	215	206	216	207
rect	230	206	231	207
rect	233	206	234	207
rect	245	206	246	207
rect	249	206	250	207
rect	251	206	252	207
rect	254	206	255	207
rect	261	206	262	207
rect	273	206	274	207
rect	278	206	279	207
rect	285	206	286	207
rect	290	206	291	207
rect	293	206	294	207
rect	296	206	297	207
rect	305	206	306	207
rect	307	206	308	207
rect	310	206	311	207
rect	312	206	313	207
rect	314	206	315	207
rect	316	206	317	207
rect	319	206	320	207
rect	325	206	326	207
rect	331	206	332	207
rect	338	206	339	207
rect	343	206	344	207
rect	353	206	354	207
rect	356	206	357	207
rect	359	206	360	207
rect	385	206	386	207
rect	388	206	389	207
rect	391	206	392	207
rect	394	206	395	207
rect	397	206	398	207
rect	8	207	9	208
rect	14	207	15	208
rect	24	207	25	208
rect	27	207	28	208
rect	30	207	31	208
rect	42	207	43	208
rect	51	207	52	208
rect	53	207	54	208
rect	56	207	57	208
rect	61	207	62	208
rect	67	207	68	208
rect	97	207	98	208
rect	116	207	117	208
rect	128	207	129	208
rect	140	207	141	208
rect	152	207	153	208
rect	159	207	160	208
rect	168	207	169	208
rect	171	207	172	208
rect	174	207	175	208
rect	186	207	187	208
rect	202	207	203	208
rect	206	207	207	208
rect	208	207	209	208
rect	212	207	213	208
rect	215	207	216	208
rect	230	207	231	208
rect	233	207	234	208
rect	249	207	250	208
rect	251	207	252	208
rect	254	207	255	208
rect	261	207	262	208
rect	273	207	274	208
rect	278	207	279	208
rect	285	207	286	208
rect	293	207	294	208
rect	296	207	297	208
rect	307	207	308	208
rect	310	207	311	208
rect	314	207	315	208
rect	316	207	317	208
rect	319	207	320	208
rect	325	207	326	208
rect	331	207	332	208
rect	338	207	339	208
rect	343	207	344	208
rect	356	207	357	208
rect	359	207	360	208
rect	385	207	386	208
rect	388	207	389	208
rect	391	207	392	208
rect	394	207	395	208
rect	397	207	398	208
rect	8	208	9	209
rect	14	208	15	209
rect	24	208	25	209
rect	27	208	28	209
rect	30	208	31	209
rect	42	208	43	209
rect	47	208	48	209
rect	51	208	52	209
rect	53	208	54	209
rect	56	208	57	209
rect	61	208	62	209
rect	67	208	68	209
rect	97	208	98	209
rect	101	208	102	209
rect	116	208	117	209
rect	126	208	127	209
rect	128	208	129	209
rect	140	208	141	209
rect	150	208	151	209
rect	152	208	153	209
rect	159	208	160	209
rect	168	208	169	209
rect	171	208	172	209
rect	174	208	175	209
rect	186	208	187	209
rect	202	208	203	209
rect	206	208	207	209
rect	208	208	209	209
rect	212	208	213	209
rect	215	208	216	209
rect	224	208	225	209
rect	230	208	231	209
rect	233	208	234	209
rect	249	208	250	209
rect	251	208	252	209
rect	254	208	255	209
rect	258	208	259	209
rect	261	208	262	209
rect	273	208	274	209
rect	278	208	279	209
rect	285	208	286	209
rect	293	208	294	209
rect	296	208	297	209
rect	304	208	305	209
rect	307	208	308	209
rect	310	208	311	209
rect	314	208	315	209
rect	316	208	317	209
rect	319	208	320	209
rect	325	208	326	209
rect	328	208	329	209
rect	331	208	332	209
rect	338	208	339	209
rect	340	208	341	209
rect	343	208	344	209
rect	356	208	357	209
rect	359	208	360	209
rect	385	208	386	209
rect	388	208	389	209
rect	391	208	392	209
rect	394	208	395	209
rect	397	208	398	209
rect	8	209	9	210
rect	14	209	15	210
rect	24	209	25	210
rect	30	209	31	210
rect	42	209	43	210
rect	47	209	48	210
rect	51	209	52	210
rect	53	209	54	210
rect	56	209	57	210
rect	61	209	62	210
rect	67	209	68	210
rect	97	209	98	210
rect	101	209	102	210
rect	116	209	117	210
rect	126	209	127	210
rect	128	209	129	210
rect	140	209	141	210
rect	150	209	151	210
rect	152	209	153	210
rect	159	209	160	210
rect	168	209	169	210
rect	171	209	172	210
rect	174	209	175	210
rect	186	209	187	210
rect	202	209	203	210
rect	206	209	207	210
rect	208	209	209	210
rect	212	209	213	210
rect	215	209	216	210
rect	224	209	225	210
rect	230	209	231	210
rect	233	209	234	210
rect	249	209	250	210
rect	251	209	252	210
rect	254	209	255	210
rect	258	209	259	210
rect	261	209	262	210
rect	273	209	274	210
rect	278	209	279	210
rect	285	209	286	210
rect	296	209	297	210
rect	304	209	305	210
rect	307	209	308	210
rect	310	209	311	210
rect	316	209	317	210
rect	319	209	320	210
rect	325	209	326	210
rect	328	209	329	210
rect	331	209	332	210
rect	338	209	339	210
rect	340	209	341	210
rect	343	209	344	210
rect	359	209	360	210
rect	385	209	386	210
rect	391	209	392	210
rect	394	209	395	210
rect	8	210	9	211
rect	14	210	15	211
rect	24	210	25	211
rect	30	210	31	211
rect	42	210	43	211
rect	47	210	48	211
rect	51	210	52	211
rect	53	210	54	211
rect	56	210	57	211
rect	61	210	62	211
rect	67	210	68	211
rect	97	210	98	211
rect	101	210	102	211
rect	116	210	117	211
rect	126	210	127	211
rect	128	210	129	211
rect	140	210	141	211
rect	150	210	151	211
rect	152	210	153	211
rect	159	210	160	211
rect	168	210	169	211
rect	171	210	172	211
rect	174	210	175	211
rect	186	210	187	211
rect	202	210	203	211
rect	206	210	207	211
rect	208	210	209	211
rect	212	210	213	211
rect	215	210	216	211
rect	224	210	225	211
rect	230	210	231	211
rect	233	210	234	211
rect	249	210	250	211
rect	251	210	252	211
rect	254	210	255	211
rect	258	210	259	211
rect	261	210	262	211
rect	264	210	265	211
rect	267	210	268	211
rect	273	210	274	211
rect	278	210	279	211
rect	285	210	286	211
rect	296	210	297	211
rect	301	210	302	211
rect	304	210	305	211
rect	307	210	308	211
rect	310	210	311	211
rect	316	210	317	211
rect	319	210	320	211
rect	322	210	323	211
rect	325	210	326	211
rect	328	210	329	211
rect	331	210	332	211
rect	338	210	339	211
rect	340	210	341	211
rect	343	210	344	211
rect	359	210	360	211
rect	385	210	386	211
rect	391	210	392	211
rect	394	210	395	211
rect	8	211	9	212
rect	24	211	25	212
rect	42	211	43	212
rect	47	211	48	212
rect	53	211	54	212
rect	56	211	57	212
rect	61	211	62	212
rect	101	211	102	212
rect	126	211	127	212
rect	150	211	151	212
rect	159	211	160	212
rect	168	211	169	212
rect	171	211	172	212
rect	186	211	187	212
rect	202	211	203	212
rect	206	211	207	212
rect	208	211	209	212
rect	212	211	213	212
rect	215	211	216	212
rect	224	211	225	212
rect	230	211	231	212
rect	249	211	250	212
rect	251	211	252	212
rect	258	211	259	212
rect	261	211	262	212
rect	264	211	265	212
rect	267	211	268	212
rect	273	211	274	212
rect	278	211	279	212
rect	285	211	286	212
rect	296	211	297	212
rect	301	211	302	212
rect	304	211	305	212
rect	307	211	308	212
rect	310	211	311	212
rect	316	211	317	212
rect	319	211	320	212
rect	322	211	323	212
rect	325	211	326	212
rect	328	211	329	212
rect	331	211	332	212
rect	340	211	341	212
rect	343	211	344	212
rect	359	211	360	212
rect	385	211	386	212
rect	394	211	395	212
rect	8	212	9	213
rect	17	212	18	213
rect	24	212	25	213
rect	26	212	27	213
rect	38	212	39	213
rect	42	212	43	213
rect	47	212	48	213
rect	53	212	54	213
rect	56	212	57	213
rect	61	212	62	213
rect	75	212	76	213
rect	98	212	99	213
rect	101	212	102	213
rect	117	212	118	213
rect	126	212	127	213
rect	135	212	136	213
rect	138	212	139	213
rect	147	212	148	213
rect	150	212	151	213
rect	159	212	160	213
rect	168	212	169	213
rect	171	212	172	213
rect	180	212	181	213
rect	186	212	187	213
rect	202	212	203	213
rect	206	212	207	213
rect	208	212	209	213
rect	212	212	213	213
rect	215	212	216	213
rect	224	212	225	213
rect	230	212	231	213
rect	246	212	247	213
rect	249	212	250	213
rect	251	212	252	213
rect	258	212	259	213
rect	261	212	262	213
rect	264	212	265	213
rect	267	212	268	213
rect	273	212	274	213
rect	278	212	279	213
rect	285	212	286	213
rect	296	212	297	213
rect	301	212	302	213
rect	304	212	305	213
rect	307	212	308	213
rect	310	212	311	213
rect	316	212	317	213
rect	319	212	320	213
rect	322	212	323	213
rect	325	212	326	213
rect	328	212	329	213
rect	331	212	332	213
rect	340	212	341	213
rect	343	212	344	213
rect	359	212	360	213
rect	368	212	369	213
rect	385	212	386	213
rect	394	212	395	213
rect	17	213	18	214
rect	24	213	25	214
rect	26	213	27	214
rect	38	213	39	214
rect	42	213	43	214
rect	47	213	48	214
rect	53	213	54	214
rect	56	213	57	214
rect	61	213	62	214
rect	75	213	76	214
rect	98	213	99	214
rect	101	213	102	214
rect	117	213	118	214
rect	126	213	127	214
rect	135	213	136	214
rect	138	213	139	214
rect	147	213	148	214
rect	150	213	151	214
rect	159	213	160	214
rect	168	213	169	214
rect	171	213	172	214
rect	180	213	181	214
rect	186	213	187	214
rect	202	213	203	214
rect	206	213	207	214
rect	208	213	209	214
rect	212	213	213	214
rect	215	213	216	214
rect	224	213	225	214
rect	230	213	231	214
rect	246	213	247	214
rect	249	213	250	214
rect	251	213	252	214
rect	258	213	259	214
rect	261	213	262	214
rect	264	213	265	214
rect	267	213	268	214
rect	273	213	274	214
rect	278	213	279	214
rect	285	213	286	214
rect	296	213	297	214
rect	301	213	302	214
rect	304	213	305	214
rect	307	213	308	214
rect	310	213	311	214
rect	316	213	317	214
rect	319	213	320	214
rect	322	213	323	214
rect	325	213	326	214
rect	328	213	329	214
rect	331	213	332	214
rect	340	213	341	214
rect	343	213	344	214
rect	368	213	369	214
rect	385	213	386	214
rect	17	214	18	215
rect	24	214	25	215
rect	26	214	27	215
rect	38	214	39	215
rect	42	214	43	215
rect	47	214	48	215
rect	53	214	54	215
rect	56	214	57	215
rect	61	214	62	215
rect	75	214	76	215
rect	98	214	99	215
rect	101	214	102	215
rect	117	214	118	215
rect	126	214	127	215
rect	135	214	136	215
rect	138	214	139	215
rect	147	214	148	215
rect	150	214	151	215
rect	159	214	160	215
rect	168	214	169	215
rect	171	214	172	215
rect	180	214	181	215
rect	186	214	187	215
rect	202	214	203	215
rect	206	214	207	215
rect	208	214	209	215
rect	212	214	213	215
rect	215	214	216	215
rect	224	214	225	215
rect	230	214	231	215
rect	246	214	247	215
rect	249	214	250	215
rect	251	214	252	215
rect	258	214	259	215
rect	261	214	262	215
rect	264	214	265	215
rect	267	214	268	215
rect	273	214	274	215
rect	278	214	279	215
rect	285	214	286	215
rect	296	214	297	215
rect	301	214	302	215
rect	304	214	305	215
rect	307	214	308	215
rect	310	214	311	215
rect	316	214	317	215
rect	319	214	320	215
rect	322	214	323	215
rect	325	214	326	215
rect	328	214	329	215
rect	331	214	332	215
rect	340	214	341	215
rect	343	214	344	215
rect	352	214	353	215
rect	368	214	369	215
rect	371	214	372	215
rect	385	214	386	215
rect	387	214	388	215
rect	17	215	18	216
rect	26	215	27	216
rect	38	215	39	216
rect	47	215	48	216
rect	53	215	54	216
rect	56	215	57	216
rect	75	215	76	216
rect	98	215	99	216
rect	101	215	102	216
rect	117	215	118	216
rect	126	215	127	216
rect	135	215	136	216
rect	138	215	139	216
rect	147	215	148	216
rect	150	215	151	216
rect	159	215	160	216
rect	168	215	169	216
rect	180	215	181	216
rect	186	215	187	216
rect	206	215	207	216
rect	212	215	213	216
rect	215	215	216	216
rect	224	215	225	216
rect	246	215	247	216
rect	249	215	250	216
rect	258	215	259	216
rect	261	215	262	216
rect	264	215	265	216
rect	267	215	268	216
rect	273	215	274	216
rect	285	215	286	216
rect	301	215	302	216
rect	304	215	305	216
rect	307	215	308	216
rect	310	215	311	216
rect	316	215	317	216
rect	319	215	320	216
rect	322	215	323	216
rect	325	215	326	216
rect	328	215	329	216
rect	331	215	332	216
rect	340	215	341	216
rect	343	215	344	216
rect	352	215	353	216
rect	368	215	369	216
rect	371	215	372	216
rect	387	215	388	216
rect	8	216	9	217
rect	14	216	15	217
rect	17	216	18	217
rect	26	216	27	217
rect	35	216	36	217
rect	38	216	39	217
rect	47	216	48	217
rect	50	216	51	217
rect	53	216	54	217
rect	56	216	57	217
rect	72	216	73	217
rect	75	216	76	217
rect	81	216	82	217
rect	98	216	99	217
rect	101	216	102	217
rect	117	216	118	217
rect	126	216	127	217
rect	135	216	136	217
rect	138	216	139	217
rect	147	216	148	217
rect	150	216	151	217
rect	159	216	160	217
rect	162	216	163	217
rect	168	216	169	217
rect	177	216	178	217
rect	180	216	181	217
rect	186	216	187	217
rect	203	216	204	217
rect	206	216	207	217
rect	212	216	213	217
rect	215	216	216	217
rect	224	216	225	217
rect	227	216	228	217
rect	243	216	244	217
rect	246	216	247	217
rect	249	216	250	217
rect	258	216	259	217
rect	261	216	262	217
rect	264	216	265	217
rect	267	216	268	217
rect	270	216	271	217
rect	273	216	274	217
rect	282	216	283	217
rect	285	216	286	217
rect	301	216	302	217
rect	304	216	305	217
rect	307	216	308	217
rect	310	216	311	217
rect	316	216	317	217
rect	319	216	320	217
rect	322	216	323	217
rect	325	216	326	217
rect	328	216	329	217
rect	331	216	332	217
rect	340	216	341	217
rect	343	216	344	217
rect	352	216	353	217
rect	368	216	369	217
rect	371	216	372	217
rect	387	216	388	217
rect	14	223	15	224
rect	17	223	18	224
rect	26	223	27	224
rect	35	223	36	224
rect	38	223	39	224
rect	47	223	48	224
rect	50	223	51	224
rect	53	223	54	224
rect	56	223	57	224
rect	66	223	67	224
rect	72	223	73	224
rect	75	223	76	224
rect	92	223	93	224
rect	98	223	99	224
rect	101	223	102	224
rect	117	223	118	224
rect	126	223	127	224
rect	135	223	136	224
rect	138	223	139	224
rect	147	223	148	224
rect	150	223	151	224
rect	159	223	160	224
rect	165	223	166	224
rect	168	223	169	224
rect	177	223	178	224
rect	180	223	181	224
rect	193	223	194	224
rect	203	223	204	224
rect	206	223	207	224
rect	215	223	216	224
rect	221	223	222	224
rect	224	223	225	224
rect	227	223	228	224
rect	240	223	241	224
rect	243	223	244	224
rect	246	223	247	224
rect	249	223	250	224
rect	252	223	253	224
rect	258	223	259	224
rect	261	223	262	224
rect	264	223	265	224
rect	267	223	268	224
rect	270	223	271	224
rect	273	223	274	224
rect	276	223	277	224
rect	282	223	283	224
rect	285	223	286	224
rect	301	223	302	224
rect	304	223	305	224
rect	307	223	308	224
rect	310	223	311	224
rect	316	223	317	224
rect	319	223	320	224
rect	322	223	323	224
rect	325	223	326	224
rect	328	223	329	224
rect	331	223	332	224
rect	334	223	335	224
rect	340	223	341	224
rect	343	223	344	224
rect	346	223	347	224
rect	349	223	350	224
rect	352	223	353	224
rect	362	223	363	224
rect	368	223	369	224
rect	371	223	372	224
rect	381	223	382	224
rect	387	223	388	224
rect	14	224	15	225
rect	17	224	18	225
rect	26	224	27	225
rect	35	224	36	225
rect	38	224	39	225
rect	47	224	48	225
rect	50	224	51	225
rect	53	224	54	225
rect	56	224	57	225
rect	66	224	67	225
rect	72	224	73	225
rect	75	224	76	225
rect	92	224	93	225
rect	98	224	99	225
rect	101	224	102	225
rect	117	224	118	225
rect	126	224	127	225
rect	135	224	136	225
rect	138	224	139	225
rect	147	224	148	225
rect	150	224	151	225
rect	159	224	160	225
rect	165	224	166	225
rect	168	224	169	225
rect	177	224	178	225
rect	180	224	181	225
rect	193	224	194	225
rect	203	224	204	225
rect	206	224	207	225
rect	215	224	216	225
rect	221	224	222	225
rect	224	224	225	225
rect	227	224	228	225
rect	243	224	244	225
rect	246	224	247	225
rect	249	224	250	225
rect	252	224	253	225
rect	258	224	259	225
rect	261	224	262	225
rect	264	224	265	225
rect	270	224	271	225
rect	273	224	274	225
rect	276	224	277	225
rect	282	224	283	225
rect	285	224	286	225
rect	301	224	302	225
rect	304	224	305	225
rect	307	224	308	225
rect	310	224	311	225
rect	316	224	317	225
rect	319	224	320	225
rect	322	224	323	225
rect	325	224	326	225
rect	328	224	329	225
rect	331	224	332	225
rect	334	224	335	225
rect	340	224	341	225
rect	343	224	344	225
rect	346	224	347	225
rect	349	224	350	225
rect	352	224	353	225
rect	362	224	363	225
rect	368	224	369	225
rect	371	224	372	225
rect	381	224	382	225
rect	387	224	388	225
rect	14	225	15	226
rect	17	225	18	226
rect	26	225	27	226
rect	35	225	36	226
rect	38	225	39	226
rect	47	225	48	226
rect	50	225	51	226
rect	53	225	54	226
rect	56	225	57	226
rect	66	225	67	226
rect	72	225	73	226
rect	75	225	76	226
rect	92	225	93	226
rect	98	225	99	226
rect	101	225	102	226
rect	117	225	118	226
rect	126	225	127	226
rect	135	225	136	226
rect	138	225	139	226
rect	147	225	148	226
rect	150	225	151	226
rect	159	225	160	226
rect	165	225	166	226
rect	168	225	169	226
rect	177	225	178	226
rect	180	225	181	226
rect	193	225	194	226
rect	203	225	204	226
rect	206	225	207	226
rect	215	225	216	226
rect	221	225	222	226
rect	224	225	225	226
rect	227	225	228	226
rect	243	225	244	226
rect	246	225	247	226
rect	249	225	250	226
rect	252	225	253	226
rect	258	225	259	226
rect	261	225	262	226
rect	264	225	265	226
rect	270	225	271	226
rect	273	225	274	226
rect	276	225	277	226
rect	282	225	283	226
rect	285	225	286	226
rect	301	225	302	226
rect	304	225	305	226
rect	307	225	308	226
rect	310	225	311	226
rect	316	225	317	226
rect	319	225	320	226
rect	322	225	323	226
rect	325	225	326	226
rect	328	225	329	226
rect	331	225	332	226
rect	334	225	335	226
rect	340	225	341	226
rect	343	225	344	226
rect	346	225	347	226
rect	349	225	350	226
rect	352	225	353	226
rect	362	225	363	226
rect	368	225	369	226
rect	371	225	372	226
rect	381	225	382	226
rect	387	225	388	226
rect	14	226	15	227
rect	17	226	18	227
rect	26	226	27	227
rect	35	226	36	227
rect	38	226	39	227
rect	47	226	48	227
rect	50	226	51	227
rect	53	226	54	227
rect	56	226	57	227
rect	66	226	67	227
rect	72	226	73	227
rect	75	226	76	227
rect	92	226	93	227
rect	98	226	99	227
rect	101	226	102	227
rect	117	226	118	227
rect	126	226	127	227
rect	135	226	136	227
rect	138	226	139	227
rect	147	226	148	227
rect	150	226	151	227
rect	159	226	160	227
rect	165	226	166	227
rect	168	226	169	227
rect	177	226	178	227
rect	180	226	181	227
rect	193	226	194	227
rect	203	226	204	227
rect	206	226	207	227
rect	215	226	216	227
rect	221	226	222	227
rect	224	226	225	227
rect	227	226	228	227
rect	243	226	244	227
rect	246	226	247	227
rect	249	226	250	227
rect	252	226	253	227
rect	258	226	259	227
rect	264	226	265	227
rect	270	226	271	227
rect	273	226	274	227
rect	276	226	277	227
rect	282	226	283	227
rect	285	226	286	227
rect	301	226	302	227
rect	304	226	305	227
rect	307	226	308	227
rect	310	226	311	227
rect	316	226	317	227
rect	319	226	320	227
rect	322	226	323	227
rect	325	226	326	227
rect	328	226	329	227
rect	331	226	332	227
rect	334	226	335	227
rect	340	226	341	227
rect	343	226	344	227
rect	346	226	347	227
rect	349	226	350	227
rect	352	226	353	227
rect	362	226	363	227
rect	368	226	369	227
rect	371	226	372	227
rect	381	226	382	227
rect	387	226	388	227
rect	14	227	15	228
rect	17	227	18	228
rect	26	227	27	228
rect	35	227	36	228
rect	38	227	39	228
rect	47	227	48	228
rect	50	227	51	228
rect	53	227	54	228
rect	56	227	57	228
rect	66	227	67	228
rect	72	227	73	228
rect	75	227	76	228
rect	92	227	93	228
rect	98	227	99	228
rect	101	227	102	228
rect	117	227	118	228
rect	126	227	127	228
rect	135	227	136	228
rect	138	227	139	228
rect	147	227	148	228
rect	150	227	151	228
rect	159	227	160	228
rect	165	227	166	228
rect	168	227	169	228
rect	177	227	178	228
rect	180	227	181	228
rect	193	227	194	228
rect	203	227	204	228
rect	206	227	207	228
rect	215	227	216	228
rect	221	227	222	228
rect	224	227	225	228
rect	227	227	228	228
rect	243	227	244	228
rect	246	227	247	228
rect	249	227	250	228
rect	252	227	253	228
rect	258	227	259	228
rect	264	227	265	228
rect	266	227	267	228
rect	270	227	271	228
rect	273	227	274	228
rect	276	227	277	228
rect	282	227	283	228
rect	285	227	286	228
rect	301	227	302	228
rect	304	227	305	228
rect	307	227	308	228
rect	310	227	311	228
rect	316	227	317	228
rect	319	227	320	228
rect	322	227	323	228
rect	325	227	326	228
rect	328	227	329	228
rect	331	227	332	228
rect	334	227	335	228
rect	340	227	341	228
rect	343	227	344	228
rect	346	227	347	228
rect	349	227	350	228
rect	352	227	353	228
rect	362	227	363	228
rect	368	227	369	228
rect	371	227	372	228
rect	381	227	382	228
rect	387	227	388	228
rect	14	228	15	229
rect	17	228	18	229
rect	26	228	27	229
rect	35	228	36	229
rect	38	228	39	229
rect	47	228	48	229
rect	50	228	51	229
rect	53	228	54	229
rect	56	228	57	229
rect	66	228	67	229
rect	72	228	73	229
rect	75	228	76	229
rect	92	228	93	229
rect	98	228	99	229
rect	101	228	102	229
rect	117	228	118	229
rect	126	228	127	229
rect	135	228	136	229
rect	138	228	139	229
rect	147	228	148	229
rect	150	228	151	229
rect	159	228	160	229
rect	165	228	166	229
rect	168	228	169	229
rect	177	228	178	229
rect	193	228	194	229
rect	203	228	204	229
rect	206	228	207	229
rect	215	228	216	229
rect	221	228	222	229
rect	224	228	225	229
rect	227	228	228	229
rect	243	228	244	229
rect	246	228	247	229
rect	264	228	265	229
rect	266	228	267	229
rect	270	228	271	229
rect	273	228	274	229
rect	282	228	283	229
rect	285	228	286	229
rect	301	228	302	229
rect	304	228	305	229
rect	307	228	308	229
rect	310	228	311	229
rect	316	228	317	229
rect	319	228	320	229
rect	322	228	323	229
rect	325	228	326	229
rect	328	228	329	229
rect	331	228	332	229
rect	334	228	335	229
rect	340	228	341	229
rect	343	228	344	229
rect	346	228	347	229
rect	349	228	350	229
rect	352	228	353	229
rect	362	228	363	229
rect	368	228	369	229
rect	371	228	372	229
rect	381	228	382	229
rect	387	228	388	229
rect	14	229	15	230
rect	17	229	18	230
rect	26	229	27	230
rect	35	229	36	230
rect	38	229	39	230
rect	47	229	48	230
rect	50	229	51	230
rect	53	229	54	230
rect	56	229	57	230
rect	66	229	67	230
rect	72	229	73	230
rect	75	229	76	230
rect	92	229	93	230
rect	98	229	99	230
rect	101	229	102	230
rect	117	229	118	230
rect	126	229	127	230
rect	135	229	136	230
rect	138	229	139	230
rect	147	229	148	230
rect	150	229	151	230
rect	159	229	160	230
rect	165	229	166	230
rect	168	229	169	230
rect	177	229	178	230
rect	188	229	189	230
rect	193	229	194	230
rect	203	229	204	230
rect	206	229	207	230
rect	215	229	216	230
rect	221	229	222	230
rect	224	229	225	230
rect	227	229	228	230
rect	243	229	244	230
rect	246	229	247	230
rect	264	229	265	230
rect	266	229	267	230
rect	270	229	271	230
rect	273	229	274	230
rect	282	229	283	230
rect	285	229	286	230
rect	301	229	302	230
rect	304	229	305	230
rect	307	229	308	230
rect	310	229	311	230
rect	316	229	317	230
rect	319	229	320	230
rect	322	229	323	230
rect	325	229	326	230
rect	328	229	329	230
rect	331	229	332	230
rect	334	229	335	230
rect	340	229	341	230
rect	343	229	344	230
rect	346	229	347	230
rect	349	229	350	230
rect	352	229	353	230
rect	362	229	363	230
rect	368	229	369	230
rect	371	229	372	230
rect	381	229	382	230
rect	387	229	388	230
rect	14	230	15	231
rect	17	230	18	231
rect	26	230	27	231
rect	35	230	36	231
rect	38	230	39	231
rect	47	230	48	231
rect	50	230	51	231
rect	53	230	54	231
rect	56	230	57	231
rect	66	230	67	231
rect	72	230	73	231
rect	75	230	76	231
rect	92	230	93	231
rect	98	230	99	231
rect	101	230	102	231
rect	117	230	118	231
rect	126	230	127	231
rect	135	230	136	231
rect	147	230	148	231
rect	159	230	160	231
rect	165	230	166	231
rect	168	230	169	231
rect	188	230	189	231
rect	193	230	194	231
rect	203	230	204	231
rect	206	230	207	231
rect	215	230	216	231
rect	227	230	228	231
rect	243	230	244	231
rect	246	230	247	231
rect	264	230	265	231
rect	266	230	267	231
rect	270	230	271	231
rect	282	230	283	231
rect	285	230	286	231
rect	301	230	302	231
rect	304	230	305	231
rect	307	230	308	231
rect	310	230	311	231
rect	316	230	317	231
rect	319	230	320	231
rect	322	230	323	231
rect	325	230	326	231
rect	328	230	329	231
rect	331	230	332	231
rect	334	230	335	231
rect	340	230	341	231
rect	343	230	344	231
rect	346	230	347	231
rect	349	230	350	231
rect	352	230	353	231
rect	362	230	363	231
rect	368	230	369	231
rect	371	230	372	231
rect	381	230	382	231
rect	387	230	388	231
rect	14	231	15	232
rect	17	231	18	232
rect	26	231	27	232
rect	35	231	36	232
rect	38	231	39	232
rect	47	231	48	232
rect	50	231	51	232
rect	53	231	54	232
rect	56	231	57	232
rect	66	231	67	232
rect	72	231	73	232
rect	75	231	76	232
rect	92	231	93	232
rect	98	231	99	232
rect	101	231	102	232
rect	117	231	118	232
rect	126	231	127	232
rect	135	231	136	232
rect	137	231	138	232
rect	147	231	148	232
rect	159	231	160	232
rect	161	231	162	232
rect	165	231	166	232
rect	168	231	169	232
rect	185	231	186	232
rect	188	231	189	232
rect	193	231	194	232
rect	203	231	204	232
rect	206	231	207	232
rect	215	231	216	232
rect	227	231	228	232
rect	243	231	244	232
rect	246	231	247	232
rect	248	231	249	232
rect	260	231	261	232
rect	264	231	265	232
rect	266	231	267	232
rect	270	231	271	232
rect	275	231	276	232
rect	282	231	283	232
rect	285	231	286	232
rect	301	231	302	232
rect	304	231	305	232
rect	307	231	308	232
rect	310	231	311	232
rect	316	231	317	232
rect	319	231	320	232
rect	322	231	323	232
rect	325	231	326	232
rect	328	231	329	232
rect	331	231	332	232
rect	334	231	335	232
rect	340	231	341	232
rect	343	231	344	232
rect	346	231	347	232
rect	349	231	350	232
rect	352	231	353	232
rect	362	231	363	232
rect	368	231	369	232
rect	371	231	372	232
rect	381	231	382	232
rect	387	231	388	232
rect	14	232	15	233
rect	17	232	18	233
rect	26	232	27	233
rect	35	232	36	233
rect	38	232	39	233
rect	47	232	48	233
rect	50	232	51	233
rect	53	232	54	233
rect	66	232	67	233
rect	72	232	73	233
rect	75	232	76	233
rect	92	232	93	233
rect	98	232	99	233
rect	101	232	102	233
rect	117	232	118	233
rect	126	232	127	233
rect	137	232	138	233
rect	147	232	148	233
rect	159	232	160	233
rect	161	232	162	233
rect	165	232	166	233
rect	168	232	169	233
rect	185	232	186	233
rect	188	232	189	233
rect	193	232	194	233
rect	206	232	207	233
rect	227	232	228	233
rect	243	232	244	233
rect	248	232	249	233
rect	260	232	261	233
rect	264	232	265	233
rect	266	232	267	233
rect	270	232	271	233
rect	275	232	276	233
rect	282	232	283	233
rect	285	232	286	233
rect	301	232	302	233
rect	304	232	305	233
rect	307	232	308	233
rect	310	232	311	233
rect	316	232	317	233
rect	319	232	320	233
rect	322	232	323	233
rect	325	232	326	233
rect	328	232	329	233
rect	331	232	332	233
rect	334	232	335	233
rect	340	232	341	233
rect	343	232	344	233
rect	346	232	347	233
rect	349	232	350	233
rect	352	232	353	233
rect	362	232	363	233
rect	368	232	369	233
rect	371	232	372	233
rect	381	232	382	233
rect	387	232	388	233
rect	14	233	15	234
rect	17	233	18	234
rect	26	233	27	234
rect	35	233	36	234
rect	38	233	39	234
rect	47	233	48	234
rect	50	233	51	234
rect	53	233	54	234
rect	60	233	61	234
rect	66	233	67	234
rect	72	233	73	234
rect	75	233	76	234
rect	92	233	93	234
rect	98	233	99	234
rect	101	233	102	234
rect	117	233	118	234
rect	126	233	127	234
rect	137	233	138	234
rect	147	233	148	234
rect	149	233	150	234
rect	159	233	160	234
rect	161	233	162	234
rect	165	233	166	234
rect	168	233	169	234
rect	170	233	171	234
rect	179	233	180	234
rect	185	233	186	234
rect	188	233	189	234
rect	193	233	194	234
rect	206	233	207	234
rect	210	233	211	234
rect	227	233	228	234
rect	232	233	233	234
rect	243	233	244	234
rect	248	233	249	234
rect	260	233	261	234
rect	264	233	265	234
rect	266	233	267	234
rect	270	233	271	234
rect	272	233	273	234
rect	275	233	276	234
rect	282	233	283	234
rect	285	233	286	234
rect	301	233	302	234
rect	304	233	305	234
rect	307	233	308	234
rect	310	233	311	234
rect	316	233	317	234
rect	319	233	320	234
rect	322	233	323	234
rect	325	233	326	234
rect	328	233	329	234
rect	331	233	332	234
rect	334	233	335	234
rect	340	233	341	234
rect	343	233	344	234
rect	346	233	347	234
rect	349	233	350	234
rect	352	233	353	234
rect	362	233	363	234
rect	368	233	369	234
rect	371	233	372	234
rect	381	233	382	234
rect	387	233	388	234
rect	14	234	15	235
rect	17	234	18	235
rect	26	234	27	235
rect	35	234	36	235
rect	38	234	39	235
rect	47	234	48	235
rect	50	234	51	235
rect	60	234	61	235
rect	66	234	67	235
rect	72	234	73	235
rect	75	234	76	235
rect	92	234	93	235
rect	98	234	99	235
rect	117	234	118	235
rect	126	234	127	235
rect	137	234	138	235
rect	149	234	150	235
rect	159	234	160	235
rect	161	234	162	235
rect	165	234	166	235
rect	170	234	171	235
rect	179	234	180	235
rect	185	234	186	235
rect	188	234	189	235
rect	193	234	194	235
rect	210	234	211	235
rect	227	234	228	235
rect	232	234	233	235
rect	248	234	249	235
rect	260	234	261	235
rect	264	234	265	235
rect	266	234	267	235
rect	270	234	271	235
rect	272	234	273	235
rect	275	234	276	235
rect	282	234	283	235
rect	285	234	286	235
rect	301	234	302	235
rect	304	234	305	235
rect	307	234	308	235
rect	310	234	311	235
rect	316	234	317	235
rect	319	234	320	235
rect	322	234	323	235
rect	328	234	329	235
rect	331	234	332	235
rect	334	234	335	235
rect	340	234	341	235
rect	343	234	344	235
rect	346	234	347	235
rect	349	234	350	235
rect	352	234	353	235
rect	362	234	363	235
rect	368	234	369	235
rect	371	234	372	235
rect	381	234	382	235
rect	387	234	388	235
rect	14	235	15	236
rect	17	235	18	236
rect	26	235	27	236
rect	35	235	36	236
rect	38	235	39	236
rect	47	235	48	236
rect	50	235	51	236
rect	57	235	58	236
rect	60	235	61	236
rect	66	235	67	236
rect	72	235	73	236
rect	75	235	76	236
rect	92	235	93	236
rect	98	235	99	236
rect	106	235	107	236
rect	117	235	118	236
rect	126	235	127	236
rect	134	235	135	236
rect	137	235	138	236
rect	149	235	150	236
rect	159	235	160	236
rect	161	235	162	236
rect	165	235	166	236
rect	170	235	171	236
rect	176	235	177	236
rect	179	235	180	236
rect	185	235	186	236
rect	188	235	189	236
rect	193	235	194	236
rect	197	235	198	236
rect	210	235	211	236
rect	214	235	215	236
rect	220	235	221	236
rect	227	235	228	236
rect	232	235	233	236
rect	248	235	249	236
rect	251	235	252	236
rect	260	235	261	236
rect	264	235	265	236
rect	266	235	267	236
rect	270	235	271	236
rect	272	235	273	236
rect	275	235	276	236
rect	282	235	283	236
rect	285	235	286	236
rect	301	235	302	236
rect	304	235	305	236
rect	307	235	308	236
rect	310	235	311	236
rect	316	235	317	236
rect	319	235	320	236
rect	322	235	323	236
rect	328	235	329	236
rect	331	235	332	236
rect	334	235	335	236
rect	336	235	337	236
rect	340	235	341	236
rect	343	235	344	236
rect	346	235	347	236
rect	349	235	350	236
rect	352	235	353	236
rect	362	235	363	236
rect	368	235	369	236
rect	371	235	372	236
rect	381	235	382	236
rect	387	235	388	236
rect	14	236	15	237
rect	17	236	18	237
rect	26	236	27	237
rect	35	236	36	237
rect	38	236	39	237
rect	47	236	48	237
rect	57	236	58	237
rect	60	236	61	237
rect	66	236	67	237
rect	72	236	73	237
rect	75	236	76	237
rect	92	236	93	237
rect	106	236	107	237
rect	134	236	135	237
rect	137	236	138	237
rect	149	236	150	237
rect	161	236	162	237
rect	165	236	166	237
rect	170	236	171	237
rect	176	236	177	237
rect	179	236	180	237
rect	185	236	186	237
rect	188	236	189	237
rect	197	236	198	237
rect	210	236	211	237
rect	214	236	215	237
rect	220	236	221	237
rect	227	236	228	237
rect	232	236	233	237
rect	248	236	249	237
rect	251	236	252	237
rect	260	236	261	237
rect	264	236	265	237
rect	266	236	267	237
rect	270	236	271	237
rect	272	236	273	237
rect	275	236	276	237
rect	282	236	283	237
rect	301	236	302	237
rect	304	236	305	237
rect	307	236	308	237
rect	310	236	311	237
rect	316	236	317	237
rect	322	236	323	237
rect	328	236	329	237
rect	331	236	332	237
rect	336	236	337	237
rect	343	236	344	237
rect	349	236	350	237
rect	352	236	353	237
rect	362	236	363	237
rect	368	236	369	237
rect	371	236	372	237
rect	381	236	382	237
rect	387	236	388	237
rect	14	237	15	238
rect	17	237	18	238
rect	26	237	27	238
rect	35	237	36	238
rect	38	237	39	238
rect	47	237	48	238
rect	54	237	55	238
rect	57	237	58	238
rect	60	237	61	238
rect	66	237	67	238
rect	72	237	73	238
rect	75	237	76	238
rect	92	237	93	238
rect	106	237	107	238
rect	109	237	110	238
rect	118	237	119	238
rect	134	237	135	238
rect	137	237	138	238
rect	140	237	141	238
rect	149	237	150	238
rect	161	237	162	238
rect	165	237	166	238
rect	170	237	171	238
rect	173	237	174	238
rect	176	237	177	238
rect	179	237	180	238
rect	185	237	186	238
rect	188	237	189	238
rect	197	237	198	238
rect	210	237	211	238
rect	214	237	215	238
rect	220	237	221	238
rect	227	237	228	238
rect	232	237	233	238
rect	248	237	249	238
rect	251	237	252	238
rect	260	237	261	238
rect	264	237	265	238
rect	266	237	267	238
rect	270	237	271	238
rect	272	237	273	238
rect	275	237	276	238
rect	282	237	283	238
rect	301	237	302	238
rect	304	237	305	238
rect	307	237	308	238
rect	310	237	311	238
rect	316	237	317	238
rect	322	237	323	238
rect	328	237	329	238
rect	331	237	332	238
rect	336	237	337	238
rect	343	237	344	238
rect	349	237	350	238
rect	352	237	353	238
rect	362	237	363	238
rect	368	237	369	238
rect	371	237	372	238
rect	381	237	382	238
rect	387	237	388	238
rect	14	238	15	239
rect	17	238	18	239
rect	26	238	27	239
rect	35	238	36	239
rect	38	238	39	239
rect	54	238	55	239
rect	57	238	58	239
rect	60	238	61	239
rect	66	238	67	239
rect	72	238	73	239
rect	75	238	76	239
rect	92	238	93	239
rect	106	238	107	239
rect	109	238	110	239
rect	118	238	119	239
rect	134	238	135	239
rect	137	238	138	239
rect	140	238	141	239
rect	149	238	150	239
rect	161	238	162	239
rect	170	238	171	239
rect	173	238	174	239
rect	176	238	177	239
rect	179	238	180	239
rect	185	238	186	239
rect	188	238	189	239
rect	197	238	198	239
rect	210	238	211	239
rect	214	238	215	239
rect	220	238	221	239
rect	227	238	228	239
rect	232	238	233	239
rect	248	238	249	239
rect	251	238	252	239
rect	260	238	261	239
rect	264	238	265	239
rect	266	238	267	239
rect	270	238	271	239
rect	272	238	273	239
rect	275	238	276	239
rect	282	238	283	239
rect	301	238	302	239
rect	304	238	305	239
rect	307	238	308	239
rect	310	238	311	239
rect	316	238	317	239
rect	322	238	323	239
rect	331	238	332	239
rect	336	238	337	239
rect	343	238	344	239
rect	349	238	350	239
rect	352	238	353	239
rect	362	238	363	239
rect	368	238	369	239
rect	371	238	372	239
rect	381	238	382	239
rect	387	238	388	239
rect	14	239	15	240
rect	17	239	18	240
rect	26	239	27	240
rect	35	239	36	240
rect	38	239	39	240
rect	51	239	52	240
rect	54	239	55	240
rect	57	239	58	240
rect	60	239	61	240
rect	66	239	67	240
rect	72	239	73	240
rect	75	239	76	240
rect	80	239	81	240
rect	92	239	93	240
rect	106	239	107	240
rect	109	239	110	240
rect	118	239	119	240
rect	134	239	135	240
rect	137	239	138	240
rect	140	239	141	240
rect	149	239	150	240
rect	158	239	159	240
rect	161	239	162	240
rect	170	239	171	240
rect	173	239	174	240
rect	176	239	177	240
rect	179	239	180	240
rect	185	239	186	240
rect	188	239	189	240
rect	197	239	198	240
rect	210	239	211	240
rect	214	239	215	240
rect	220	239	221	240
rect	227	239	228	240
rect	232	239	233	240
rect	248	239	249	240
rect	251	239	252	240
rect	260	239	261	240
rect	264	239	265	240
rect	266	239	267	240
rect	270	239	271	240
rect	272	239	273	240
rect	275	239	276	240
rect	282	239	283	240
rect	301	239	302	240
rect	304	239	305	240
rect	307	239	308	240
rect	310	239	311	240
rect	316	239	317	240
rect	322	239	323	240
rect	324	239	325	240
rect	331	239	332	240
rect	336	239	337	240
rect	339	239	340	240
rect	343	239	344	240
rect	349	239	350	240
rect	352	239	353	240
rect	362	239	363	240
rect	368	239	369	240
rect	371	239	372	240
rect	381	239	382	240
rect	387	239	388	240
rect	14	240	15	241
rect	17	240	18	241
rect	38	240	39	241
rect	51	240	52	241
rect	54	240	55	241
rect	57	240	58	241
rect	60	240	61	241
rect	66	240	67	241
rect	72	240	73	241
rect	80	240	81	241
rect	92	240	93	241
rect	106	240	107	241
rect	109	240	110	241
rect	118	240	119	241
rect	134	240	135	241
rect	137	240	138	241
rect	140	240	141	241
rect	149	240	150	241
rect	158	240	159	241
rect	161	240	162	241
rect	170	240	171	241
rect	173	240	174	241
rect	176	240	177	241
rect	179	240	180	241
rect	185	240	186	241
rect	188	240	189	241
rect	197	240	198	241
rect	210	240	211	241
rect	214	240	215	241
rect	220	240	221	241
rect	227	240	228	241
rect	232	240	233	241
rect	248	240	249	241
rect	251	240	252	241
rect	260	240	261	241
rect	264	240	265	241
rect	266	240	267	241
rect	270	240	271	241
rect	272	240	273	241
rect	275	240	276	241
rect	282	240	283	241
rect	301	240	302	241
rect	304	240	305	241
rect	307	240	308	241
rect	310	240	311	241
rect	316	240	317	241
rect	322	240	323	241
rect	324	240	325	241
rect	336	240	337	241
rect	339	240	340	241
rect	343	240	344	241
rect	349	240	350	241
rect	352	240	353	241
rect	368	240	369	241
rect	371	240	372	241
rect	381	240	382	241
rect	387	240	388	241
rect	14	241	15	242
rect	17	241	18	242
rect	24	241	25	242
rect	38	241	39	242
rect	48	241	49	242
rect	51	241	52	242
rect	54	241	55	242
rect	57	241	58	242
rect	60	241	61	242
rect	66	241	67	242
rect	72	241	73	242
rect	80	241	81	242
rect	92	241	93	242
rect	106	241	107	242
rect	109	241	110	242
rect	118	241	119	242
rect	134	241	135	242
rect	137	241	138	242
rect	140	241	141	242
rect	149	241	150	242
rect	158	241	159	242
rect	161	241	162	242
rect	170	241	171	242
rect	173	241	174	242
rect	176	241	177	242
rect	179	241	180	242
rect	185	241	186	242
rect	188	241	189	242
rect	197	241	198	242
rect	210	241	211	242
rect	214	241	215	242
rect	220	241	221	242
rect	227	241	228	242
rect	232	241	233	242
rect	248	241	249	242
rect	251	241	252	242
rect	260	241	261	242
rect	264	241	265	242
rect	266	241	267	242
rect	270	241	271	242
rect	272	241	273	242
rect	275	241	276	242
rect	282	241	283	242
rect	301	241	302	242
rect	304	241	305	242
rect	307	241	308	242
rect	310	241	311	242
rect	316	241	317	242
rect	322	241	323	242
rect	324	241	325	242
rect	327	241	328	242
rect	336	241	337	242
rect	339	241	340	242
rect	343	241	344	242
rect	349	241	350	242
rect	352	241	353	242
rect	368	241	369	242
rect	371	241	372	242
rect	381	241	382	242
rect	387	241	388	242
rect	14	242	15	243
rect	24	242	25	243
rect	48	242	49	243
rect	51	242	52	243
rect	54	242	55	243
rect	57	242	58	243
rect	60	242	61	243
rect	66	242	67	243
rect	80	242	81	243
rect	106	242	107	243
rect	109	242	110	243
rect	118	242	119	243
rect	134	242	135	243
rect	137	242	138	243
rect	140	242	141	243
rect	149	242	150	243
rect	158	242	159	243
rect	161	242	162	243
rect	170	242	171	243
rect	173	242	174	243
rect	176	242	177	243
rect	179	242	180	243
rect	185	242	186	243
rect	188	242	189	243
rect	197	242	198	243
rect	210	242	211	243
rect	214	242	215	243
rect	220	242	221	243
rect	227	242	228	243
rect	232	242	233	243
rect	248	242	249	243
rect	251	242	252	243
rect	260	242	261	243
rect	264	242	265	243
rect	266	242	267	243
rect	270	242	271	243
rect	272	242	273	243
rect	275	242	276	243
rect	282	242	283	243
rect	301	242	302	243
rect	304	242	305	243
rect	307	242	308	243
rect	310	242	311	243
rect	316	242	317	243
rect	322	242	323	243
rect	324	242	325	243
rect	327	242	328	243
rect	336	242	337	243
rect	339	242	340	243
rect	352	242	353	243
rect	381	242	382	243
rect	387	242	388	243
rect	14	243	15	244
rect	24	243	25	244
rect	27	243	28	244
rect	30	243	31	244
rect	48	243	49	244
rect	51	243	52	244
rect	54	243	55	244
rect	57	243	58	244
rect	60	243	61	244
rect	66	243	67	244
rect	80	243	81	244
rect	83	243	84	244
rect	106	243	107	244
rect	109	243	110	244
rect	118	243	119	244
rect	134	243	135	244
rect	137	243	138	244
rect	140	243	141	244
rect	149	243	150	244
rect	158	243	159	244
rect	161	243	162	244
rect	170	243	171	244
rect	173	243	174	244
rect	176	243	177	244
rect	179	243	180	244
rect	185	243	186	244
rect	188	243	189	244
rect	197	243	198	244
rect	210	243	211	244
rect	214	243	215	244
rect	220	243	221	244
rect	227	243	228	244
rect	232	243	233	244
rect	248	243	249	244
rect	251	243	252	244
rect	260	243	261	244
rect	264	243	265	244
rect	266	243	267	244
rect	270	243	271	244
rect	272	243	273	244
rect	275	243	276	244
rect	282	243	283	244
rect	301	243	302	244
rect	304	243	305	244
rect	307	243	308	244
rect	310	243	311	244
rect	316	243	317	244
rect	322	243	323	244
rect	324	243	325	244
rect	327	243	328	244
rect	333	243	334	244
rect	336	243	337	244
rect	339	243	340	244
rect	352	243	353	244
rect	360	243	361	244
rect	376	243	377	244
rect	381	243	382	244
rect	387	243	388	244
rect	24	244	25	245
rect	27	244	28	245
rect	30	244	31	245
rect	48	244	49	245
rect	51	244	52	245
rect	54	244	55	245
rect	57	244	58	245
rect	60	244	61	245
rect	80	244	81	245
rect	83	244	84	245
rect	106	244	107	245
rect	109	244	110	245
rect	118	244	119	245
rect	134	244	135	245
rect	137	244	138	245
rect	140	244	141	245
rect	149	244	150	245
rect	158	244	159	245
rect	161	244	162	245
rect	170	244	171	245
rect	173	244	174	245
rect	176	244	177	245
rect	179	244	180	245
rect	185	244	186	245
rect	188	244	189	245
rect	197	244	198	245
rect	210	244	211	245
rect	214	244	215	245
rect	220	244	221	245
rect	232	244	233	245
rect	248	244	249	245
rect	251	244	252	245
rect	260	244	261	245
rect	264	244	265	245
rect	266	244	267	245
rect	272	244	273	245
rect	275	244	276	245
rect	282	244	283	245
rect	301	244	302	245
rect	304	244	305	245
rect	310	244	311	245
rect	322	244	323	245
rect	324	244	325	245
rect	327	244	328	245
rect	333	244	334	245
rect	336	244	337	245
rect	339	244	340	245
rect	352	244	353	245
rect	360	244	361	245
rect	376	244	377	245
rect	387	244	388	245
rect	21	245	22	246
rect	24	245	25	246
rect	27	245	28	246
rect	30	245	31	246
rect	36	245	37	246
rect	39	245	40	246
rect	48	245	49	246
rect	51	245	52	246
rect	54	245	55	246
rect	57	245	58	246
rect	60	245	61	246
rect	80	245	81	246
rect	83	245	84	246
rect	106	245	107	246
rect	109	245	110	246
rect	118	245	119	246
rect	134	245	135	246
rect	137	245	138	246
rect	140	245	141	246
rect	149	245	150	246
rect	158	245	159	246
rect	161	245	162	246
rect	170	245	171	246
rect	173	245	174	246
rect	176	245	177	246
rect	179	245	180	246
rect	185	245	186	246
rect	188	245	189	246
rect	197	245	198	246
rect	210	245	211	246
rect	214	245	215	246
rect	220	245	221	246
rect	223	245	224	246
rect	232	245	233	246
rect	248	245	249	246
rect	251	245	252	246
rect	254	245	255	246
rect	260	245	261	246
rect	264	245	265	246
rect	266	245	267	246
rect	272	245	273	246
rect	275	245	276	246
rect	282	245	283	246
rect	287	245	288	246
rect	301	245	302	246
rect	304	245	305	246
rect	308	245	309	246
rect	310	245	311	246
rect	322	245	323	246
rect	324	245	325	246
rect	327	245	328	246
rect	333	245	334	246
rect	336	245	337	246
rect	339	245	340	246
rect	352	245	353	246
rect	360	245	361	246
rect	376	245	377	246
rect	387	245	388	246
rect	21	246	22	247
rect	24	246	25	247
rect	27	246	28	247
rect	30	246	31	247
rect	36	246	37	247
rect	39	246	40	247
rect	48	246	49	247
rect	51	246	52	247
rect	54	246	55	247
rect	57	246	58	247
rect	60	246	61	247
rect	80	246	81	247
rect	83	246	84	247
rect	106	246	107	247
rect	109	246	110	247
rect	118	246	119	247
rect	134	246	135	247
rect	137	246	138	247
rect	140	246	141	247
rect	149	246	150	247
rect	158	246	159	247
rect	161	246	162	247
rect	170	246	171	247
rect	173	246	174	247
rect	176	246	177	247
rect	179	246	180	247
rect	185	246	186	247
rect	188	246	189	247
rect	197	246	198	247
rect	210	246	211	247
rect	214	246	215	247
rect	220	246	221	247
rect	223	246	224	247
rect	232	246	233	247
rect	248	246	249	247
rect	251	246	252	247
rect	254	246	255	247
rect	260	246	261	247
rect	266	246	267	247
rect	272	246	273	247
rect	275	246	276	247
rect	287	246	288	247
rect	308	246	309	247
rect	324	246	325	247
rect	327	246	328	247
rect	333	246	334	247
rect	336	246	337	247
rect	339	246	340	247
rect	360	246	361	247
rect	376	246	377	247
rect	4	247	5	248
rect	21	247	22	248
rect	24	247	25	248
rect	27	247	28	248
rect	30	247	31	248
rect	36	247	37	248
rect	39	247	40	248
rect	48	247	49	248
rect	51	247	52	248
rect	54	247	55	248
rect	57	247	58	248
rect	60	247	61	248
rect	80	247	81	248
rect	83	247	84	248
rect	106	247	107	248
rect	109	247	110	248
rect	118	247	119	248
rect	134	247	135	248
rect	137	247	138	248
rect	140	247	141	248
rect	149	247	150	248
rect	158	247	159	248
rect	161	247	162	248
rect	170	247	171	248
rect	173	247	174	248
rect	176	247	177	248
rect	179	247	180	248
rect	185	247	186	248
rect	188	247	189	248
rect	197	247	198	248
rect	210	247	211	248
rect	214	247	215	248
rect	220	247	221	248
rect	223	247	224	248
rect	232	247	233	248
rect	248	247	249	248
rect	251	247	252	248
rect	254	247	255	248
rect	257	247	258	248
rect	260	247	261	248
rect	266	247	267	248
rect	269	247	270	248
rect	272	247	273	248
rect	275	247	276	248
rect	284	247	285	248
rect	287	247	288	248
rect	296	247	297	248
rect	305	247	306	248
rect	308	247	309	248
rect	324	247	325	248
rect	327	247	328	248
rect	333	247	334	248
rect	336	247	337	248
rect	339	247	340	248
rect	348	247	349	248
rect	357	247	358	248
rect	360	247	361	248
rect	363	247	364	248
rect	370	247	371	248
rect	373	247	374	248
rect	376	247	377	248
rect	379	247	380	248
rect	4	254	5	255
rect	21	254	22	255
rect	24	254	25	255
rect	27	254	28	255
rect	30	254	31	255
rect	39	254	40	255
rect	48	254	49	255
rect	51	254	52	255
rect	54	254	55	255
rect	57	254	58	255
rect	60	254	61	255
rect	83	254	84	255
rect	89	254	90	255
rect	103	254	104	255
rect	106	254	107	255
rect	109	254	110	255
rect	112	254	113	255
rect	118	254	119	255
rect	134	254	135	255
rect	137	254	138	255
rect	140	254	141	255
rect	149	254	150	255
rect	158	254	159	255
rect	161	254	162	255
rect	164	254	165	255
rect	170	254	171	255
rect	173	254	174	255
rect	176	254	177	255
rect	179	254	180	255
rect	185	254	186	255
rect	188	254	189	255
rect	194	254	195	255
rect	197	254	198	255
rect	220	254	221	255
rect	223	254	224	255
rect	232	254	233	255
rect	248	254	249	255
rect	251	254	252	255
rect	254	254	255	255
rect	257	254	258	255
rect	266	254	267	255
rect	269	254	270	255
rect	272	254	273	255
rect	275	254	276	255
rect	281	254	282	255
rect	284	254	285	255
rect	287	254	288	255
rect	296	254	297	255
rect	305	254	306	255
rect	308	254	309	255
rect	314	254	315	255
rect	324	254	325	255
rect	333	254	334	255
rect	336	254	337	255
rect	339	254	340	255
rect	348	254	349	255
rect	357	254	358	255
rect	373	254	374	255
rect	376	254	377	255
rect	379	254	380	255
rect	4	255	5	256
rect	21	255	22	256
rect	24	255	25	256
rect	27	255	28	256
rect	30	255	31	256
rect	39	255	40	256
rect	48	255	49	256
rect	51	255	52	256
rect	54	255	55	256
rect	57	255	58	256
rect	60	255	61	256
rect	83	255	84	256
rect	89	255	90	256
rect	103	255	104	256
rect	106	255	107	256
rect	109	255	110	256
rect	112	255	113	256
rect	118	255	119	256
rect	134	255	135	256
rect	137	255	138	256
rect	140	255	141	256
rect	149	255	150	256
rect	158	255	159	256
rect	161	255	162	256
rect	164	255	165	256
rect	170	255	171	256
rect	173	255	174	256
rect	176	255	177	256
rect	179	255	180	256
rect	185	255	186	256
rect	188	255	189	256
rect	194	255	195	256
rect	197	255	198	256
rect	220	255	221	256
rect	223	255	224	256
rect	232	255	233	256
rect	248	255	249	256
rect	251	255	252	256
rect	254	255	255	256
rect	257	255	258	256
rect	266	255	267	256
rect	269	255	270	256
rect	272	255	273	256
rect	275	255	276	256
rect	284	255	285	256
rect	287	255	288	256
rect	296	255	297	256
rect	305	255	306	256
rect	308	255	309	256
rect	314	255	315	256
rect	324	255	325	256
rect	333	255	334	256
rect	336	255	337	256
rect	339	255	340	256
rect	348	255	349	256
rect	357	255	358	256
rect	373	255	374	256
rect	376	255	377	256
rect	379	255	380	256
rect	4	256	5	257
rect	21	256	22	257
rect	24	256	25	257
rect	27	256	28	257
rect	30	256	31	257
rect	39	256	40	257
rect	48	256	49	257
rect	51	256	52	257
rect	54	256	55	257
rect	57	256	58	257
rect	60	256	61	257
rect	83	256	84	257
rect	89	256	90	257
rect	103	256	104	257
rect	106	256	107	257
rect	109	256	110	257
rect	112	256	113	257
rect	118	256	119	257
rect	134	256	135	257
rect	137	256	138	257
rect	140	256	141	257
rect	149	256	150	257
rect	158	256	159	257
rect	161	256	162	257
rect	164	256	165	257
rect	170	256	171	257
rect	173	256	174	257
rect	176	256	177	257
rect	179	256	180	257
rect	185	256	186	257
rect	188	256	189	257
rect	194	256	195	257
rect	197	256	198	257
rect	220	256	221	257
rect	223	256	224	257
rect	232	256	233	257
rect	248	256	249	257
rect	251	256	252	257
rect	254	256	255	257
rect	257	256	258	257
rect	266	256	267	257
rect	269	256	270	257
rect	272	256	273	257
rect	275	256	276	257
rect	284	256	285	257
rect	287	256	288	257
rect	296	256	297	257
rect	305	256	306	257
rect	308	256	309	257
rect	314	256	315	257
rect	324	256	325	257
rect	333	256	334	257
rect	336	256	337	257
rect	339	256	340	257
rect	348	256	349	257
rect	357	256	358	257
rect	366	256	367	257
rect	373	256	374	257
rect	376	256	377	257
rect	379	256	380	257
rect	4	257	5	258
rect	21	257	22	258
rect	24	257	25	258
rect	27	257	28	258
rect	30	257	31	258
rect	39	257	40	258
rect	48	257	49	258
rect	51	257	52	258
rect	54	257	55	258
rect	57	257	58	258
rect	60	257	61	258
rect	83	257	84	258
rect	89	257	90	258
rect	103	257	104	258
rect	106	257	107	258
rect	109	257	110	258
rect	112	257	113	258
rect	118	257	119	258
rect	134	257	135	258
rect	137	257	138	258
rect	140	257	141	258
rect	149	257	150	258
rect	158	257	159	258
rect	161	257	162	258
rect	164	257	165	258
rect	170	257	171	258
rect	173	257	174	258
rect	176	257	177	258
rect	188	257	189	258
rect	194	257	195	258
rect	197	257	198	258
rect	220	257	221	258
rect	223	257	224	258
rect	232	257	233	258
rect	248	257	249	258
rect	251	257	252	258
rect	254	257	255	258
rect	257	257	258	258
rect	266	257	267	258
rect	269	257	270	258
rect	272	257	273	258
rect	284	257	285	258
rect	287	257	288	258
rect	296	257	297	258
rect	305	257	306	258
rect	308	257	309	258
rect	314	257	315	258
rect	324	257	325	258
rect	333	257	334	258
rect	336	257	337	258
rect	339	257	340	258
rect	348	257	349	258
rect	357	257	358	258
rect	366	257	367	258
rect	373	257	374	258
rect	376	257	377	258
rect	379	257	380	258
rect	4	258	5	259
rect	21	258	22	259
rect	24	258	25	259
rect	27	258	28	259
rect	30	258	31	259
rect	39	258	40	259
rect	48	258	49	259
rect	51	258	52	259
rect	54	258	55	259
rect	57	258	58	259
rect	60	258	61	259
rect	83	258	84	259
rect	89	258	90	259
rect	103	258	104	259
rect	106	258	107	259
rect	109	258	110	259
rect	112	258	113	259
rect	118	258	119	259
rect	134	258	135	259
rect	137	258	138	259
rect	140	258	141	259
rect	149	258	150	259
rect	158	258	159	259
rect	161	258	162	259
rect	164	258	165	259
rect	170	258	171	259
rect	173	258	174	259
rect	176	258	177	259
rect	188	258	189	259
rect	194	258	195	259
rect	197	258	198	259
rect	220	258	221	259
rect	223	258	224	259
rect	232	258	233	259
rect	248	258	249	259
rect	251	258	252	259
rect	254	258	255	259
rect	257	258	258	259
rect	266	258	267	259
rect	269	258	270	259
rect	272	258	273	259
rect	280	258	281	259
rect	284	258	285	259
rect	287	258	288	259
rect	296	258	297	259
rect	305	258	306	259
rect	308	258	309	259
rect	314	258	315	259
rect	324	258	325	259
rect	333	258	334	259
rect	336	258	337	259
rect	339	258	340	259
rect	348	258	349	259
rect	357	258	358	259
rect	366	258	367	259
rect	373	258	374	259
rect	376	258	377	259
rect	379	258	380	259
rect	4	259	5	260
rect	21	259	22	260
rect	24	259	25	260
rect	27	259	28	260
rect	30	259	31	260
rect	39	259	40	260
rect	48	259	49	260
rect	51	259	52	260
rect	54	259	55	260
rect	60	259	61	260
rect	83	259	84	260
rect	89	259	90	260
rect	103	259	104	260
rect	106	259	107	260
rect	109	259	110	260
rect	112	259	113	260
rect	118	259	119	260
rect	134	259	135	260
rect	137	259	138	260
rect	140	259	141	260
rect	149	259	150	260
rect	161	259	162	260
rect	170	259	171	260
rect	176	259	177	260
rect	188	259	189	260
rect	194	259	195	260
rect	197	259	198	260
rect	220	259	221	260
rect	223	259	224	260
rect	232	259	233	260
rect	248	259	249	260
rect	251	259	252	260
rect	254	259	255	260
rect	269	259	270	260
rect	272	259	273	260
rect	280	259	281	260
rect	284	259	285	260
rect	287	259	288	260
rect	296	259	297	260
rect	305	259	306	260
rect	308	259	309	260
rect	314	259	315	260
rect	324	259	325	260
rect	333	259	334	260
rect	336	259	337	260
rect	339	259	340	260
rect	348	259	349	260
rect	357	259	358	260
rect	366	259	367	260
rect	373	259	374	260
rect	376	259	377	260
rect	4	260	5	261
rect	21	260	22	261
rect	24	260	25	261
rect	27	260	28	261
rect	30	260	31	261
rect	39	260	40	261
rect	48	260	49	261
rect	51	260	52	261
rect	54	260	55	261
rect	60	260	61	261
rect	63	260	64	261
rect	83	260	84	261
rect	89	260	90	261
rect	103	260	104	261
rect	106	260	107	261
rect	109	260	110	261
rect	112	260	113	261
rect	118	260	119	261
rect	134	260	135	261
rect	137	260	138	261
rect	140	260	141	261
rect	149	260	150	261
rect	161	260	162	261
rect	170	260	171	261
rect	176	260	177	261
rect	188	260	189	261
rect	194	260	195	261
rect	197	260	198	261
rect	200	260	201	261
rect	220	260	221	261
rect	223	260	224	261
rect	232	260	233	261
rect	248	260	249	261
rect	251	260	252	261
rect	254	260	255	261
rect	262	260	263	261
rect	269	260	270	261
rect	272	260	273	261
rect	280	260	281	261
rect	284	260	285	261
rect	287	260	288	261
rect	289	260	290	261
rect	296	260	297	261
rect	305	260	306	261
rect	308	260	309	261
rect	314	260	315	261
rect	324	260	325	261
rect	333	260	334	261
rect	336	260	337	261
rect	339	260	340	261
rect	348	260	349	261
rect	357	260	358	261
rect	366	260	367	261
rect	373	260	374	261
rect	376	260	377	261
rect	381	260	382	261
rect	4	261	5	262
rect	24	261	25	262
rect	27	261	28	262
rect	30	261	31	262
rect	39	261	40	262
rect	48	261	49	262
rect	51	261	52	262
rect	60	261	61	262
rect	63	261	64	262
rect	83	261	84	262
rect	89	261	90	262
rect	103	261	104	262
rect	106	261	107	262
rect	109	261	110	262
rect	112	261	113	262
rect	118	261	119	262
rect	134	261	135	262
rect	137	261	138	262
rect	149	261	150	262
rect	161	261	162	262
rect	170	261	171	262
rect	188	261	189	262
rect	194	261	195	262
rect	197	261	198	262
rect	200	261	201	262
rect	220	261	221	262
rect	223	261	224	262
rect	232	261	233	262
rect	248	261	249	262
rect	251	261	252	262
rect	262	261	263	262
rect	269	261	270	262
rect	280	261	281	262
rect	287	261	288	262
rect	289	261	290	262
rect	296	261	297	262
rect	305	261	306	262
rect	308	261	309	262
rect	314	261	315	262
rect	324	261	325	262
rect	336	261	337	262
rect	339	261	340	262
rect	348	261	349	262
rect	366	261	367	262
rect	373	261	374	262
rect	376	261	377	262
rect	381	261	382	262
rect	4	262	5	263
rect	24	262	25	263
rect	27	262	28	263
rect	30	262	31	263
rect	33	262	34	263
rect	39	262	40	263
rect	48	262	49	263
rect	51	262	52	263
rect	57	262	58	263
rect	60	262	61	263
rect	63	262	64	263
rect	83	262	84	263
rect	89	262	90	263
rect	103	262	104	263
rect	106	262	107	263
rect	109	262	110	263
rect	112	262	113	263
rect	118	262	119	263
rect	134	262	135	263
rect	137	262	138	263
rect	149	262	150	263
rect	151	262	152	263
rect	161	262	162	263
rect	163	262	164	263
rect	170	262	171	263
rect	172	262	173	263
rect	185	262	186	263
rect	188	262	189	263
rect	194	262	195	263
rect	197	262	198	263
rect	200	262	201	263
rect	220	262	221	263
rect	223	262	224	263
rect	232	262	233	263
rect	248	262	249	263
rect	251	262	252	263
rect	262	262	263	263
rect	265	262	266	263
rect	269	262	270	263
rect	277	262	278	263
rect	280	262	281	263
rect	287	262	288	263
rect	289	262	290	263
rect	296	262	297	263
rect	298	262	299	263
rect	305	262	306	263
rect	308	262	309	263
rect	314	262	315	263
rect	324	262	325	263
rect	336	262	337	263
rect	339	262	340	263
rect	341	262	342	263
rect	348	262	349	263
rect	366	262	367	263
rect	373	262	374	263
rect	376	262	377	263
rect	378	262	379	263
rect	381	262	382	263
rect	4	263	5	264
rect	30	263	31	264
rect	33	263	34	264
rect	39	263	40	264
rect	48	263	49	264
rect	57	263	58	264
rect	63	263	64	264
rect	83	263	84	264
rect	89	263	90	264
rect	103	263	104	264
rect	106	263	107	264
rect	109	263	110	264
rect	118	263	119	264
rect	137	263	138	264
rect	149	263	150	264
rect	151	263	152	264
rect	163	263	164	264
rect	170	263	171	264
rect	172	263	173	264
rect	185	263	186	264
rect	188	263	189	264
rect	197	263	198	264
rect	200	263	201	264
rect	220	263	221	264
rect	223	263	224	264
rect	232	263	233	264
rect	248	263	249	264
rect	251	263	252	264
rect	262	263	263	264
rect	265	263	266	264
rect	269	263	270	264
rect	277	263	278	264
rect	280	263	281	264
rect	287	263	288	264
rect	289	263	290	264
rect	296	263	297	264
rect	298	263	299	264
rect	305	263	306	264
rect	308	263	309	264
rect	314	263	315	264
rect	324	263	325	264
rect	341	263	342	264
rect	366	263	367	264
rect	373	263	374	264
rect	376	263	377	264
rect	378	263	379	264
rect	381	263	382	264
rect	4	264	5	265
rect	21	264	22	265
rect	30	264	31	265
rect	33	264	34	265
rect	36	264	37	265
rect	39	264	40	265
rect	48	264	49	265
rect	54	264	55	265
rect	57	264	58	265
rect	63	264	64	265
rect	66	264	67	265
rect	83	264	84	265
rect	89	264	90	265
rect	103	264	104	265
rect	106	264	107	265
rect	109	264	110	265
rect	118	264	119	265
rect	124	264	125	265
rect	137	264	138	265
rect	139	264	140	265
rect	149	264	150	265
rect	151	264	152	265
rect	163	264	164	265
rect	170	264	171	265
rect	172	264	173	265
rect	175	264	176	265
rect	185	264	186	265
rect	188	264	189	265
rect	197	264	198	265
rect	200	264	201	265
rect	220	264	221	265
rect	223	264	224	265
rect	232	264	233	265
rect	248	264	249	265
rect	251	264	252	265
rect	262	264	263	265
rect	265	264	266	265
rect	269	264	270	265
rect	277	264	278	265
rect	280	264	281	265
rect	287	264	288	265
rect	289	264	290	265
rect	296	264	297	265
rect	298	264	299	265
rect	305	264	306	265
rect	308	264	309	265
rect	314	264	315	265
rect	320	264	321	265
rect	324	264	325	265
rect	326	264	327	265
rect	341	264	342	265
rect	344	264	345	265
rect	360	264	361	265
rect	366	264	367	265
rect	373	264	374	265
rect	376	264	377	265
rect	378	264	379	265
rect	381	264	382	265
rect	4	265	5	266
rect	21	265	22	266
rect	33	265	34	266
rect	36	265	37	266
rect	54	265	55	266
rect	57	265	58	266
rect	63	265	64	266
rect	66	265	67	266
rect	83	265	84	266
rect	106	265	107	266
rect	109	265	110	266
rect	118	265	119	266
rect	124	265	125	266
rect	137	265	138	266
rect	139	265	140	266
rect	149	265	150	266
rect	151	265	152	266
rect	163	265	164	266
rect	172	265	173	266
rect	175	265	176	266
rect	185	265	186	266
rect	188	265	189	266
rect	200	265	201	266
rect	220	265	221	266
rect	232	265	233	266
rect	248	265	249	266
rect	262	265	263	266
rect	265	265	266	266
rect	269	265	270	266
rect	277	265	278	266
rect	280	265	281	266
rect	289	265	290	266
rect	296	265	297	266
rect	298	265	299	266
rect	305	265	306	266
rect	308	265	309	266
rect	320	265	321	266
rect	324	265	325	266
rect	326	265	327	266
rect	341	265	342	266
rect	344	265	345	266
rect	360	265	361	266
rect	366	265	367	266
rect	376	265	377	266
rect	378	265	379	266
rect	381	265	382	266
rect	4	266	5	267
rect	21	266	22	267
rect	24	266	25	267
rect	33	266	34	267
rect	36	266	37	267
rect	45	266	46	267
rect	54	266	55	267
rect	57	266	58	267
rect	63	266	64	267
rect	66	266	67	267
rect	75	266	76	267
rect	83	266	84	267
rect	91	266	92	267
rect	106	266	107	267
rect	109	266	110	267
rect	112	266	113	267
rect	118	266	119	267
rect	124	266	125	267
rect	133	266	134	267
rect	137	266	138	267
rect	139	266	140	267
rect	142	266	143	267
rect	149	266	150	267
rect	151	266	152	267
rect	160	266	161	267
rect	163	266	164	267
rect	172	266	173	267
rect	175	266	176	267
rect	185	266	186	267
rect	188	266	189	267
rect	191	266	192	267
rect	200	266	201	267
rect	220	266	221	267
rect	227	266	228	267
rect	232	266	233	267
rect	248	266	249	267
rect	262	266	263	267
rect	265	266	266	267
rect	269	266	270	267
rect	274	266	275	267
rect	277	266	278	267
rect	280	266	281	267
rect	283	266	284	267
rect	289	266	290	267
rect	296	266	297	267
rect	298	266	299	267
rect	305	266	306	267
rect	308	266	309	267
rect	320	266	321	267
rect	324	266	325	267
rect	326	266	327	267
rect	341	266	342	267
rect	344	266	345	267
rect	360	266	361	267
rect	363	266	364	267
rect	366	266	367	267
rect	376	266	377	267
rect	378	266	379	267
rect	381	266	382	267
rect	387	266	388	267
rect	21	267	22	268
rect	24	267	25	268
rect	33	267	34	268
rect	36	267	37	268
rect	45	267	46	268
rect	54	267	55	268
rect	57	267	58	268
rect	63	267	64	268
rect	66	267	67	268
rect	75	267	76	268
rect	91	267	92	268
rect	112	267	113	268
rect	124	267	125	268
rect	133	267	134	268
rect	139	267	140	268
rect	142	267	143	268
rect	151	267	152	268
rect	160	267	161	268
rect	163	267	164	268
rect	172	267	173	268
rect	175	267	176	268
rect	185	267	186	268
rect	191	267	192	268
rect	200	267	201	268
rect	227	267	228	268
rect	262	267	263	268
rect	265	267	266	268
rect	274	267	275	268
rect	277	267	278	268
rect	280	267	281	268
rect	283	267	284	268
rect	289	267	290	268
rect	298	267	299	268
rect	308	267	309	268
rect	320	267	321	268
rect	326	267	327	268
rect	341	267	342	268
rect	344	267	345	268
rect	360	267	361	268
rect	363	267	364	268
rect	366	267	367	268
rect	378	267	379	268
rect	381	267	382	268
rect	387	267	388	268
rect	21	268	22	269
rect	24	268	25	269
rect	33	268	34	269
rect	36	268	37	269
rect	45	268	46	269
rect	54	268	55	269
rect	57	268	58	269
rect	60	268	61	269
rect	63	268	64	269
rect	66	268	67	269
rect	75	268	76	269
rect	91	268	92	269
rect	100	268	101	269
rect	103	268	104	269
rect	112	268	113	269
rect	115	268	116	269
rect	124	268	125	269
rect	127	268	128	269
rect	130	268	131	269
rect	133	268	134	269
rect	139	268	140	269
rect	142	268	143	269
rect	151	268	152	269
rect	160	268	161	269
rect	163	268	164	269
rect	169	268	170	269
rect	172	268	173	269
rect	175	268	176	269
rect	185	268	186	269
rect	191	268	192	269
rect	194	268	195	269
rect	200	268	201	269
rect	224	268	225	269
rect	227	268	228	269
rect	236	268	237	269
rect	259	268	260	269
rect	262	268	263	269
rect	265	268	266	269
rect	274	268	275	269
rect	277	268	278	269
rect	280	268	281	269
rect	283	268	284	269
rect	289	268	290	269
rect	292	268	293	269
rect	298	268	299	269
rect	302	268	303	269
rect	308	268	309	269
rect	317	268	318	269
rect	320	268	321	269
rect	323	268	324	269
rect	326	268	327	269
rect	329	268	330	269
rect	335	268	336	269
rect	338	268	339	269
rect	341	268	342	269
rect	344	268	345	269
rect	357	268	358	269
rect	360	268	361	269
rect	363	268	364	269
rect	366	268	367	269
rect	369	268	370	269
rect	378	268	379	269
rect	381	268	382	269
rect	387	268	388	269
rect	1	275	2	276
rect	11	275	12	276
rect	21	275	22	276
rect	24	275	25	276
rect	33	275	34	276
rect	36	275	37	276
rect	45	275	46	276
rect	54	275	55	276
rect	57	275	58	276
rect	60	275	61	276
rect	63	275	64	276
rect	66	275	67	276
rect	75	275	76	276
rect	91	275	92	276
rect	100	275	101	276
rect	103	275	104	276
rect	112	275	113	276
rect	115	275	116	276
rect	118	275	119	276
rect	124	275	125	276
rect	127	275	128	276
rect	130	275	131	276
rect	139	275	140	276
rect	142	275	143	276
rect	145	275	146	276
rect	151	275	152	276
rect	154	275	155	276
rect	160	275	161	276
rect	169	275	170	276
rect	172	275	173	276
rect	175	275	176	276
rect	178	275	179	276
rect	185	275	186	276
rect	191	275	192	276
rect	194	275	195	276
rect	197	275	198	276
rect	224	275	225	276
rect	227	275	228	276
rect	236	275	237	276
rect	259	275	260	276
rect	262	275	263	276
rect	265	275	266	276
rect	274	275	275	276
rect	277	275	278	276
rect	280	275	281	276
rect	283	275	284	276
rect	292	275	293	276
rect	308	275	309	276
rect	317	275	318	276
rect	320	275	321	276
rect	323	275	324	276
rect	326	275	327	276
rect	335	275	336	276
rect	338	275	339	276
rect	341	275	342	276
rect	344	275	345	276
rect	350	275	351	276
rect	360	275	361	276
rect	363	275	364	276
rect	366	275	367	276
rect	369	275	370	276
rect	372	275	373	276
rect	378	275	379	276
rect	381	275	382	276
rect	1	276	2	277
rect	11	276	12	277
rect	21	276	22	277
rect	24	276	25	277
rect	33	276	34	277
rect	36	276	37	277
rect	45	276	46	277
rect	54	276	55	277
rect	57	276	58	277
rect	60	276	61	277
rect	63	276	64	277
rect	66	276	67	277
rect	75	276	76	277
rect	91	276	92	277
rect	100	276	101	277
rect	103	276	104	277
rect	112	276	113	277
rect	115	276	116	277
rect	118	276	119	277
rect	124	276	125	277
rect	127	276	128	277
rect	130	276	131	277
rect	139	276	140	277
rect	142	276	143	277
rect	145	276	146	277
rect	151	276	152	277
rect	154	276	155	277
rect	160	276	161	277
rect	169	276	170	277
rect	172	276	173	277
rect	175	276	176	277
rect	178	276	179	277
rect	185	276	186	277
rect	191	276	192	277
rect	194	276	195	277
rect	197	276	198	277
rect	224	276	225	277
rect	227	276	228	277
rect	236	276	237	277
rect	259	276	260	277
rect	262	276	263	277
rect	265	276	266	277
rect	274	276	275	277
rect	277	276	278	277
rect	280	276	281	277
rect	283	276	284	277
rect	308	276	309	277
rect	317	276	318	277
rect	320	276	321	277
rect	323	276	324	277
rect	326	276	327	277
rect	335	276	336	277
rect	338	276	339	277
rect	341	276	342	277
rect	344	276	345	277
rect	350	276	351	277
rect	360	276	361	277
rect	363	276	364	277
rect	366	276	367	277
rect	369	276	370	277
rect	372	276	373	277
rect	378	276	379	277
rect	1	277	2	278
rect	11	277	12	278
rect	21	277	22	278
rect	24	277	25	278
rect	33	277	34	278
rect	36	277	37	278
rect	45	277	46	278
rect	54	277	55	278
rect	57	277	58	278
rect	60	277	61	278
rect	63	277	64	278
rect	66	277	67	278
rect	75	277	76	278
rect	91	277	92	278
rect	100	277	101	278
rect	103	277	104	278
rect	112	277	113	278
rect	115	277	116	278
rect	118	277	119	278
rect	124	277	125	278
rect	127	277	128	278
rect	130	277	131	278
rect	139	277	140	278
rect	142	277	143	278
rect	145	277	146	278
rect	151	277	152	278
rect	154	277	155	278
rect	160	277	161	278
rect	169	277	170	278
rect	172	277	173	278
rect	175	277	176	278
rect	178	277	179	278
rect	185	277	186	278
rect	191	277	192	278
rect	194	277	195	278
rect	197	277	198	278
rect	224	277	225	278
rect	227	277	228	278
rect	236	277	237	278
rect	259	277	260	278
rect	262	277	263	278
rect	265	277	266	278
rect	274	277	275	278
rect	277	277	278	278
rect	280	277	281	278
rect	283	277	284	278
rect	308	277	309	278
rect	311	277	312	278
rect	317	277	318	278
rect	320	277	321	278
rect	323	277	324	278
rect	326	277	327	278
rect	335	277	336	278
rect	338	277	339	278
rect	341	277	342	278
rect	344	277	345	278
rect	350	277	351	278
rect	360	277	361	278
rect	363	277	364	278
rect	366	277	367	278
rect	369	277	370	278
rect	372	277	373	278
rect	378	277	379	278
rect	387	277	388	278
rect	1	278	2	279
rect	11	278	12	279
rect	21	278	22	279
rect	24	278	25	279
rect	33	278	34	279
rect	36	278	37	279
rect	45	278	46	279
rect	54	278	55	279
rect	57	278	58	279
rect	60	278	61	279
rect	63	278	64	279
rect	66	278	67	279
rect	75	278	76	279
rect	91	278	92	279
rect	100	278	101	279
rect	103	278	104	279
rect	112	278	113	279
rect	115	278	116	279
rect	118	278	119	279
rect	124	278	125	279
rect	127	278	128	279
rect	130	278	131	279
rect	139	278	140	279
rect	142	278	143	279
rect	145	278	146	279
rect	151	278	152	279
rect	154	278	155	279
rect	160	278	161	279
rect	169	278	170	279
rect	172	278	173	279
rect	175	278	176	279
rect	178	278	179	279
rect	185	278	186	279
rect	191	278	192	279
rect	194	278	195	279
rect	197	278	198	279
rect	224	278	225	279
rect	227	278	228	279
rect	236	278	237	279
rect	259	278	260	279
rect	262	278	263	279
rect	265	278	266	279
rect	274	278	275	279
rect	277	278	278	279
rect	280	278	281	279
rect	283	278	284	279
rect	311	278	312	279
rect	317	278	318	279
rect	320	278	321	279
rect	323	278	324	279
rect	326	278	327	279
rect	335	278	336	279
rect	341	278	342	279
rect	344	278	345	279
rect	350	278	351	279
rect	363	278	364	279
rect	366	278	367	279
rect	369	278	370	279
rect	372	278	373	279
rect	378	278	379	279
rect	387	278	388	279
rect	1	279	2	280
rect	11	279	12	280
rect	21	279	22	280
rect	24	279	25	280
rect	33	279	34	280
rect	36	279	37	280
rect	45	279	46	280
rect	54	279	55	280
rect	57	279	58	280
rect	60	279	61	280
rect	63	279	64	280
rect	66	279	67	280
rect	75	279	76	280
rect	91	279	92	280
rect	100	279	101	280
rect	103	279	104	280
rect	112	279	113	280
rect	115	279	116	280
rect	118	279	119	280
rect	124	279	125	280
rect	127	279	128	280
rect	130	279	131	280
rect	139	279	140	280
rect	142	279	143	280
rect	145	279	146	280
rect	151	279	152	280
rect	154	279	155	280
rect	160	279	161	280
rect	169	279	170	280
rect	172	279	173	280
rect	175	279	176	280
rect	178	279	179	280
rect	185	279	186	280
rect	191	279	192	280
rect	194	279	195	280
rect	197	279	198	280
rect	224	279	225	280
rect	227	279	228	280
rect	236	279	237	280
rect	259	279	260	280
rect	262	279	263	280
rect	265	279	266	280
rect	274	279	275	280
rect	277	279	278	280
rect	280	279	281	280
rect	283	279	284	280
rect	289	279	290	280
rect	311	279	312	280
rect	317	279	318	280
rect	320	279	321	280
rect	323	279	324	280
rect	326	279	327	280
rect	335	279	336	280
rect	341	279	342	280
rect	344	279	345	280
rect	350	279	351	280
rect	357	279	358	280
rect	363	279	364	280
rect	366	279	367	280
rect	369	279	370	280
rect	372	279	373	280
rect	378	279	379	280
rect	381	279	382	280
rect	387	279	388	280
rect	1	280	2	281
rect	11	280	12	281
rect	21	280	22	281
rect	24	280	25	281
rect	33	280	34	281
rect	36	280	37	281
rect	45	280	46	281
rect	54	280	55	281
rect	57	280	58	281
rect	60	280	61	281
rect	63	280	64	281
rect	66	280	67	281
rect	75	280	76	281
rect	91	280	92	281
rect	100	280	101	281
rect	103	280	104	281
rect	112	280	113	281
rect	115	280	116	281
rect	118	280	119	281
rect	124	280	125	281
rect	127	280	128	281
rect	130	280	131	281
rect	139	280	140	281
rect	142	280	143	281
rect	145	280	146	281
rect	151	280	152	281
rect	154	280	155	281
rect	160	280	161	281
rect	169	280	170	281
rect	172	280	173	281
rect	175	280	176	281
rect	185	280	186	281
rect	194	280	195	281
rect	197	280	198	281
rect	224	280	225	281
rect	227	280	228	281
rect	236	280	237	281
rect	259	280	260	281
rect	262	280	263	281
rect	265	280	266	281
rect	277	280	278	281
rect	280	280	281	281
rect	283	280	284	281
rect	289	280	290	281
rect	311	280	312	281
rect	317	280	318	281
rect	320	280	321	281
rect	323	280	324	281
rect	326	280	327	281
rect	341	280	342	281
rect	344	280	345	281
rect	350	280	351	281
rect	357	280	358	281
rect	363	280	364	281
rect	366	280	367	281
rect	369	280	370	281
rect	372	280	373	281
rect	378	280	379	281
rect	381	280	382	281
rect	387	280	388	281
rect	1	281	2	282
rect	11	281	12	282
rect	21	281	22	282
rect	24	281	25	282
rect	33	281	34	282
rect	36	281	37	282
rect	45	281	46	282
rect	54	281	55	282
rect	57	281	58	282
rect	60	281	61	282
rect	63	281	64	282
rect	66	281	67	282
rect	75	281	76	282
rect	91	281	92	282
rect	100	281	101	282
rect	103	281	104	282
rect	112	281	113	282
rect	115	281	116	282
rect	118	281	119	282
rect	124	281	125	282
rect	127	281	128	282
rect	130	281	131	282
rect	139	281	140	282
rect	142	281	143	282
rect	145	281	146	282
rect	151	281	152	282
rect	154	281	155	282
rect	160	281	161	282
rect	169	281	170	282
rect	172	281	173	282
rect	175	281	176	282
rect	179	281	180	282
rect	185	281	186	282
rect	188	281	189	282
rect	194	281	195	282
rect	197	281	198	282
rect	224	281	225	282
rect	227	281	228	282
rect	236	281	237	282
rect	259	281	260	282
rect	262	281	263	282
rect	265	281	266	282
rect	277	281	278	282
rect	280	281	281	282
rect	283	281	284	282
rect	289	281	290	282
rect	308	281	309	282
rect	311	281	312	282
rect	317	281	318	282
rect	320	281	321	282
rect	323	281	324	282
rect	326	281	327	282
rect	341	281	342	282
rect	344	281	345	282
rect	350	281	351	282
rect	357	281	358	282
rect	360	281	361	282
rect	363	281	364	282
rect	366	281	367	282
rect	369	281	370	282
rect	372	281	373	282
rect	378	281	379	282
rect	381	281	382	282
rect	387	281	388	282
rect	1	282	2	283
rect	11	282	12	283
rect	21	282	22	283
rect	24	282	25	283
rect	33	282	34	283
rect	36	282	37	283
rect	45	282	46	283
rect	54	282	55	283
rect	57	282	58	283
rect	60	282	61	283
rect	66	282	67	283
rect	75	282	76	283
rect	91	282	92	283
rect	100	282	101	283
rect	103	282	104	283
rect	112	282	113	283
rect	118	282	119	283
rect	124	282	125	283
rect	127	282	128	283
rect	139	282	140	283
rect	142	282	143	283
rect	151	282	152	283
rect	154	282	155	283
rect	160	282	161	283
rect	169	282	170	283
rect	175	282	176	283
rect	179	282	180	283
rect	188	282	189	283
rect	194	282	195	283
rect	197	282	198	283
rect	224	282	225	283
rect	227	282	228	283
rect	236	282	237	283
rect	259	282	260	283
rect	262	282	263	283
rect	265	282	266	283
rect	283	282	284	283
rect	289	282	290	283
rect	308	282	309	283
rect	311	282	312	283
rect	317	282	318	283
rect	320	282	321	283
rect	323	282	324	283
rect	341	282	342	283
rect	350	282	351	283
rect	357	282	358	283
rect	360	282	361	283
rect	363	282	364	283
rect	366	282	367	283
rect	369	282	370	283
rect	378	282	379	283
rect	381	282	382	283
rect	387	282	388	283
rect	1	283	2	284
rect	11	283	12	284
rect	21	283	22	284
rect	24	283	25	284
rect	33	283	34	284
rect	36	283	37	284
rect	45	283	46	284
rect	54	283	55	284
rect	57	283	58	284
rect	60	283	61	284
rect	66	283	67	284
rect	69	283	70	284
rect	75	283	76	284
rect	91	283	92	284
rect	100	283	101	284
rect	103	283	104	284
rect	107	283	108	284
rect	112	283	113	284
rect	118	283	119	284
rect	124	283	125	284
rect	127	283	128	284
rect	133	283	134	284
rect	139	283	140	284
rect	142	283	143	284
rect	151	283	152	284
rect	154	283	155	284
rect	160	283	161	284
rect	167	283	168	284
rect	169	283	170	284
rect	175	283	176	284
rect	179	283	180	284
rect	182	283	183	284
rect	188	283	189	284
rect	194	283	195	284
rect	197	283	198	284
rect	200	283	201	284
rect	224	283	225	284
rect	227	283	228	284
rect	236	283	237	284
rect	259	283	260	284
rect	262	283	263	284
rect	265	283	266	284
rect	274	283	275	284
rect	283	283	284	284
rect	289	283	290	284
rect	292	283	293	284
rect	308	283	309	284
rect	311	283	312	284
rect	317	283	318	284
rect	320	283	321	284
rect	323	283	324	284
rect	330	283	331	284
rect	336	283	337	284
rect	341	283	342	284
rect	350	283	351	284
rect	357	283	358	284
rect	360	283	361	284
rect	363	283	364	284
rect	366	283	367	284
rect	369	283	370	284
rect	378	283	379	284
rect	381	283	382	284
rect	387	283	388	284
rect	393	283	394	284
rect	1	284	2	285
rect	11	284	12	285
rect	21	284	22	285
rect	24	284	25	285
rect	33	284	34	285
rect	36	284	37	285
rect	45	284	46	285
rect	54	284	55	285
rect	57	284	58	285
rect	69	284	70	285
rect	75	284	76	285
rect	91	284	92	285
rect	100	284	101	285
rect	103	284	104	285
rect	107	284	108	285
rect	118	284	119	285
rect	124	284	125	285
rect	133	284	134	285
rect	139	284	140	285
rect	151	284	152	285
rect	154	284	155	285
rect	167	284	168	285
rect	175	284	176	285
rect	179	284	180	285
rect	182	284	183	285
rect	188	284	189	285
rect	194	284	195	285
rect	197	284	198	285
rect	200	284	201	285
rect	224	284	225	285
rect	262	284	263	285
rect	265	284	266	285
rect	274	284	275	285
rect	289	284	290	285
rect	292	284	293	285
rect	308	284	309	285
rect	311	284	312	285
rect	317	284	318	285
rect	323	284	324	285
rect	330	284	331	285
rect	336	284	337	285
rect	341	284	342	285
rect	350	284	351	285
rect	357	284	358	285
rect	360	284	361	285
rect	363	284	364	285
rect	369	284	370	285
rect	378	284	379	285
rect	381	284	382	285
rect	387	284	388	285
rect	393	284	394	285
rect	1	285	2	286
rect	11	285	12	286
rect	21	285	22	286
rect	24	285	25	286
rect	33	285	34	286
rect	36	285	37	286
rect	45	285	46	286
rect	54	285	55	286
rect	57	285	58	286
rect	63	285	64	286
rect	69	285	70	286
rect	72	285	73	286
rect	75	285	76	286
rect	91	285	92	286
rect	100	285	101	286
rect	103	285	104	286
rect	107	285	108	286
rect	109	285	110	286
rect	118	285	119	286
rect	124	285	125	286
rect	130	285	131	286
rect	133	285	134	286
rect	139	285	140	286
rect	148	285	149	286
rect	151	285	152	286
rect	154	285	155	286
rect	164	285	165	286
rect	167	285	168	286
rect	175	285	176	286
rect	179	285	180	286
rect	182	285	183	286
rect	188	285	189	286
rect	194	285	195	286
rect	197	285	198	286
rect	200	285	201	286
rect	203	285	204	286
rect	206	285	207	286
rect	215	285	216	286
rect	224	285	225	286
rect	230	285	231	286
rect	246	285	247	286
rect	262	285	263	286
rect	265	285	266	286
rect	271	285	272	286
rect	274	285	275	286
rect	277	285	278	286
rect	289	285	290	286
rect	292	285	293	286
rect	308	285	309	286
rect	311	285	312	286
rect	317	285	318	286
rect	323	285	324	286
rect	330	285	331	286
rect	336	285	337	286
rect	341	285	342	286
rect	345	285	346	286
rect	350	285	351	286
rect	357	285	358	286
rect	360	285	361	286
rect	363	285	364	286
rect	369	285	370	286
rect	375	285	376	286
rect	378	285	379	286
rect	381	285	382	286
rect	387	285	388	286
rect	393	285	394	286
rect	1	286	2	287
rect	11	286	12	287
rect	21	286	22	287
rect	33	286	34	287
rect	45	286	46	287
rect	54	286	55	287
rect	63	286	64	287
rect	69	286	70	287
rect	72	286	73	287
rect	75	286	76	287
rect	91	286	92	287
rect	103	286	104	287
rect	107	286	108	287
rect	109	286	110	287
rect	130	286	131	287
rect	133	286	134	287
rect	139	286	140	287
rect	148	286	149	287
rect	154	286	155	287
rect	164	286	165	287
rect	167	286	168	287
rect	179	286	180	287
rect	182	286	183	287
rect	188	286	189	287
rect	194	286	195	287
rect	200	286	201	287
rect	203	286	204	287
rect	206	286	207	287
rect	215	286	216	287
rect	224	286	225	287
rect	230	286	231	287
rect	246	286	247	287
rect	271	286	272	287
rect	274	286	275	287
rect	277	286	278	287
rect	289	286	290	287
rect	292	286	293	287
rect	308	286	309	287
rect	311	286	312	287
rect	330	286	331	287
rect	336	286	337	287
rect	345	286	346	287
rect	357	286	358	287
rect	360	286	361	287
rect	369	286	370	287
rect	375	286	376	287
rect	378	286	379	287
rect	381	286	382	287
rect	387	286	388	287
rect	393	286	394	287
rect	1	287	2	288
rect	11	287	12	288
rect	21	287	22	288
rect	23	287	24	288
rect	33	287	34	288
rect	42	287	43	288
rect	45	287	46	288
rect	54	287	55	288
rect	63	287	64	288
rect	66	287	67	288
rect	69	287	70	288
rect	72	287	73	288
rect	75	287	76	288
rect	91	287	92	288
rect	103	287	104	288
rect	107	287	108	288
rect	109	287	110	288
rect	112	287	113	288
rect	115	287	116	288
rect	130	287	131	288
rect	133	287	134	288
rect	139	287	140	288
rect	145	287	146	288
rect	148	287	149	288
rect	154	287	155	288
rect	164	287	165	288
rect	167	287	168	288
rect	170	287	171	288
rect	179	287	180	288
rect	182	287	183	288
rect	188	287	189	288
rect	191	287	192	288
rect	194	287	195	288
rect	200	287	201	288
rect	203	287	204	288
rect	206	287	207	288
rect	215	287	216	288
rect	218	287	219	288
rect	224	287	225	288
rect	227	287	228	288
rect	230	287	231	288
rect	236	287	237	288
rect	246	287	247	288
rect	255	287	256	288
rect	271	287	272	288
rect	274	287	275	288
rect	277	287	278	288
rect	280	287	281	288
rect	289	287	290	288
rect	292	287	293	288
rect	308	287	309	288
rect	311	287	312	288
rect	318	287	319	288
rect	324	287	325	288
rect	330	287	331	288
rect	333	287	334	288
rect	336	287	337	288
rect	345	287	346	288
rect	354	287	355	288
rect	357	287	358	288
rect	360	287	361	288
rect	369	287	370	288
rect	372	287	373	288
rect	375	287	376	288
rect	378	287	379	288
rect	381	287	382	288
rect	387	287	388	288
rect	393	287	394	288
rect	23	288	24	289
rect	42	288	43	289
rect	63	288	64	289
rect	66	288	67	289
rect	69	288	70	289
rect	72	288	73	289
rect	109	288	110	289
rect	112	288	113	289
rect	115	288	116	289
rect	130	288	131	289
rect	133	288	134	289
rect	139	288	140	289
rect	145	288	146	289
rect	148	288	149	289
rect	164	288	165	289
rect	167	288	168	289
rect	170	288	171	289
rect	179	288	180	289
rect	182	288	183	289
rect	188	288	189	289
rect	191	288	192	289
rect	200	288	201	289
rect	203	288	204	289
rect	206	288	207	289
rect	215	288	216	289
rect	218	288	219	289
rect	227	288	228	289
rect	230	288	231	289
rect	236	288	237	289
rect	246	288	247	289
rect	255	288	256	289
rect	271	288	272	289
rect	274	288	275	289
rect	277	288	278	289
rect	280	288	281	289
rect	289	288	290	289
rect	292	288	293	289
rect	308	288	309	289
rect	311	288	312	289
rect	318	288	319	289
rect	324	288	325	289
rect	330	288	331	289
rect	333	288	334	289
rect	336	288	337	289
rect	345	288	346	289
rect	354	288	355	289
rect	357	288	358	289
rect	360	288	361	289
rect	372	288	373	289
rect	375	288	376	289
rect	378	288	379	289
rect	381	288	382	289
rect	387	288	388	289
rect	393	288	394	289
rect	14	289	15	290
rect	23	289	24	290
rect	39	289	40	290
rect	42	289	43	290
rect	51	289	52	290
rect	60	289	61	290
rect	63	289	64	290
rect	66	289	67	290
rect	69	289	70	290
rect	72	289	73	290
rect	81	289	82	290
rect	97	289	98	290
rect	100	289	101	290
rect	109	289	110	290
rect	112	289	113	290
rect	115	289	116	290
rect	118	289	119	290
rect	121	289	122	290
rect	127	289	128	290
rect	130	289	131	290
rect	133	289	134	290
rect	139	289	140	290
rect	142	289	143	290
rect	145	289	146	290
rect	148	289	149	290
rect	151	289	152	290
rect	164	289	165	290
rect	167	289	168	290
rect	170	289	171	290
rect	179	289	180	290
rect	182	289	183	290
rect	185	289	186	290
rect	188	289	189	290
rect	191	289	192	290
rect	200	289	201	290
rect	203	289	204	290
rect	206	289	207	290
rect	209	289	210	290
rect	215	289	216	290
rect	218	289	219	290
rect	227	289	228	290
rect	230	289	231	290
rect	236	289	237	290
rect	246	289	247	290
rect	255	289	256	290
rect	271	289	272	290
rect	274	289	275	290
rect	277	289	278	290
rect	280	289	281	290
rect	289	289	290	290
rect	292	289	293	290
rect	308	289	309	290
rect	311	289	312	290
rect	318	289	319	290
rect	324	289	325	290
rect	330	289	331	290
rect	333	289	334	290
rect	336	289	337	290
rect	345	289	346	290
rect	351	289	352	290
rect	354	289	355	290
rect	357	289	358	290
rect	360	289	361	290
rect	363	289	364	290
rect	372	289	373	290
rect	375	289	376	290
rect	378	289	379	290
rect	381	289	382	290
rect	387	289	388	290
rect	393	289	394	290
rect	4	296	5	297
rect	8	296	9	297
rect	14	296	15	297
rect	23	296	24	297
rect	39	296	40	297
rect	42	296	43	297
rect	51	296	52	297
rect	60	296	61	297
rect	63	296	64	297
rect	66	296	67	297
rect	69	296	70	297
rect	72	296	73	297
rect	81	296	82	297
rect	97	296	98	297
rect	100	296	101	297
rect	109	296	110	297
rect	112	296	113	297
rect	115	296	116	297
rect	118	296	119	297
rect	121	296	122	297
rect	124	296	125	297
rect	127	296	128	297
rect	130	296	131	297
rect	133	296	134	297
rect	139	296	140	297
rect	142	296	143	297
rect	145	296	146	297
rect	148	296	149	297
rect	158	296	159	297
rect	164	296	165	297
rect	167	296	168	297
rect	170	296	171	297
rect	176	296	177	297
rect	179	296	180	297
rect	182	296	183	297
rect	185	296	186	297
rect	188	296	189	297
rect	191	296	192	297
rect	197	296	198	297
rect	200	296	201	297
rect	203	296	204	297
rect	206	296	207	297
rect	209	296	210	297
rect	218	296	219	297
rect	224	296	225	297
rect	227	296	228	297
rect	230	296	231	297
rect	233	296	234	297
rect	246	296	247	297
rect	255	296	256	297
rect	271	296	272	297
rect	274	296	275	297
rect	277	296	278	297
rect	280	296	281	297
rect	289	296	290	297
rect	292	296	293	297
rect	308	296	309	297
rect	311	296	312	297
rect	324	296	325	297
rect	333	296	334	297
rect	336	296	337	297
rect	345	296	346	297
rect	348	296	349	297
rect	354	296	355	297
rect	357	296	358	297
rect	360	296	361	297
rect	363	296	364	297
rect	366	296	367	297
rect	372	296	373	297
rect	375	296	376	297
rect	378	296	379	297
rect	384	296	385	297
rect	387	296	388	297
rect	390	296	391	297
rect	400	296	401	297
rect	4	297	5	298
rect	8	297	9	298
rect	14	297	15	298
rect	23	297	24	298
rect	39	297	40	298
rect	42	297	43	298
rect	51	297	52	298
rect	60	297	61	298
rect	63	297	64	298
rect	66	297	67	298
rect	69	297	70	298
rect	72	297	73	298
rect	81	297	82	298
rect	97	297	98	298
rect	100	297	101	298
rect	109	297	110	298
rect	112	297	113	298
rect	115	297	116	298
rect	118	297	119	298
rect	121	297	122	298
rect	124	297	125	298
rect	127	297	128	298
rect	130	297	131	298
rect	139	297	140	298
rect	142	297	143	298
rect	145	297	146	298
rect	148	297	149	298
rect	158	297	159	298
rect	164	297	165	298
rect	167	297	168	298
rect	170	297	171	298
rect	176	297	177	298
rect	179	297	180	298
rect	182	297	183	298
rect	185	297	186	298
rect	188	297	189	298
rect	191	297	192	298
rect	197	297	198	298
rect	200	297	201	298
rect	206	297	207	298
rect	209	297	210	298
rect	218	297	219	298
rect	224	297	225	298
rect	227	297	228	298
rect	230	297	231	298
rect	233	297	234	298
rect	255	297	256	298
rect	271	297	272	298
rect	274	297	275	298
rect	277	297	278	298
rect	280	297	281	298
rect	289	297	290	298
rect	292	297	293	298
rect	308	297	309	298
rect	311	297	312	298
rect	324	297	325	298
rect	333	297	334	298
rect	336	297	337	298
rect	345	297	346	298
rect	348	297	349	298
rect	354	297	355	298
rect	357	297	358	298
rect	360	297	361	298
rect	363	297	364	298
rect	366	297	367	298
rect	372	297	373	298
rect	375	297	376	298
rect	378	297	379	298
rect	384	297	385	298
rect	387	297	388	298
rect	390	297	391	298
rect	400	297	401	298
rect	4	298	5	299
rect	8	298	9	299
rect	14	298	15	299
rect	23	298	24	299
rect	39	298	40	299
rect	42	298	43	299
rect	51	298	52	299
rect	60	298	61	299
rect	63	298	64	299
rect	66	298	67	299
rect	69	298	70	299
rect	72	298	73	299
rect	81	298	82	299
rect	97	298	98	299
rect	100	298	101	299
rect	109	298	110	299
rect	112	298	113	299
rect	115	298	116	299
rect	118	298	119	299
rect	121	298	122	299
rect	124	298	125	299
rect	127	298	128	299
rect	130	298	131	299
rect	137	298	138	299
rect	139	298	140	299
rect	142	298	143	299
rect	145	298	146	299
rect	148	298	149	299
rect	158	298	159	299
rect	164	298	165	299
rect	167	298	168	299
rect	170	298	171	299
rect	176	298	177	299
rect	179	298	180	299
rect	182	298	183	299
rect	185	298	186	299
rect	188	298	189	299
rect	191	298	192	299
rect	197	298	198	299
rect	200	298	201	299
rect	206	298	207	299
rect	209	298	210	299
rect	218	298	219	299
rect	224	298	225	299
rect	227	298	228	299
rect	230	298	231	299
rect	233	298	234	299
rect	242	298	243	299
rect	251	298	252	299
rect	255	298	256	299
rect	271	298	272	299
rect	274	298	275	299
rect	277	298	278	299
rect	280	298	281	299
rect	289	298	290	299
rect	292	298	293	299
rect	308	298	309	299
rect	311	298	312	299
rect	324	298	325	299
rect	333	298	334	299
rect	336	298	337	299
rect	345	298	346	299
rect	348	298	349	299
rect	354	298	355	299
rect	357	298	358	299
rect	360	298	361	299
rect	363	298	364	299
rect	366	298	367	299
rect	372	298	373	299
rect	375	298	376	299
rect	378	298	379	299
rect	384	298	385	299
rect	387	298	388	299
rect	390	298	391	299
rect	400	298	401	299
rect	4	299	5	300
rect	8	299	9	300
rect	14	299	15	300
rect	23	299	24	300
rect	39	299	40	300
rect	42	299	43	300
rect	51	299	52	300
rect	60	299	61	300
rect	63	299	64	300
rect	66	299	67	300
rect	69	299	70	300
rect	72	299	73	300
rect	81	299	82	300
rect	97	299	98	300
rect	100	299	101	300
rect	109	299	110	300
rect	112	299	113	300
rect	115	299	116	300
rect	118	299	119	300
rect	121	299	122	300
rect	124	299	125	300
rect	127	299	128	300
rect	137	299	138	300
rect	139	299	140	300
rect	142	299	143	300
rect	145	299	146	300
rect	148	299	149	300
rect	158	299	159	300
rect	164	299	165	300
rect	167	299	168	300
rect	170	299	171	300
rect	176	299	177	300
rect	179	299	180	300
rect	182	299	183	300
rect	188	299	189	300
rect	191	299	192	300
rect	197	299	198	300
rect	200	299	201	300
rect	206	299	207	300
rect	209	299	210	300
rect	224	299	225	300
rect	227	299	228	300
rect	230	299	231	300
rect	233	299	234	300
rect	242	299	243	300
rect	251	299	252	300
rect	255	299	256	300
rect	271	299	272	300
rect	274	299	275	300
rect	277	299	278	300
rect	280	299	281	300
rect	289	299	290	300
rect	292	299	293	300
rect	308	299	309	300
rect	311	299	312	300
rect	324	299	325	300
rect	333	299	334	300
rect	336	299	337	300
rect	345	299	346	300
rect	348	299	349	300
rect	354	299	355	300
rect	357	299	358	300
rect	360	299	361	300
rect	363	299	364	300
rect	366	299	367	300
rect	372	299	373	300
rect	375	299	376	300
rect	378	299	379	300
rect	384	299	385	300
rect	387	299	388	300
rect	390	299	391	300
rect	400	299	401	300
rect	4	300	5	301
rect	8	300	9	301
rect	14	300	15	301
rect	23	300	24	301
rect	39	300	40	301
rect	42	300	43	301
rect	51	300	52	301
rect	60	300	61	301
rect	63	300	64	301
rect	66	300	67	301
rect	69	300	70	301
rect	72	300	73	301
rect	81	300	82	301
rect	97	300	98	301
rect	100	300	101	301
rect	109	300	110	301
rect	112	300	113	301
rect	115	300	116	301
rect	118	300	119	301
rect	121	300	122	301
rect	124	300	125	301
rect	127	300	128	301
rect	134	300	135	301
rect	137	300	138	301
rect	139	300	140	301
rect	142	300	143	301
rect	145	300	146	301
rect	148	300	149	301
rect	158	300	159	301
rect	164	300	165	301
rect	167	300	168	301
rect	170	300	171	301
rect	176	300	177	301
rect	179	300	180	301
rect	182	300	183	301
rect	188	300	189	301
rect	191	300	192	301
rect	197	300	198	301
rect	200	300	201	301
rect	203	300	204	301
rect	206	300	207	301
rect	209	300	210	301
rect	224	300	225	301
rect	227	300	228	301
rect	230	300	231	301
rect	233	300	234	301
rect	242	300	243	301
rect	245	300	246	301
rect	251	300	252	301
rect	255	300	256	301
rect	271	300	272	301
rect	274	300	275	301
rect	277	300	278	301
rect	280	300	281	301
rect	289	300	290	301
rect	292	300	293	301
rect	308	300	309	301
rect	311	300	312	301
rect	324	300	325	301
rect	333	300	334	301
rect	336	300	337	301
rect	345	300	346	301
rect	348	300	349	301
rect	354	300	355	301
rect	357	300	358	301
rect	360	300	361	301
rect	363	300	364	301
rect	366	300	367	301
rect	372	300	373	301
rect	375	300	376	301
rect	378	300	379	301
rect	384	300	385	301
rect	387	300	388	301
rect	390	300	391	301
rect	400	300	401	301
rect	4	301	5	302
rect	8	301	9	302
rect	14	301	15	302
rect	23	301	24	302
rect	39	301	40	302
rect	42	301	43	302
rect	51	301	52	302
rect	60	301	61	302
rect	63	301	64	302
rect	66	301	67	302
rect	69	301	70	302
rect	72	301	73	302
rect	81	301	82	302
rect	97	301	98	302
rect	100	301	101	302
rect	109	301	110	302
rect	115	301	116	302
rect	118	301	119	302
rect	121	301	122	302
rect	124	301	125	302
rect	127	301	128	302
rect	134	301	135	302
rect	137	301	138	302
rect	139	301	140	302
rect	142	301	143	302
rect	145	301	146	302
rect	148	301	149	302
rect	158	301	159	302
rect	164	301	165	302
rect	167	301	168	302
rect	170	301	171	302
rect	179	301	180	302
rect	182	301	183	302
rect	188	301	189	302
rect	191	301	192	302
rect	197	301	198	302
rect	200	301	201	302
rect	203	301	204	302
rect	209	301	210	302
rect	224	301	225	302
rect	227	301	228	302
rect	230	301	231	302
rect	233	301	234	302
rect	242	301	243	302
rect	245	301	246	302
rect	251	301	252	302
rect	255	301	256	302
rect	271	301	272	302
rect	274	301	275	302
rect	277	301	278	302
rect	280	301	281	302
rect	289	301	290	302
rect	308	301	309	302
rect	311	301	312	302
rect	324	301	325	302
rect	333	301	334	302
rect	336	301	337	302
rect	345	301	346	302
rect	348	301	349	302
rect	354	301	355	302
rect	357	301	358	302
rect	360	301	361	302
rect	363	301	364	302
rect	366	301	367	302
rect	372	301	373	302
rect	375	301	376	302
rect	378	301	379	302
rect	384	301	385	302
rect	390	301	391	302
rect	400	301	401	302
rect	4	302	5	303
rect	8	302	9	303
rect	14	302	15	303
rect	23	302	24	303
rect	39	302	40	303
rect	42	302	43	303
rect	51	302	52	303
rect	60	302	61	303
rect	63	302	64	303
rect	66	302	67	303
rect	69	302	70	303
rect	72	302	73	303
rect	81	302	82	303
rect	97	302	98	303
rect	100	302	101	303
rect	109	302	110	303
rect	115	302	116	303
rect	118	302	119	303
rect	121	302	122	303
rect	124	302	125	303
rect	127	302	128	303
rect	131	302	132	303
rect	134	302	135	303
rect	137	302	138	303
rect	139	302	140	303
rect	142	302	143	303
rect	145	302	146	303
rect	148	302	149	303
rect	158	302	159	303
rect	164	302	165	303
rect	167	302	168	303
rect	170	302	171	303
rect	179	302	180	303
rect	182	302	183	303
rect	185	302	186	303
rect	188	302	189	303
rect	191	302	192	303
rect	197	302	198	303
rect	200	302	201	303
rect	203	302	204	303
rect	209	302	210	303
rect	221	302	222	303
rect	224	302	225	303
rect	227	302	228	303
rect	230	302	231	303
rect	233	302	234	303
rect	242	302	243	303
rect	245	302	246	303
rect	251	302	252	303
rect	255	302	256	303
rect	271	302	272	303
rect	274	302	275	303
rect	277	302	278	303
rect	280	302	281	303
rect	287	302	288	303
rect	289	302	290	303
rect	308	302	309	303
rect	311	302	312	303
rect	324	302	325	303
rect	333	302	334	303
rect	336	302	337	303
rect	345	302	346	303
rect	348	302	349	303
rect	354	302	355	303
rect	357	302	358	303
rect	360	302	361	303
rect	363	302	364	303
rect	366	302	367	303
rect	372	302	373	303
rect	375	302	376	303
rect	378	302	379	303
rect	384	302	385	303
rect	390	302	391	303
rect	394	302	395	303
rect	400	302	401	303
rect	4	303	5	304
rect	8	303	9	304
rect	14	303	15	304
rect	23	303	24	304
rect	39	303	40	304
rect	42	303	43	304
rect	51	303	52	304
rect	60	303	61	304
rect	63	303	64	304
rect	66	303	67	304
rect	69	303	70	304
rect	72	303	73	304
rect	81	303	82	304
rect	97	303	98	304
rect	100	303	101	304
rect	109	303	110	304
rect	115	303	116	304
rect	118	303	119	304
rect	121	303	122	304
rect	127	303	128	304
rect	131	303	132	304
rect	134	303	135	304
rect	137	303	138	304
rect	139	303	140	304
rect	142	303	143	304
rect	145	303	146	304
rect	148	303	149	304
rect	158	303	159	304
rect	164	303	165	304
rect	167	303	168	304
rect	170	303	171	304
rect	179	303	180	304
rect	182	303	183	304
rect	185	303	186	304
rect	191	303	192	304
rect	197	303	198	304
rect	203	303	204	304
rect	209	303	210	304
rect	221	303	222	304
rect	224	303	225	304
rect	227	303	228	304
rect	230	303	231	304
rect	233	303	234	304
rect	242	303	243	304
rect	245	303	246	304
rect	251	303	252	304
rect	255	303	256	304
rect	274	303	275	304
rect	277	303	278	304
rect	287	303	288	304
rect	289	303	290	304
rect	308	303	309	304
rect	311	303	312	304
rect	324	303	325	304
rect	333	303	334	304
rect	336	303	337	304
rect	345	303	346	304
rect	348	303	349	304
rect	354	303	355	304
rect	360	303	361	304
rect	363	303	364	304
rect	366	303	367	304
rect	372	303	373	304
rect	375	303	376	304
rect	378	303	379	304
rect	384	303	385	304
rect	390	303	391	304
rect	394	303	395	304
rect	400	303	401	304
rect	4	304	5	305
rect	8	304	9	305
rect	14	304	15	305
rect	23	304	24	305
rect	39	304	40	305
rect	42	304	43	305
rect	51	304	52	305
rect	60	304	61	305
rect	63	304	64	305
rect	66	304	67	305
rect	69	304	70	305
rect	72	304	73	305
rect	81	304	82	305
rect	97	304	98	305
rect	100	304	101	305
rect	109	304	110	305
rect	113	304	114	305
rect	115	304	116	305
rect	118	304	119	305
rect	121	304	122	305
rect	127	304	128	305
rect	131	304	132	305
rect	134	304	135	305
rect	137	304	138	305
rect	139	304	140	305
rect	142	304	143	305
rect	145	304	146	305
rect	148	304	149	305
rect	158	304	159	305
rect	164	304	165	305
rect	167	304	168	305
rect	170	304	171	305
rect	176	304	177	305
rect	179	304	180	305
rect	182	304	183	305
rect	185	304	186	305
rect	191	304	192	305
rect	197	304	198	305
rect	203	304	204	305
rect	209	304	210	305
rect	218	304	219	305
rect	221	304	222	305
rect	224	304	225	305
rect	227	304	228	305
rect	230	304	231	305
rect	233	304	234	305
rect	242	304	243	305
rect	245	304	246	305
rect	251	304	252	305
rect	255	304	256	305
rect	269	304	270	305
rect	274	304	275	305
rect	277	304	278	305
rect	287	304	288	305
rect	289	304	290	305
rect	293	304	294	305
rect	308	304	309	305
rect	311	304	312	305
rect	324	304	325	305
rect	333	304	334	305
rect	336	304	337	305
rect	345	304	346	305
rect	348	304	349	305
rect	354	304	355	305
rect	360	304	361	305
rect	363	304	364	305
rect	366	304	367	305
rect	372	304	373	305
rect	375	304	376	305
rect	378	304	379	305
rect	384	304	385	305
rect	388	304	389	305
rect	390	304	391	305
rect	394	304	395	305
rect	400	304	401	305
rect	4	305	5	306
rect	8	305	9	306
rect	14	305	15	306
rect	23	305	24	306
rect	39	305	40	306
rect	42	305	43	306
rect	51	305	52	306
rect	60	305	61	306
rect	63	305	64	306
rect	66	305	67	306
rect	69	305	70	306
rect	72	305	73	306
rect	81	305	82	306
rect	97	305	98	306
rect	100	305	101	306
rect	109	305	110	306
rect	113	305	114	306
rect	115	305	116	306
rect	118	305	119	306
rect	121	305	122	306
rect	131	305	132	306
rect	134	305	135	306
rect	137	305	138	306
rect	142	305	143	306
rect	145	305	146	306
rect	148	305	149	306
rect	158	305	159	306
rect	164	305	165	306
rect	167	305	168	306
rect	176	305	177	306
rect	179	305	180	306
rect	182	305	183	306
rect	185	305	186	306
rect	191	305	192	306
rect	203	305	204	306
rect	209	305	210	306
rect	218	305	219	306
rect	221	305	222	306
rect	224	305	225	306
rect	227	305	228	306
rect	230	305	231	306
rect	242	305	243	306
rect	245	305	246	306
rect	251	305	252	306
rect	255	305	256	306
rect	269	305	270	306
rect	274	305	275	306
rect	277	305	278	306
rect	287	305	288	306
rect	289	305	290	306
rect	293	305	294	306
rect	308	305	309	306
rect	311	305	312	306
rect	324	305	325	306
rect	333	305	334	306
rect	336	305	337	306
rect	345	305	346	306
rect	348	305	349	306
rect	354	305	355	306
rect	360	305	361	306
rect	366	305	367	306
rect	372	305	373	306
rect	375	305	376	306
rect	378	305	379	306
rect	384	305	385	306
rect	388	305	389	306
rect	390	305	391	306
rect	394	305	395	306
rect	400	305	401	306
rect	4	306	5	307
rect	8	306	9	307
rect	14	306	15	307
rect	23	306	24	307
rect	39	306	40	307
rect	42	306	43	307
rect	51	306	52	307
rect	60	306	61	307
rect	63	306	64	307
rect	66	306	67	307
rect	69	306	70	307
rect	72	306	73	307
rect	81	306	82	307
rect	97	306	98	307
rect	100	306	101	307
rect	109	306	110	307
rect	113	306	114	307
rect	115	306	116	307
rect	118	306	119	307
rect	121	306	122	307
rect	125	306	126	307
rect	131	306	132	307
rect	134	306	135	307
rect	137	306	138	307
rect	142	306	143	307
rect	145	306	146	307
rect	148	306	149	307
rect	152	306	153	307
rect	158	306	159	307
rect	164	306	165	307
rect	167	306	168	307
rect	176	306	177	307
rect	179	306	180	307
rect	182	306	183	307
rect	185	306	186	307
rect	188	306	189	307
rect	191	306	192	307
rect	203	306	204	307
rect	209	306	210	307
rect	215	306	216	307
rect	218	306	219	307
rect	221	306	222	307
rect	224	306	225	307
rect	227	306	228	307
rect	230	306	231	307
rect	242	306	243	307
rect	245	306	246	307
rect	251	306	252	307
rect	255	306	256	307
rect	269	306	270	307
rect	274	306	275	307
rect	277	306	278	307
rect	281	306	282	307
rect	287	306	288	307
rect	289	306	290	307
rect	293	306	294	307
rect	308	306	309	307
rect	311	306	312	307
rect	324	306	325	307
rect	333	306	334	307
rect	336	306	337	307
rect	345	306	346	307
rect	348	306	349	307
rect	354	306	355	307
rect	358	306	359	307
rect	360	306	361	307
rect	366	306	367	307
rect	372	306	373	307
rect	375	306	376	307
rect	378	306	379	307
rect	384	306	385	307
rect	388	306	389	307
rect	390	306	391	307
rect	394	306	395	307
rect	400	306	401	307
rect	4	307	5	308
rect	8	307	9	308
rect	14	307	15	308
rect	23	307	24	308
rect	39	307	40	308
rect	42	307	43	308
rect	51	307	52	308
rect	60	307	61	308
rect	63	307	64	308
rect	66	307	67	308
rect	69	307	70	308
rect	81	307	82	308
rect	97	307	98	308
rect	109	307	110	308
rect	113	307	114	308
rect	115	307	116	308
rect	118	307	119	308
rect	121	307	122	308
rect	125	307	126	308
rect	131	307	132	308
rect	134	307	135	308
rect	137	307	138	308
rect	142	307	143	308
rect	145	307	146	308
rect	152	307	153	308
rect	158	307	159	308
rect	167	307	168	308
rect	176	307	177	308
rect	179	307	180	308
rect	182	307	183	308
rect	185	307	186	308
rect	188	307	189	308
rect	203	307	204	308
rect	209	307	210	308
rect	215	307	216	308
rect	218	307	219	308
rect	221	307	222	308
rect	224	307	225	308
rect	227	307	228	308
rect	230	307	231	308
rect	242	307	243	308
rect	245	307	246	308
rect	251	307	252	308
rect	255	307	256	308
rect	269	307	270	308
rect	274	307	275	308
rect	277	307	278	308
rect	281	307	282	308
rect	287	307	288	308
rect	293	307	294	308
rect	308	307	309	308
rect	311	307	312	308
rect	324	307	325	308
rect	333	307	334	308
rect	336	307	337	308
rect	345	307	346	308
rect	354	307	355	308
rect	358	307	359	308
rect	366	307	367	308
rect	372	307	373	308
rect	375	307	376	308
rect	378	307	379	308
rect	384	307	385	308
rect	388	307	389	308
rect	390	307	391	308
rect	394	307	395	308
rect	400	307	401	308
rect	4	308	5	309
rect	8	308	9	309
rect	14	308	15	309
rect	23	308	24	309
rect	39	308	40	309
rect	42	308	43	309
rect	51	308	52	309
rect	60	308	61	309
rect	63	308	64	309
rect	66	308	67	309
rect	69	308	70	309
rect	81	308	82	309
rect	83	308	84	309
rect	95	308	96	309
rect	97	308	98	309
rect	109	308	110	309
rect	113	308	114	309
rect	115	308	116	309
rect	118	308	119	309
rect	121	308	122	309
rect	125	308	126	309
rect	128	308	129	309
rect	131	308	132	309
rect	134	308	135	309
rect	137	308	138	309
rect	142	308	143	309
rect	145	308	146	309
rect	152	308	153	309
rect	158	308	159	309
rect	167	308	168	309
rect	170	308	171	309
rect	176	308	177	309
rect	179	308	180	309
rect	182	308	183	309
rect	185	308	186	309
rect	188	308	189	309
rect	203	308	204	309
rect	206	308	207	309
rect	209	308	210	309
rect	215	308	216	309
rect	218	308	219	309
rect	221	308	222	309
rect	224	308	225	309
rect	227	308	228	309
rect	230	308	231	309
rect	233	308	234	309
rect	239	308	240	309
rect	242	308	243	309
rect	245	308	246	309
rect	251	308	252	309
rect	255	308	256	309
rect	269	308	270	309
rect	272	308	273	309
rect	274	308	275	309
rect	277	308	278	309
rect	281	308	282	309
rect	287	308	288	309
rect	293	308	294	309
rect	308	308	309	309
rect	311	308	312	309
rect	324	308	325	309
rect	333	308	334	309
rect	336	308	337	309
rect	345	308	346	309
rect	354	308	355	309
rect	358	308	359	309
rect	366	308	367	309
rect	372	308	373	309
rect	375	308	376	309
rect	378	308	379	309
rect	384	308	385	309
rect	388	308	389	309
rect	390	308	391	309
rect	394	308	395	309
rect	400	308	401	309
rect	4	309	5	310
rect	8	309	9	310
rect	14	309	15	310
rect	23	309	24	310
rect	39	309	40	310
rect	42	309	43	310
rect	51	309	52	310
rect	60	309	61	310
rect	63	309	64	310
rect	69	309	70	310
rect	81	309	82	310
rect	83	309	84	310
rect	95	309	96	310
rect	97	309	98	310
rect	113	309	114	310
rect	115	309	116	310
rect	118	309	119	310
rect	125	309	126	310
rect	128	309	129	310
rect	131	309	132	310
rect	134	309	135	310
rect	137	309	138	310
rect	142	309	143	310
rect	145	309	146	310
rect	152	309	153	310
rect	158	309	159	310
rect	167	309	168	310
rect	170	309	171	310
rect	176	309	177	310
rect	179	309	180	310
rect	182	309	183	310
rect	185	309	186	310
rect	188	309	189	310
rect	203	309	204	310
rect	206	309	207	310
rect	209	309	210	310
rect	215	309	216	310
rect	218	309	219	310
rect	221	309	222	310
rect	224	309	225	310
rect	227	309	228	310
rect	230	309	231	310
rect	233	309	234	310
rect	239	309	240	310
rect	242	309	243	310
rect	245	309	246	310
rect	251	309	252	310
rect	255	309	256	310
rect	269	309	270	310
rect	272	309	273	310
rect	274	309	275	310
rect	277	309	278	310
rect	281	309	282	310
rect	287	309	288	310
rect	293	309	294	310
rect	308	309	309	310
rect	311	309	312	310
rect	324	309	325	310
rect	333	309	334	310
rect	336	309	337	310
rect	345	309	346	310
rect	354	309	355	310
rect	358	309	359	310
rect	366	309	367	310
rect	372	309	373	310
rect	375	309	376	310
rect	378	309	379	310
rect	384	309	385	310
rect	388	309	389	310
rect	390	309	391	310
rect	394	309	395	310
rect	400	309	401	310
rect	4	310	5	311
rect	8	310	9	311
rect	14	310	15	311
rect	23	310	24	311
rect	39	310	40	311
rect	42	310	43	311
rect	51	310	52	311
rect	60	310	61	311
rect	63	310	64	311
rect	69	310	70	311
rect	77	310	78	311
rect	81	310	82	311
rect	83	310	84	311
rect	95	310	96	311
rect	97	310	98	311
rect	101	310	102	311
rect	113	310	114	311
rect	115	310	116	311
rect	118	310	119	311
rect	125	310	126	311
rect	128	310	129	311
rect	131	310	132	311
rect	134	310	135	311
rect	137	310	138	311
rect	142	310	143	311
rect	145	310	146	311
rect	152	310	153	311
rect	158	310	159	311
rect	167	310	168	311
rect	170	310	171	311
rect	176	310	177	311
rect	179	310	180	311
rect	182	310	183	311
rect	185	310	186	311
rect	188	310	189	311
rect	203	310	204	311
rect	206	310	207	311
rect	209	310	210	311
rect	215	310	216	311
rect	218	310	219	311
rect	221	310	222	311
rect	224	310	225	311
rect	227	310	228	311
rect	230	310	231	311
rect	233	310	234	311
rect	239	310	240	311
rect	242	310	243	311
rect	245	310	246	311
rect	251	310	252	311
rect	255	310	256	311
rect	269	310	270	311
rect	272	310	273	311
rect	274	310	275	311
rect	277	310	278	311
rect	281	310	282	311
rect	287	310	288	311
rect	293	310	294	311
rect	308	310	309	311
rect	311	310	312	311
rect	324	310	325	311
rect	333	310	334	311
rect	336	310	337	311
rect	345	310	346	311
rect	354	310	355	311
rect	358	310	359	311
rect	366	310	367	311
rect	372	310	373	311
rect	375	310	376	311
rect	378	310	379	311
rect	384	310	385	311
rect	388	310	389	311
rect	390	310	391	311
rect	394	310	395	311
rect	400	310	401	311
rect	413	310	414	311
rect	4	311	5	312
rect	8	311	9	312
rect	23	311	24	312
rect	39	311	40	312
rect	51	311	52	312
rect	60	311	61	312
rect	69	311	70	312
rect	77	311	78	312
rect	83	311	84	312
rect	97	311	98	312
rect	101	311	102	312
rect	113	311	114	312
rect	115	311	116	312
rect	118	311	119	312
rect	125	311	126	312
rect	128	311	129	312
rect	131	311	132	312
rect	134	311	135	312
rect	137	311	138	312
rect	152	311	153	312
rect	158	311	159	312
rect	167	311	168	312
rect	170	311	171	312
rect	176	311	177	312
rect	179	311	180	312
rect	185	311	186	312
rect	188	311	189	312
rect	203	311	204	312
rect	206	311	207	312
rect	209	311	210	312
rect	215	311	216	312
rect	218	311	219	312
rect	221	311	222	312
rect	227	311	228	312
rect	230	311	231	312
rect	233	311	234	312
rect	239	311	240	312
rect	242	311	243	312
rect	245	311	246	312
rect	251	311	252	312
rect	255	311	256	312
rect	269	311	270	312
rect	272	311	273	312
rect	274	311	275	312
rect	277	311	278	312
rect	281	311	282	312
rect	287	311	288	312
rect	293	311	294	312
rect	308	311	309	312
rect	311	311	312	312
rect	324	311	325	312
rect	333	311	334	312
rect	336	311	337	312
rect	345	311	346	312
rect	354	311	355	312
rect	358	311	359	312
rect	366	311	367	312
rect	372	311	373	312
rect	375	311	376	312
rect	384	311	385	312
rect	388	311	389	312
rect	390	311	391	312
rect	394	311	395	312
rect	400	311	401	312
rect	413	311	414	312
rect	1	312	2	313
rect	4	312	5	313
rect	8	312	9	313
rect	23	312	24	313
rect	39	312	40	313
rect	47	312	48	313
rect	51	312	52	313
rect	60	312	61	313
rect	69	312	70	313
rect	74	312	75	313
rect	77	312	78	313
rect	83	312	84	313
rect	92	312	93	313
rect	97	312	98	313
rect	101	312	102	313
rect	110	312	111	313
rect	113	312	114	313
rect	115	312	116	313
rect	118	312	119	313
rect	122	312	123	313
rect	125	312	126	313
rect	128	312	129	313
rect	131	312	132	313
rect	134	312	135	313
rect	137	312	138	313
rect	152	312	153	313
rect	155	312	156	313
rect	158	312	159	313
rect	161	312	162	313
rect	164	312	165	313
rect	167	312	168	313
rect	170	312	171	313
rect	176	312	177	313
rect	179	312	180	313
rect	185	312	186	313
rect	188	312	189	313
rect	200	312	201	313
rect	203	312	204	313
rect	206	312	207	313
rect	209	312	210	313
rect	215	312	216	313
rect	218	312	219	313
rect	221	312	222	313
rect	227	312	228	313
rect	230	312	231	313
rect	233	312	234	313
rect	239	312	240	313
rect	242	312	243	313
rect	245	312	246	313
rect	251	312	252	313
rect	255	312	256	313
rect	269	312	270	313
rect	272	312	273	313
rect	274	312	275	313
rect	277	312	278	313
rect	281	312	282	313
rect	287	312	288	313
rect	293	312	294	313
rect	308	312	309	313
rect	311	312	312	313
rect	324	312	325	313
rect	333	312	334	313
rect	336	312	337	313
rect	345	312	346	313
rect	354	312	355	313
rect	358	312	359	313
rect	361	312	362	313
rect	366	312	367	313
rect	372	312	373	313
rect	375	312	376	313
rect	379	312	380	313
rect	384	312	385	313
rect	388	312	389	313
rect	390	312	391	313
rect	394	312	395	313
rect	400	312	401	313
rect	413	312	414	313
rect	1	313	2	314
rect	47	313	48	314
rect	74	313	75	314
rect	77	313	78	314
rect	83	313	84	314
rect	92	313	93	314
rect	101	313	102	314
rect	110	313	111	314
rect	113	313	114	314
rect	122	313	123	314
rect	125	313	126	314
rect	128	313	129	314
rect	131	313	132	314
rect	134	313	135	314
rect	137	313	138	314
rect	152	313	153	314
rect	155	313	156	314
rect	161	313	162	314
rect	164	313	165	314
rect	167	313	168	314
rect	170	313	171	314
rect	176	313	177	314
rect	185	313	186	314
rect	188	313	189	314
rect	200	313	201	314
rect	203	313	204	314
rect	206	313	207	314
rect	215	313	216	314
rect	218	313	219	314
rect	221	313	222	314
rect	227	313	228	314
rect	233	313	234	314
rect	239	313	240	314
rect	242	313	243	314
rect	245	313	246	314
rect	251	313	252	314
rect	255	313	256	314
rect	269	313	270	314
rect	272	313	273	314
rect	274	313	275	314
rect	281	313	282	314
rect	287	313	288	314
rect	293	313	294	314
rect	308	313	309	314
rect	311	313	312	314
rect	324	313	325	314
rect	333	313	334	314
rect	345	313	346	314
rect	358	313	359	314
rect	361	313	362	314
rect	375	313	376	314
rect	379	313	380	314
rect	388	313	389	314
rect	394	313	395	314
rect	400	313	401	314
rect	413	313	414	314
rect	1	314	2	315
rect	14	314	15	315
rect	44	314	45	315
rect	47	314	48	315
rect	56	314	57	315
rect	65	314	66	315
rect	74	314	75	315
rect	77	314	78	315
rect	80	314	81	315
rect	83	314	84	315
rect	92	314	93	315
rect	101	314	102	315
rect	104	314	105	315
rect	107	314	108	315
rect	110	314	111	315
rect	113	314	114	315
rect	122	314	123	315
rect	125	314	126	315
rect	128	314	129	315
rect	131	314	132	315
rect	134	314	135	315
rect	137	314	138	315
rect	140	314	141	315
rect	146	314	147	315
rect	149	314	150	315
rect	152	314	153	315
rect	155	314	156	315
rect	161	314	162	315
rect	164	314	165	315
rect	167	314	168	315
rect	170	314	171	315
rect	173	314	174	315
rect	176	314	177	315
rect	185	314	186	315
rect	188	314	189	315
rect	197	314	198	315
rect	200	314	201	315
rect	203	314	204	315
rect	206	314	207	315
rect	215	314	216	315
rect	218	314	219	315
rect	221	314	222	315
rect	224	314	225	315
rect	227	314	228	315
rect	233	314	234	315
rect	236	314	237	315
rect	239	314	240	315
rect	242	314	243	315
rect	245	314	246	315
rect	251	314	252	315
rect	255	314	256	315
rect	269	314	270	315
rect	272	314	273	315
rect	274	314	275	315
rect	281	314	282	315
rect	287	314	288	315
rect	290	314	291	315
rect	293	314	294	315
rect	308	314	309	315
rect	311	314	312	315
rect	324	314	325	315
rect	333	314	334	315
rect	335	314	336	315
rect	345	314	346	315
rect	358	314	359	315
rect	361	314	362	315
rect	375	314	376	315
rect	379	314	380	315
rect	388	314	389	315
rect	394	314	395	315
rect	400	314	401	315
rect	410	314	411	315
rect	413	314	414	315
rect	1	315	2	316
rect	14	315	15	316
rect	44	315	45	316
rect	47	315	48	316
rect	56	315	57	316
rect	65	315	66	316
rect	74	315	75	316
rect	77	315	78	316
rect	80	315	81	316
rect	83	315	84	316
rect	92	315	93	316
rect	101	315	102	316
rect	104	315	105	316
rect	107	315	108	316
rect	110	315	111	316
rect	113	315	114	316
rect	122	315	123	316
rect	125	315	126	316
rect	128	315	129	316
rect	131	315	132	316
rect	134	315	135	316
rect	137	315	138	316
rect	140	315	141	316
rect	146	315	147	316
rect	149	315	150	316
rect	152	315	153	316
rect	155	315	156	316
rect	161	315	162	316
rect	164	315	165	316
rect	167	315	168	316
rect	170	315	171	316
rect	173	315	174	316
rect	176	315	177	316
rect	185	315	186	316
rect	188	315	189	316
rect	197	315	198	316
rect	200	315	201	316
rect	203	315	204	316
rect	206	315	207	316
rect	215	315	216	316
rect	218	315	219	316
rect	221	315	222	316
rect	224	315	225	316
rect	233	315	234	316
rect	236	315	237	316
rect	239	315	240	316
rect	242	315	243	316
rect	245	315	246	316
rect	251	315	252	316
rect	269	315	270	316
rect	272	315	273	316
rect	281	315	282	316
rect	287	315	288	316
rect	290	315	291	316
rect	293	315	294	316
rect	335	315	336	316
rect	358	315	359	316
rect	361	315	362	316
rect	379	315	380	316
rect	388	315	389	316
rect	394	315	395	316
rect	410	315	411	316
rect	413	315	414	316
rect	1	316	2	317
rect	4	316	5	317
rect	14	316	15	317
rect	44	316	45	317
rect	47	316	48	317
rect	56	316	57	317
rect	65	316	66	317
rect	74	316	75	317
rect	77	316	78	317
rect	80	316	81	317
rect	83	316	84	317
rect	92	316	93	317
rect	101	316	102	317
rect	104	316	105	317
rect	107	316	108	317
rect	110	316	111	317
rect	113	316	114	317
rect	122	316	123	317
rect	125	316	126	317
rect	128	316	129	317
rect	131	316	132	317
rect	134	316	135	317
rect	137	316	138	317
rect	140	316	141	317
rect	146	316	147	317
rect	149	316	150	317
rect	152	316	153	317
rect	155	316	156	317
rect	161	316	162	317
rect	164	316	165	317
rect	167	316	168	317
rect	170	316	171	317
rect	173	316	174	317
rect	176	316	177	317
rect	185	316	186	317
rect	188	316	189	317
rect	197	316	198	317
rect	200	316	201	317
rect	203	316	204	317
rect	206	316	207	317
rect	212	316	213	317
rect	215	316	216	317
rect	218	316	219	317
rect	221	316	222	317
rect	224	316	225	317
rect	233	316	234	317
rect	236	316	237	317
rect	239	316	240	317
rect	242	316	243	317
rect	245	316	246	317
rect	248	316	249	317
rect	251	316	252	317
rect	260	316	261	317
rect	269	316	270	317
rect	272	316	273	317
rect	281	316	282	317
rect	284	316	285	317
rect	287	316	288	317
rect	290	316	291	317
rect	293	316	294	317
rect	323	316	324	317
rect	332	316	333	317
rect	335	316	336	317
rect	358	316	359	317
rect	361	316	362	317
rect	370	316	371	317
rect	379	316	380	317
rect	388	316	389	317
rect	391	316	392	317
rect	394	316	395	317
rect	410	316	411	317
rect	413	316	414	317
rect	419	316	420	317
rect	14	323	15	324
rect	44	323	45	324
rect	47	323	48	324
rect	56	323	57	324
rect	65	323	66	324
rect	74	323	75	324
rect	77	323	78	324
rect	80	323	81	324
rect	83	323	84	324
rect	92	323	93	324
rect	101	323	102	324
rect	104	323	105	324
rect	107	323	108	324
rect	110	323	111	324
rect	113	323	114	324
rect	116	323	117	324
rect	122	323	123	324
rect	125	323	126	324
rect	128	323	129	324
rect	131	323	132	324
rect	134	323	135	324
rect	137	323	138	324
rect	140	323	141	324
rect	149	323	150	324
rect	152	323	153	324
rect	155	323	156	324
rect	164	323	165	324
rect	167	323	168	324
rect	170	323	171	324
rect	173	323	174	324
rect	176	323	177	324
rect	179	323	180	324
rect	185	323	186	324
rect	188	323	189	324
rect	191	323	192	324
rect	197	323	198	324
rect	200	323	201	324
rect	203	323	204	324
rect	206	323	207	324
rect	215	323	216	324
rect	218	323	219	324
rect	221	323	222	324
rect	224	323	225	324
rect	230	323	231	324
rect	233	323	234	324
rect	236	323	237	324
rect	245	323	246	324
rect	248	323	249	324
rect	251	323	252	324
rect	260	323	261	324
rect	269	323	270	324
rect	272	323	273	324
rect	281	323	282	324
rect	284	323	285	324
rect	287	323	288	324
rect	290	323	291	324
rect	293	323	294	324
rect	323	323	324	324
rect	332	323	333	324
rect	335	323	336	324
rect	338	323	339	324
rect	348	323	349	324
rect	358	323	359	324
rect	361	323	362	324
rect	370	323	371	324
rect	376	323	377	324
rect	379	323	380	324
rect	382	323	383	324
rect	388	323	389	324
rect	391	323	392	324
rect	394	323	395	324
rect	400	323	401	324
rect	410	323	411	324
rect	416	323	417	324
rect	419	323	420	324
rect	14	324	15	325
rect	44	324	45	325
rect	47	324	48	325
rect	56	324	57	325
rect	65	324	66	325
rect	74	324	75	325
rect	77	324	78	325
rect	80	324	81	325
rect	83	324	84	325
rect	92	324	93	325
rect	101	324	102	325
rect	104	324	105	325
rect	107	324	108	325
rect	110	324	111	325
rect	113	324	114	325
rect	116	324	117	325
rect	122	324	123	325
rect	125	324	126	325
rect	128	324	129	325
rect	131	324	132	325
rect	134	324	135	325
rect	137	324	138	325
rect	140	324	141	325
rect	149	324	150	325
rect	152	324	153	325
rect	155	324	156	325
rect	164	324	165	325
rect	167	324	168	325
rect	170	324	171	325
rect	173	324	174	325
rect	176	324	177	325
rect	179	324	180	325
rect	185	324	186	325
rect	188	324	189	325
rect	191	324	192	325
rect	197	324	198	325
rect	200	324	201	325
rect	203	324	204	325
rect	206	324	207	325
rect	215	324	216	325
rect	218	324	219	325
rect	221	324	222	325
rect	224	324	225	325
rect	233	324	234	325
rect	236	324	237	325
rect	245	324	246	325
rect	248	324	249	325
rect	251	324	252	325
rect	260	324	261	325
rect	269	324	270	325
rect	272	324	273	325
rect	281	324	282	325
rect	284	324	285	325
rect	287	324	288	325
rect	290	324	291	325
rect	293	324	294	325
rect	323	324	324	325
rect	332	324	333	325
rect	335	324	336	325
rect	338	324	339	325
rect	348	324	349	325
rect	358	324	359	325
rect	361	324	362	325
rect	370	324	371	325
rect	376	324	377	325
rect	379	324	380	325
rect	382	324	383	325
rect	388	324	389	325
rect	391	324	392	325
rect	394	324	395	325
rect	400	324	401	325
rect	410	324	411	325
rect	416	324	417	325
rect	419	324	420	325
rect	14	325	15	326
rect	44	325	45	326
rect	47	325	48	326
rect	56	325	57	326
rect	65	325	66	326
rect	74	325	75	326
rect	77	325	78	326
rect	80	325	81	326
rect	83	325	84	326
rect	92	325	93	326
rect	101	325	102	326
rect	104	325	105	326
rect	107	325	108	326
rect	110	325	111	326
rect	113	325	114	326
rect	116	325	117	326
rect	122	325	123	326
rect	125	325	126	326
rect	128	325	129	326
rect	131	325	132	326
rect	134	325	135	326
rect	137	325	138	326
rect	140	325	141	326
rect	149	325	150	326
rect	152	325	153	326
rect	155	325	156	326
rect	164	325	165	326
rect	167	325	168	326
rect	170	325	171	326
rect	173	325	174	326
rect	176	325	177	326
rect	179	325	180	326
rect	185	325	186	326
rect	188	325	189	326
rect	191	325	192	326
rect	197	325	198	326
rect	200	325	201	326
rect	203	325	204	326
rect	206	325	207	326
rect	213	325	214	326
rect	215	325	216	326
rect	218	325	219	326
rect	221	325	222	326
rect	224	325	225	326
rect	233	325	234	326
rect	236	325	237	326
rect	245	325	246	326
rect	248	325	249	326
rect	251	325	252	326
rect	260	325	261	326
rect	269	325	270	326
rect	272	325	273	326
rect	281	325	282	326
rect	284	325	285	326
rect	287	325	288	326
rect	290	325	291	326
rect	293	325	294	326
rect	323	325	324	326
rect	332	325	333	326
rect	335	325	336	326
rect	338	325	339	326
rect	348	325	349	326
rect	358	325	359	326
rect	361	325	362	326
rect	370	325	371	326
rect	376	325	377	326
rect	379	325	380	326
rect	382	325	383	326
rect	388	325	389	326
rect	391	325	392	326
rect	394	325	395	326
rect	400	325	401	326
rect	410	325	411	326
rect	416	325	417	326
rect	419	325	420	326
rect	14	326	15	327
rect	44	326	45	327
rect	47	326	48	327
rect	56	326	57	327
rect	65	326	66	327
rect	74	326	75	327
rect	77	326	78	327
rect	80	326	81	327
rect	83	326	84	327
rect	92	326	93	327
rect	101	326	102	327
rect	104	326	105	327
rect	107	326	108	327
rect	110	326	111	327
rect	113	326	114	327
rect	116	326	117	327
rect	122	326	123	327
rect	125	326	126	327
rect	128	326	129	327
rect	131	326	132	327
rect	134	326	135	327
rect	137	326	138	327
rect	140	326	141	327
rect	149	326	150	327
rect	152	326	153	327
rect	155	326	156	327
rect	164	326	165	327
rect	167	326	168	327
rect	170	326	171	327
rect	173	326	174	327
rect	176	326	177	327
rect	179	326	180	327
rect	185	326	186	327
rect	188	326	189	327
rect	191	326	192	327
rect	197	326	198	327
rect	200	326	201	327
rect	203	326	204	327
rect	206	326	207	327
rect	213	326	214	327
rect	215	326	216	327
rect	218	326	219	327
rect	221	326	222	327
rect	224	326	225	327
rect	233	326	234	327
rect	245	326	246	327
rect	248	326	249	327
rect	251	326	252	327
rect	260	326	261	327
rect	269	326	270	327
rect	272	326	273	327
rect	281	326	282	327
rect	284	326	285	327
rect	287	326	288	327
rect	290	326	291	327
rect	293	326	294	327
rect	323	326	324	327
rect	332	326	333	327
rect	335	326	336	327
rect	338	326	339	327
rect	348	326	349	327
rect	358	326	359	327
rect	361	326	362	327
rect	370	326	371	327
rect	376	326	377	327
rect	379	326	380	327
rect	382	326	383	327
rect	388	326	389	327
rect	391	326	392	327
rect	394	326	395	327
rect	400	326	401	327
rect	410	326	411	327
rect	416	326	417	327
rect	419	326	420	327
rect	14	327	15	328
rect	44	327	45	328
rect	47	327	48	328
rect	56	327	57	328
rect	65	327	66	328
rect	74	327	75	328
rect	77	327	78	328
rect	80	327	81	328
rect	83	327	84	328
rect	92	327	93	328
rect	101	327	102	328
rect	104	327	105	328
rect	107	327	108	328
rect	110	327	111	328
rect	113	327	114	328
rect	116	327	117	328
rect	122	327	123	328
rect	125	327	126	328
rect	128	327	129	328
rect	131	327	132	328
rect	134	327	135	328
rect	137	327	138	328
rect	140	327	141	328
rect	149	327	150	328
rect	152	327	153	328
rect	155	327	156	328
rect	164	327	165	328
rect	167	327	168	328
rect	170	327	171	328
rect	173	327	174	328
rect	176	327	177	328
rect	179	327	180	328
rect	185	327	186	328
rect	188	327	189	328
rect	191	327	192	328
rect	197	327	198	328
rect	200	327	201	328
rect	203	327	204	328
rect	206	327	207	328
rect	213	327	214	328
rect	215	327	216	328
rect	218	327	219	328
rect	221	327	222	328
rect	224	327	225	328
rect	229	327	230	328
rect	233	327	234	328
rect	245	327	246	328
rect	248	327	249	328
rect	251	327	252	328
rect	260	327	261	328
rect	269	327	270	328
rect	272	327	273	328
rect	281	327	282	328
rect	284	327	285	328
rect	287	327	288	328
rect	290	327	291	328
rect	293	327	294	328
rect	323	327	324	328
rect	332	327	333	328
rect	335	327	336	328
rect	338	327	339	328
rect	348	327	349	328
rect	358	327	359	328
rect	361	327	362	328
rect	370	327	371	328
rect	376	327	377	328
rect	379	327	380	328
rect	382	327	383	328
rect	388	327	389	328
rect	391	327	392	328
rect	394	327	395	328
rect	400	327	401	328
rect	410	327	411	328
rect	416	327	417	328
rect	419	327	420	328
rect	14	328	15	329
rect	44	328	45	329
rect	47	328	48	329
rect	56	328	57	329
rect	65	328	66	329
rect	74	328	75	329
rect	77	328	78	329
rect	80	328	81	329
rect	83	328	84	329
rect	92	328	93	329
rect	101	328	102	329
rect	104	328	105	329
rect	107	328	108	329
rect	110	328	111	329
rect	113	328	114	329
rect	116	328	117	329
rect	122	328	123	329
rect	125	328	126	329
rect	128	328	129	329
rect	131	328	132	329
rect	134	328	135	329
rect	137	328	138	329
rect	140	328	141	329
rect	149	328	150	329
rect	152	328	153	329
rect	155	328	156	329
rect	164	328	165	329
rect	167	328	168	329
rect	170	328	171	329
rect	176	328	177	329
rect	179	328	180	329
rect	185	328	186	329
rect	188	328	189	329
rect	191	328	192	329
rect	197	328	198	329
rect	200	328	201	329
rect	203	328	204	329
rect	206	328	207	329
rect	215	328	216	329
rect	218	328	219	329
rect	221	328	222	329
rect	224	328	225	329
rect	229	328	230	329
rect	233	328	234	329
rect	245	328	246	329
rect	248	328	249	329
rect	251	328	252	329
rect	260	328	261	329
rect	269	328	270	329
rect	272	328	273	329
rect	281	328	282	329
rect	284	328	285	329
rect	287	328	288	329
rect	290	328	291	329
rect	323	328	324	329
rect	332	328	333	329
rect	335	328	336	329
rect	338	328	339	329
rect	358	328	359	329
rect	361	328	362	329
rect	370	328	371	329
rect	376	328	377	329
rect	379	328	380	329
rect	382	328	383	329
rect	388	328	389	329
rect	391	328	392	329
rect	394	328	395	329
rect	400	328	401	329
rect	410	328	411	329
rect	416	328	417	329
rect	419	328	420	329
rect	14	329	15	330
rect	44	329	45	330
rect	47	329	48	330
rect	56	329	57	330
rect	65	329	66	330
rect	74	329	75	330
rect	77	329	78	330
rect	80	329	81	330
rect	83	329	84	330
rect	92	329	93	330
rect	101	329	102	330
rect	104	329	105	330
rect	107	329	108	330
rect	110	329	111	330
rect	113	329	114	330
rect	116	329	117	330
rect	122	329	123	330
rect	125	329	126	330
rect	128	329	129	330
rect	131	329	132	330
rect	134	329	135	330
rect	137	329	138	330
rect	140	329	141	330
rect	147	329	148	330
rect	149	329	150	330
rect	152	329	153	330
rect	155	329	156	330
rect	164	329	165	330
rect	167	329	168	330
rect	170	329	171	330
rect	176	329	177	330
rect	179	329	180	330
rect	185	329	186	330
rect	188	329	189	330
rect	191	329	192	330
rect	197	329	198	330
rect	200	329	201	330
rect	203	329	204	330
rect	206	329	207	330
rect	215	329	216	330
rect	218	329	219	330
rect	221	329	222	330
rect	224	329	225	330
rect	229	329	230	330
rect	233	329	234	330
rect	235	329	236	330
rect	245	329	246	330
rect	248	329	249	330
rect	251	329	252	330
rect	260	329	261	330
rect	269	329	270	330
rect	272	329	273	330
rect	281	329	282	330
rect	284	329	285	330
rect	287	329	288	330
rect	290	329	291	330
rect	323	329	324	330
rect	332	329	333	330
rect	335	329	336	330
rect	338	329	339	330
rect	358	329	359	330
rect	361	329	362	330
rect	370	329	371	330
rect	376	329	377	330
rect	379	329	380	330
rect	382	329	383	330
rect	388	329	389	330
rect	391	329	392	330
rect	394	329	395	330
rect	400	329	401	330
rect	410	329	411	330
rect	416	329	417	330
rect	419	329	420	330
rect	14	330	15	331
rect	44	330	45	331
rect	47	330	48	331
rect	56	330	57	331
rect	65	330	66	331
rect	74	330	75	331
rect	77	330	78	331
rect	80	330	81	331
rect	83	330	84	331
rect	92	330	93	331
rect	101	330	102	331
rect	104	330	105	331
rect	107	330	108	331
rect	110	330	111	331
rect	113	330	114	331
rect	116	330	117	331
rect	122	330	123	331
rect	125	330	126	331
rect	128	330	129	331
rect	131	330	132	331
rect	134	330	135	331
rect	137	330	138	331
rect	140	330	141	331
rect	147	330	148	331
rect	149	330	150	331
rect	152	330	153	331
rect	155	330	156	331
rect	164	330	165	331
rect	167	330	168	331
rect	170	330	171	331
rect	176	330	177	331
rect	179	330	180	331
rect	185	330	186	331
rect	188	330	189	331
rect	197	330	198	331
rect	200	330	201	331
rect	203	330	204	331
rect	206	330	207	331
rect	215	330	216	331
rect	218	330	219	331
rect	221	330	222	331
rect	224	330	225	331
rect	229	330	230	331
rect	235	330	236	331
rect	245	330	246	331
rect	248	330	249	331
rect	251	330	252	331
rect	260	330	261	331
rect	269	330	270	331
rect	272	330	273	331
rect	281	330	282	331
rect	284	330	285	331
rect	287	330	288	331
rect	290	330	291	331
rect	332	330	333	331
rect	335	330	336	331
rect	338	330	339	331
rect	358	330	359	331
rect	370	330	371	331
rect	376	330	377	331
rect	379	330	380	331
rect	382	330	383	331
rect	388	330	389	331
rect	391	330	392	331
rect	394	330	395	331
rect	400	330	401	331
rect	410	330	411	331
rect	416	330	417	331
rect	419	330	420	331
rect	14	331	15	332
rect	44	331	45	332
rect	47	331	48	332
rect	56	331	57	332
rect	65	331	66	332
rect	74	331	75	332
rect	77	331	78	332
rect	80	331	81	332
rect	83	331	84	332
rect	92	331	93	332
rect	101	331	102	332
rect	104	331	105	332
rect	107	331	108	332
rect	110	331	111	332
rect	113	331	114	332
rect	116	331	117	332
rect	122	331	123	332
rect	125	331	126	332
rect	128	331	129	332
rect	131	331	132	332
rect	134	331	135	332
rect	137	331	138	332
rect	140	331	141	332
rect	147	331	148	332
rect	149	331	150	332
rect	152	331	153	332
rect	155	331	156	332
rect	164	331	165	332
rect	167	331	168	332
rect	170	331	171	332
rect	174	331	175	332
rect	176	331	177	332
rect	179	331	180	332
rect	185	331	186	332
rect	188	331	189	332
rect	197	331	198	332
rect	200	331	201	332
rect	203	331	204	332
rect	206	331	207	332
rect	215	331	216	332
rect	218	331	219	332
rect	221	331	222	332
rect	224	331	225	332
rect	226	331	227	332
rect	229	331	230	332
rect	235	331	236	332
rect	245	331	246	332
rect	248	331	249	332
rect	251	331	252	332
rect	260	331	261	332
rect	269	331	270	332
rect	272	331	273	332
rect	281	331	282	332
rect	284	331	285	332
rect	287	331	288	332
rect	290	331	291	332
rect	305	331	306	332
rect	332	331	333	332
rect	335	331	336	332
rect	338	331	339	332
rect	349	331	350	332
rect	358	331	359	332
rect	370	331	371	332
rect	376	331	377	332
rect	379	331	380	332
rect	382	331	383	332
rect	388	331	389	332
rect	391	331	392	332
rect	394	331	395	332
rect	400	331	401	332
rect	410	331	411	332
rect	416	331	417	332
rect	419	331	420	332
rect	14	332	15	333
rect	44	332	45	333
rect	47	332	48	333
rect	56	332	57	333
rect	65	332	66	333
rect	74	332	75	333
rect	77	332	78	333
rect	80	332	81	333
rect	83	332	84	333
rect	92	332	93	333
rect	101	332	102	333
rect	104	332	105	333
rect	107	332	108	333
rect	110	332	111	333
rect	113	332	114	333
rect	116	332	117	333
rect	122	332	123	333
rect	125	332	126	333
rect	128	332	129	333
rect	131	332	132	333
rect	134	332	135	333
rect	137	332	138	333
rect	140	332	141	333
rect	147	332	148	333
rect	149	332	150	333
rect	152	332	153	333
rect	155	332	156	333
rect	164	332	165	333
rect	167	332	168	333
rect	170	332	171	333
rect	174	332	175	333
rect	176	332	177	333
rect	179	332	180	333
rect	185	332	186	333
rect	188	332	189	333
rect	197	332	198	333
rect	203	332	204	333
rect	206	332	207	333
rect	215	332	216	333
rect	218	332	219	333
rect	221	332	222	333
rect	224	332	225	333
rect	226	332	227	333
rect	229	332	230	333
rect	235	332	236	333
rect	245	332	246	333
rect	251	332	252	333
rect	269	332	270	333
rect	272	332	273	333
rect	281	332	282	333
rect	284	332	285	333
rect	287	332	288	333
rect	290	332	291	333
rect	305	332	306	333
rect	332	332	333	333
rect	335	332	336	333
rect	338	332	339	333
rect	349	332	350	333
rect	358	332	359	333
rect	370	332	371	333
rect	376	332	377	333
rect	379	332	380	333
rect	382	332	383	333
rect	388	332	389	333
rect	391	332	392	333
rect	394	332	395	333
rect	400	332	401	333
rect	410	332	411	333
rect	416	332	417	333
rect	419	332	420	333
rect	14	333	15	334
rect	44	333	45	334
rect	47	333	48	334
rect	56	333	57	334
rect	65	333	66	334
rect	74	333	75	334
rect	77	333	78	334
rect	80	333	81	334
rect	83	333	84	334
rect	92	333	93	334
rect	101	333	102	334
rect	104	333	105	334
rect	107	333	108	334
rect	110	333	111	334
rect	113	333	114	334
rect	116	333	117	334
rect	122	333	123	334
rect	125	333	126	334
rect	128	333	129	334
rect	131	333	132	334
rect	134	333	135	334
rect	137	333	138	334
rect	140	333	141	334
rect	147	333	148	334
rect	149	333	150	334
rect	152	333	153	334
rect	155	333	156	334
rect	164	333	165	334
rect	167	333	168	334
rect	170	333	171	334
rect	174	333	175	334
rect	176	333	177	334
rect	179	333	180	334
rect	185	333	186	334
rect	188	333	189	334
rect	192	333	193	334
rect	197	333	198	334
rect	203	333	204	334
rect	206	333	207	334
rect	215	333	216	334
rect	218	333	219	334
rect	221	333	222	334
rect	224	333	225	334
rect	226	333	227	334
rect	229	333	230	334
rect	232	333	233	334
rect	235	333	236	334
rect	245	333	246	334
rect	251	333	252	334
rect	256	333	257	334
rect	269	333	270	334
rect	272	333	273	334
rect	281	333	282	334
rect	284	333	285	334
rect	287	333	288	334
rect	290	333	291	334
rect	305	333	306	334
rect	323	333	324	334
rect	332	333	333	334
rect	335	333	336	334
rect	338	333	339	334
rect	349	333	350	334
rect	358	333	359	334
rect	361	333	362	334
rect	370	333	371	334
rect	376	333	377	334
rect	379	333	380	334
rect	382	333	383	334
rect	388	333	389	334
rect	391	333	392	334
rect	394	333	395	334
rect	400	333	401	334
rect	410	333	411	334
rect	416	333	417	334
rect	419	333	420	334
rect	14	334	15	335
rect	44	334	45	335
rect	47	334	48	335
rect	56	334	57	335
rect	65	334	66	335
rect	74	334	75	335
rect	77	334	78	335
rect	80	334	81	335
rect	83	334	84	335
rect	92	334	93	335
rect	101	334	102	335
rect	104	334	105	335
rect	107	334	108	335
rect	110	334	111	335
rect	113	334	114	335
rect	116	334	117	335
rect	122	334	123	335
rect	125	334	126	335
rect	128	334	129	335
rect	131	334	132	335
rect	134	334	135	335
rect	137	334	138	335
rect	140	334	141	335
rect	147	334	148	335
rect	149	334	150	335
rect	152	334	153	335
rect	155	334	156	335
rect	164	334	165	335
rect	167	334	168	335
rect	170	334	171	335
rect	174	334	175	335
rect	176	334	177	335
rect	179	334	180	335
rect	185	334	186	335
rect	188	334	189	335
rect	192	334	193	335
rect	197	334	198	335
rect	203	334	204	335
rect	206	334	207	335
rect	218	334	219	335
rect	221	334	222	335
rect	224	334	225	335
rect	226	334	227	335
rect	229	334	230	335
rect	232	334	233	335
rect	235	334	236	335
rect	251	334	252	335
rect	256	334	257	335
rect	272	334	273	335
rect	284	334	285	335
rect	287	334	288	335
rect	290	334	291	335
rect	305	334	306	335
rect	323	334	324	335
rect	335	334	336	335
rect	338	334	339	335
rect	349	334	350	335
rect	361	334	362	335
rect	370	334	371	335
rect	376	334	377	335
rect	379	334	380	335
rect	382	334	383	335
rect	388	334	389	335
rect	391	334	392	335
rect	394	334	395	335
rect	400	334	401	335
rect	410	334	411	335
rect	416	334	417	335
rect	419	334	420	335
rect	14	335	15	336
rect	44	335	45	336
rect	47	335	48	336
rect	56	335	57	336
rect	65	335	66	336
rect	74	335	75	336
rect	77	335	78	336
rect	80	335	81	336
rect	83	335	84	336
rect	92	335	93	336
rect	101	335	102	336
rect	104	335	105	336
rect	107	335	108	336
rect	110	335	111	336
rect	113	335	114	336
rect	116	335	117	336
rect	122	335	123	336
rect	125	335	126	336
rect	128	335	129	336
rect	131	335	132	336
rect	134	335	135	336
rect	137	335	138	336
rect	140	335	141	336
rect	147	335	148	336
rect	149	335	150	336
rect	152	335	153	336
rect	155	335	156	336
rect	164	335	165	336
rect	167	335	168	336
rect	170	335	171	336
rect	174	335	175	336
rect	176	335	177	336
rect	179	335	180	336
rect	185	335	186	336
rect	188	335	189	336
rect	192	335	193	336
rect	197	335	198	336
rect	201	335	202	336
rect	203	335	204	336
rect	206	335	207	336
rect	218	335	219	336
rect	221	335	222	336
rect	224	335	225	336
rect	226	335	227	336
rect	229	335	230	336
rect	232	335	233	336
rect	235	335	236	336
rect	247	335	248	336
rect	251	335	252	336
rect	256	335	257	336
rect	259	335	260	336
rect	272	335	273	336
rect	277	335	278	336
rect	284	335	285	336
rect	287	335	288	336
rect	290	335	291	336
rect	305	335	306	336
rect	320	335	321	336
rect	323	335	324	336
rect	335	335	336	336
rect	338	335	339	336
rect	346	335	347	336
rect	349	335	350	336
rect	361	335	362	336
rect	370	335	371	336
rect	376	335	377	336
rect	379	335	380	336
rect	382	335	383	336
rect	388	335	389	336
rect	391	335	392	336
rect	394	335	395	336
rect	400	335	401	336
rect	410	335	411	336
rect	416	335	417	336
rect	419	335	420	336
rect	14	336	15	337
rect	44	336	45	337
rect	47	336	48	337
rect	56	336	57	337
rect	65	336	66	337
rect	74	336	75	337
rect	77	336	78	337
rect	80	336	81	337
rect	83	336	84	337
rect	92	336	93	337
rect	101	336	102	337
rect	104	336	105	337
rect	107	336	108	337
rect	110	336	111	337
rect	113	336	114	337
rect	116	336	117	337
rect	122	336	123	337
rect	125	336	126	337
rect	128	336	129	337
rect	134	336	135	337
rect	137	336	138	337
rect	140	336	141	337
rect	147	336	148	337
rect	149	336	150	337
rect	152	336	153	337
rect	155	336	156	337
rect	164	336	165	337
rect	167	336	168	337
rect	170	336	171	337
rect	174	336	175	337
rect	176	336	177	337
rect	179	336	180	337
rect	185	336	186	337
rect	188	336	189	337
rect	192	336	193	337
rect	197	336	198	337
rect	201	336	202	337
rect	203	336	204	337
rect	206	336	207	337
rect	218	336	219	337
rect	221	336	222	337
rect	224	336	225	337
rect	226	336	227	337
rect	229	336	230	337
rect	232	336	233	337
rect	235	336	236	337
rect	247	336	248	337
rect	251	336	252	337
rect	256	336	257	337
rect	259	336	260	337
rect	272	336	273	337
rect	277	336	278	337
rect	284	336	285	337
rect	287	336	288	337
rect	290	336	291	337
rect	305	336	306	337
rect	320	336	321	337
rect	323	336	324	337
rect	335	336	336	337
rect	338	336	339	337
rect	346	336	347	337
rect	349	336	350	337
rect	361	336	362	337
rect	370	336	371	337
rect	376	336	377	337
rect	391	336	392	337
rect	394	336	395	337
rect	400	336	401	337
rect	410	336	411	337
rect	416	336	417	337
rect	419	336	420	337
rect	14	337	15	338
rect	44	337	45	338
rect	47	337	48	338
rect	56	337	57	338
rect	65	337	66	338
rect	74	337	75	338
rect	77	337	78	338
rect	80	337	81	338
rect	83	337	84	338
rect	92	337	93	338
rect	101	337	102	338
rect	104	337	105	338
rect	107	337	108	338
rect	110	337	111	338
rect	113	337	114	338
rect	116	337	117	338
rect	122	337	123	338
rect	125	337	126	338
rect	128	337	129	338
rect	134	337	135	338
rect	137	337	138	338
rect	140	337	141	338
rect	147	337	148	338
rect	149	337	150	338
rect	152	337	153	338
rect	155	337	156	338
rect	164	337	165	338
rect	167	337	168	338
rect	170	337	171	338
rect	174	337	175	338
rect	176	337	177	338
rect	179	337	180	338
rect	185	337	186	338
rect	188	337	189	338
rect	192	337	193	338
rect	197	337	198	338
rect	201	337	202	338
rect	203	337	204	338
rect	206	337	207	338
rect	218	337	219	338
rect	221	337	222	338
rect	224	337	225	338
rect	226	337	227	338
rect	229	337	230	338
rect	232	337	233	338
rect	235	337	236	338
rect	247	337	248	338
rect	251	337	252	338
rect	256	337	257	338
rect	259	337	260	338
rect	272	337	273	338
rect	277	337	278	338
rect	284	337	285	338
rect	287	337	288	338
rect	290	337	291	338
rect	305	337	306	338
rect	320	337	321	338
rect	323	337	324	338
rect	333	337	334	338
rect	335	337	336	338
rect	338	337	339	338
rect	346	337	347	338
rect	349	337	350	338
rect	358	337	359	338
rect	361	337	362	338
rect	370	337	371	338
rect	376	337	377	338
rect	391	337	392	338
rect	394	337	395	338
rect	400	337	401	338
rect	410	337	411	338
rect	416	337	417	338
rect	419	337	420	338
rect	14	338	15	339
rect	44	338	45	339
rect	47	338	48	339
rect	56	338	57	339
rect	65	338	66	339
rect	74	338	75	339
rect	77	338	78	339
rect	80	338	81	339
rect	92	338	93	339
rect	101	338	102	339
rect	104	338	105	339
rect	107	338	108	339
rect	110	338	111	339
rect	113	338	114	339
rect	116	338	117	339
rect	122	338	123	339
rect	125	338	126	339
rect	128	338	129	339
rect	134	338	135	339
rect	137	338	138	339
rect	140	338	141	339
rect	147	338	148	339
rect	149	338	150	339
rect	155	338	156	339
rect	164	338	165	339
rect	167	338	168	339
rect	174	338	175	339
rect	176	338	177	339
rect	179	338	180	339
rect	185	338	186	339
rect	188	338	189	339
rect	192	338	193	339
rect	197	338	198	339
rect	201	338	202	339
rect	218	338	219	339
rect	221	338	222	339
rect	224	338	225	339
rect	226	338	227	339
rect	229	338	230	339
rect	232	338	233	339
rect	235	338	236	339
rect	247	338	248	339
rect	251	338	252	339
rect	256	338	257	339
rect	259	338	260	339
rect	272	338	273	339
rect	277	338	278	339
rect	284	338	285	339
rect	287	338	288	339
rect	290	338	291	339
rect	305	338	306	339
rect	320	338	321	339
rect	323	338	324	339
rect	333	338	334	339
rect	335	338	336	339
rect	338	338	339	339
rect	346	338	347	339
rect	349	338	350	339
rect	358	338	359	339
rect	361	338	362	339
rect	370	338	371	339
rect	376	338	377	339
rect	391	338	392	339
rect	394	338	395	339
rect	400	338	401	339
rect	416	338	417	339
rect	419	338	420	339
rect	14	339	15	340
rect	44	339	45	340
rect	47	339	48	340
rect	56	339	57	340
rect	65	339	66	340
rect	74	339	75	340
rect	77	339	78	340
rect	80	339	81	340
rect	87	339	88	340
rect	92	339	93	340
rect	101	339	102	340
rect	104	339	105	340
rect	107	339	108	340
rect	110	339	111	340
rect	113	339	114	340
rect	116	339	117	340
rect	122	339	123	340
rect	125	339	126	340
rect	128	339	129	340
rect	132	339	133	340
rect	134	339	135	340
rect	137	339	138	340
rect	140	339	141	340
rect	147	339	148	340
rect	149	339	150	340
rect	155	339	156	340
rect	164	339	165	340
rect	167	339	168	340
rect	174	339	175	340
rect	176	339	177	340
rect	179	339	180	340
rect	183	339	184	340
rect	185	339	186	340
rect	188	339	189	340
rect	192	339	193	340
rect	195	339	196	340
rect	197	339	198	340
rect	201	339	202	340
rect	210	339	211	340
rect	216	339	217	340
rect	218	339	219	340
rect	221	339	222	340
rect	224	339	225	340
rect	226	339	227	340
rect	229	339	230	340
rect	232	339	233	340
rect	235	339	236	340
rect	247	339	248	340
rect	251	339	252	340
rect	256	339	257	340
rect	259	339	260	340
rect	272	339	273	340
rect	277	339	278	340
rect	284	339	285	340
rect	287	339	288	340
rect	290	339	291	340
rect	305	339	306	340
rect	320	339	321	340
rect	323	339	324	340
rect	333	339	334	340
rect	335	339	336	340
rect	338	339	339	340
rect	346	339	347	340
rect	349	339	350	340
rect	358	339	359	340
rect	361	339	362	340
rect	370	339	371	340
rect	376	339	377	340
rect	391	339	392	340
rect	394	339	395	340
rect	400	339	401	340
rect	416	339	417	340
rect	419	339	420	340
rect	14	340	15	341
rect	44	340	45	341
rect	47	340	48	341
rect	56	340	57	341
rect	65	340	66	341
rect	74	340	75	341
rect	77	340	78	341
rect	87	340	88	341
rect	92	340	93	341
rect	101	340	102	341
rect	107	340	108	341
rect	110	340	111	341
rect	116	340	117	341
rect	122	340	123	341
rect	125	340	126	341
rect	128	340	129	341
rect	132	340	133	341
rect	134	340	135	341
rect	137	340	138	341
rect	140	340	141	341
rect	147	340	148	341
rect	164	340	165	341
rect	167	340	168	341
rect	174	340	175	341
rect	176	340	177	341
rect	179	340	180	341
rect	183	340	184	341
rect	185	340	186	341
rect	188	340	189	341
rect	192	340	193	341
rect	195	340	196	341
rect	201	340	202	341
rect	210	340	211	341
rect	216	340	217	341
rect	218	340	219	341
rect	224	340	225	341
rect	226	340	227	341
rect	229	340	230	341
rect	232	340	233	341
rect	235	340	236	341
rect	247	340	248	341
rect	256	340	257	341
rect	259	340	260	341
rect	272	340	273	341
rect	277	340	278	341
rect	284	340	285	341
rect	290	340	291	341
rect	305	340	306	341
rect	320	340	321	341
rect	323	340	324	341
rect	333	340	334	341
rect	335	340	336	341
rect	338	340	339	341
rect	346	340	347	341
rect	349	340	350	341
rect	358	340	359	341
rect	361	340	362	341
rect	370	340	371	341
rect	376	340	377	341
rect	391	340	392	341
rect	394	340	395	341
rect	400	340	401	341
rect	416	340	417	341
rect	419	340	420	341
rect	14	341	15	342
rect	44	341	45	342
rect	47	341	48	342
rect	56	341	57	342
rect	65	341	66	342
rect	74	341	75	342
rect	77	341	78	342
rect	84	341	85	342
rect	87	341	88	342
rect	92	341	93	342
rect	99	341	100	342
rect	101	341	102	342
rect	107	341	108	342
rect	110	341	111	342
rect	114	341	115	342
rect	116	341	117	342
rect	122	341	123	342
rect	125	341	126	342
rect	128	341	129	342
rect	132	341	133	342
rect	134	341	135	342
rect	137	341	138	342
rect	140	341	141	342
rect	144	341	145	342
rect	147	341	148	342
rect	153	341	154	342
rect	164	341	165	342
rect	167	341	168	342
rect	171	341	172	342
rect	174	341	175	342
rect	176	341	177	342
rect	179	341	180	342
rect	183	341	184	342
rect	185	341	186	342
rect	188	341	189	342
rect	192	341	193	342
rect	195	341	196	342
rect	201	341	202	342
rect	207	341	208	342
rect	210	341	211	342
rect	216	341	217	342
rect	218	341	219	342
rect	224	341	225	342
rect	226	341	227	342
rect	229	341	230	342
rect	232	341	233	342
rect	235	341	236	342
rect	244	341	245	342
rect	247	341	248	342
rect	256	341	257	342
rect	259	341	260	342
rect	268	341	269	342
rect	272	341	273	342
rect	277	341	278	342
rect	284	341	285	342
rect	290	341	291	342
rect	305	341	306	342
rect	311	341	312	342
rect	320	341	321	342
rect	323	341	324	342
rect	333	341	334	342
rect	335	341	336	342
rect	338	341	339	342
rect	346	341	347	342
rect	349	341	350	342
rect	358	341	359	342
rect	361	341	362	342
rect	370	341	371	342
rect	376	341	377	342
rect	382	341	383	342
rect	391	341	392	342
rect	394	341	395	342
rect	400	341	401	342
rect	416	341	417	342
rect	419	341	420	342
rect	14	342	15	343
rect	44	342	45	343
rect	47	342	48	343
rect	56	342	57	343
rect	65	342	66	343
rect	74	342	75	343
rect	77	342	78	343
rect	84	342	85	343
rect	87	342	88	343
rect	92	342	93	343
rect	99	342	100	343
rect	107	342	108	343
rect	110	342	111	343
rect	114	342	115	343
rect	116	342	117	343
rect	125	342	126	343
rect	128	342	129	343
rect	132	342	133	343
rect	137	342	138	343
rect	140	342	141	343
rect	144	342	145	343
rect	147	342	148	343
rect	153	342	154	343
rect	164	342	165	343
rect	167	342	168	343
rect	171	342	172	343
rect	174	342	175	343
rect	176	342	177	343
rect	179	342	180	343
rect	183	342	184	343
rect	185	342	186	343
rect	188	342	189	343
rect	192	342	193	343
rect	195	342	196	343
rect	201	342	202	343
rect	207	342	208	343
rect	210	342	211	343
rect	216	342	217	343
rect	218	342	219	343
rect	224	342	225	343
rect	226	342	227	343
rect	229	342	230	343
rect	232	342	233	343
rect	235	342	236	343
rect	244	342	245	343
rect	247	342	248	343
rect	256	342	257	343
rect	259	342	260	343
rect	268	342	269	343
rect	272	342	273	343
rect	277	342	278	343
rect	284	342	285	343
rect	290	342	291	343
rect	305	342	306	343
rect	311	342	312	343
rect	320	342	321	343
rect	323	342	324	343
rect	333	342	334	343
rect	335	342	336	343
rect	338	342	339	343
rect	346	342	347	343
rect	349	342	350	343
rect	358	342	359	343
rect	361	342	362	343
rect	370	342	371	343
rect	376	342	377	343
rect	382	342	383	343
rect	391	342	392	343
rect	394	342	395	343
rect	400	342	401	343
rect	416	342	417	343
rect	419	342	420	343
rect	14	343	15	344
rect	44	343	45	344
rect	47	343	48	344
rect	56	343	57	344
rect	65	343	66	344
rect	72	343	73	344
rect	74	343	75	344
rect	77	343	78	344
rect	84	343	85	344
rect	87	343	88	344
rect	92	343	93	344
rect	99	343	100	344
rect	105	343	106	344
rect	107	343	108	344
rect	110	343	111	344
rect	114	343	115	344
rect	116	343	117	344
rect	125	343	126	344
rect	128	343	129	344
rect	132	343	133	344
rect	137	343	138	344
rect	140	343	141	344
rect	144	343	145	344
rect	147	343	148	344
rect	153	343	154	344
rect	164	343	165	344
rect	167	343	168	344
rect	171	343	172	344
rect	174	343	175	344
rect	176	343	177	344
rect	179	343	180	344
rect	183	343	184	344
rect	185	343	186	344
rect	188	343	189	344
rect	192	343	193	344
rect	195	343	196	344
rect	201	343	202	344
rect	207	343	208	344
rect	210	343	211	344
rect	216	343	217	344
rect	218	343	219	344
rect	224	343	225	344
rect	226	343	227	344
rect	229	343	230	344
rect	232	343	233	344
rect	235	343	236	344
rect	244	343	245	344
rect	247	343	248	344
rect	256	343	257	344
rect	259	343	260	344
rect	268	343	269	344
rect	272	343	273	344
rect	277	343	278	344
rect	284	343	285	344
rect	290	343	291	344
rect	305	343	306	344
rect	311	343	312	344
rect	320	343	321	344
rect	323	343	324	344
rect	333	343	334	344
rect	335	343	336	344
rect	338	343	339	344
rect	346	343	347	344
rect	349	343	350	344
rect	358	343	359	344
rect	361	343	362	344
rect	370	343	371	344
rect	376	343	377	344
rect	378	343	379	344
rect	382	343	383	344
rect	391	343	392	344
rect	394	343	395	344
rect	400	343	401	344
rect	416	343	417	344
rect	419	343	420	344
rect	14	344	15	345
rect	44	344	45	345
rect	47	344	48	345
rect	56	344	57	345
rect	65	344	66	345
rect	72	344	73	345
rect	74	344	75	345
rect	84	344	85	345
rect	87	344	88	345
rect	92	344	93	345
rect	99	344	100	345
rect	105	344	106	345
rect	114	344	115	345
rect	116	344	117	345
rect	125	344	126	345
rect	132	344	133	345
rect	137	344	138	345
rect	140	344	141	345
rect	144	344	145	345
rect	147	344	148	345
rect	153	344	154	345
rect	164	344	165	345
rect	167	344	168	345
rect	171	344	172	345
rect	174	344	175	345
rect	179	344	180	345
rect	183	344	184	345
rect	185	344	186	345
rect	188	344	189	345
rect	192	344	193	345
rect	195	344	196	345
rect	201	344	202	345
rect	207	344	208	345
rect	210	344	211	345
rect	216	344	217	345
rect	226	344	227	345
rect	229	344	230	345
rect	232	344	233	345
rect	235	344	236	345
rect	244	344	245	345
rect	247	344	248	345
rect	256	344	257	345
rect	259	344	260	345
rect	268	344	269	345
rect	272	344	273	345
rect	277	344	278	345
rect	284	344	285	345
rect	290	344	291	345
rect	305	344	306	345
rect	311	344	312	345
rect	320	344	321	345
rect	323	344	324	345
rect	333	344	334	345
rect	335	344	336	345
rect	338	344	339	345
rect	346	344	347	345
rect	349	344	350	345
rect	358	344	359	345
rect	361	344	362	345
rect	370	344	371	345
rect	376	344	377	345
rect	378	344	379	345
rect	382	344	383	345
rect	391	344	392	345
rect	394	344	395	345
rect	400	344	401	345
rect	416	344	417	345
rect	419	344	420	345
rect	14	345	15	346
rect	44	345	45	346
rect	47	345	48	346
rect	56	345	57	346
rect	65	345	66	346
rect	72	345	73	346
rect	74	345	75	346
rect	81	345	82	346
rect	84	345	85	346
rect	87	345	88	346
rect	92	345	93	346
rect	99	345	100	346
rect	102	345	103	346
rect	105	345	106	346
rect	114	345	115	346
rect	116	345	117	346
rect	123	345	124	346
rect	125	345	126	346
rect	132	345	133	346
rect	135	345	136	346
rect	137	345	138	346
rect	140	345	141	346
rect	144	345	145	346
rect	147	345	148	346
rect	150	345	151	346
rect	153	345	154	346
rect	164	345	165	346
rect	167	345	168	346
rect	171	345	172	346
rect	174	345	175	346
rect	179	345	180	346
rect	183	345	184	346
rect	185	345	186	346
rect	188	345	189	346
rect	192	345	193	346
rect	195	345	196	346
rect	201	345	202	346
rect	204	345	205	346
rect	207	345	208	346
rect	210	345	211	346
rect	216	345	217	346
rect	226	345	227	346
rect	229	345	230	346
rect	232	345	233	346
rect	235	345	236	346
rect	244	345	245	346
rect	247	345	248	346
rect	256	345	257	346
rect	259	345	260	346
rect	268	345	269	346
rect	272	345	273	346
rect	277	345	278	346
rect	284	345	285	346
rect	290	345	291	346
rect	305	345	306	346
rect	311	345	312	346
rect	320	345	321	346
rect	323	345	324	346
rect	333	345	334	346
rect	335	345	336	346
rect	338	345	339	346
rect	343	345	344	346
rect	346	345	347	346
rect	349	345	350	346
rect	358	345	359	346
rect	361	345	362	346
rect	370	345	371	346
rect	376	345	377	346
rect	378	345	379	346
rect	382	345	383	346
rect	391	345	392	346
rect	394	345	395	346
rect	400	345	401	346
rect	416	345	417	346
rect	419	345	420	346
rect	14	346	15	347
rect	44	346	45	347
rect	56	346	57	347
rect	72	346	73	347
rect	74	346	75	347
rect	81	346	82	347
rect	84	346	85	347
rect	87	346	88	347
rect	92	346	93	347
rect	99	346	100	347
rect	102	346	103	347
rect	105	346	106	347
rect	114	346	115	347
rect	123	346	124	347
rect	132	346	133	347
rect	135	346	136	347
rect	137	346	138	347
rect	144	346	145	347
rect	147	346	148	347
rect	150	346	151	347
rect	153	346	154	347
rect	164	346	165	347
rect	171	346	172	347
rect	174	346	175	347
rect	183	346	184	347
rect	185	346	186	347
rect	188	346	189	347
rect	192	346	193	347
rect	195	346	196	347
rect	201	346	202	347
rect	204	346	205	347
rect	207	346	208	347
rect	210	346	211	347
rect	216	346	217	347
rect	226	346	227	347
rect	229	346	230	347
rect	232	346	233	347
rect	235	346	236	347
rect	244	346	245	347
rect	247	346	248	347
rect	256	346	257	347
rect	259	346	260	347
rect	268	346	269	347
rect	277	346	278	347
rect	305	346	306	347
rect	311	346	312	347
rect	320	346	321	347
rect	323	346	324	347
rect	333	346	334	347
rect	338	346	339	347
rect	343	346	344	347
rect	346	346	347	347
rect	349	346	350	347
rect	358	346	359	347
rect	361	346	362	347
rect	370	346	371	347
rect	376	346	377	347
rect	378	346	379	347
rect	382	346	383	347
rect	391	346	392	347
rect	400	346	401	347
rect	416	346	417	347
rect	419	346	420	347
rect	14	347	15	348
rect	44	347	45	348
rect	54	347	55	348
rect	56	347	57	348
rect	72	347	73	348
rect	74	347	75	348
rect	78	347	79	348
rect	81	347	82	348
rect	84	347	85	348
rect	87	347	88	348
rect	92	347	93	348
rect	96	347	97	348
rect	99	347	100	348
rect	102	347	103	348
rect	105	347	106	348
rect	114	347	115	348
rect	123	347	124	348
rect	126	347	127	348
rect	132	347	133	348
rect	135	347	136	348
rect	137	347	138	348
rect	144	347	145	348
rect	147	347	148	348
rect	150	347	151	348
rect	153	347	154	348
rect	156	347	157	348
rect	164	347	165	348
rect	168	347	169	348
rect	171	347	172	348
rect	174	347	175	348
rect	180	347	181	348
rect	183	347	184	348
rect	185	347	186	348
rect	188	347	189	348
rect	192	347	193	348
rect	195	347	196	348
rect	198	347	199	348
rect	201	347	202	348
rect	204	347	205	348
rect	207	347	208	348
rect	210	347	211	348
rect	216	347	217	348
rect	226	347	227	348
rect	229	347	230	348
rect	232	347	233	348
rect	235	347	236	348
rect	244	347	245	348
rect	247	347	248	348
rect	256	347	257	348
rect	259	347	260	348
rect	268	347	269	348
rect	277	347	278	348
rect	280	347	281	348
rect	289	347	290	348
rect	305	347	306	348
rect	308	347	309	348
rect	311	347	312	348
rect	320	347	321	348
rect	323	347	324	348
rect	333	347	334	348
rect	338	347	339	348
rect	343	347	344	348
rect	346	347	347	348
rect	349	347	350	348
rect	358	347	359	348
rect	361	347	362	348
rect	370	347	371	348
rect	376	347	377	348
rect	378	347	379	348
rect	382	347	383	348
rect	391	347	392	348
rect	395	347	396	348
rect	400	347	401	348
rect	416	347	417	348
rect	419	347	420	348
rect	54	348	55	349
rect	72	348	73	349
rect	78	348	79	349
rect	81	348	82	349
rect	84	348	85	349
rect	87	348	88	349
rect	96	348	97	349
rect	99	348	100	349
rect	102	348	103	349
rect	105	348	106	349
rect	114	348	115	349
rect	123	348	124	349
rect	126	348	127	349
rect	132	348	133	349
rect	135	348	136	349
rect	144	348	145	349
rect	147	348	148	349
rect	150	348	151	349
rect	153	348	154	349
rect	156	348	157	349
rect	168	348	169	349
rect	171	348	172	349
rect	174	348	175	349
rect	180	348	181	349
rect	183	348	184	349
rect	192	348	193	349
rect	195	348	196	349
rect	198	348	199	349
rect	201	348	202	349
rect	204	348	205	349
rect	207	348	208	349
rect	210	348	211	349
rect	216	348	217	349
rect	226	348	227	349
rect	229	348	230	349
rect	232	348	233	349
rect	235	348	236	349
rect	244	348	245	349
rect	247	348	248	349
rect	256	348	257	349
rect	259	348	260	349
rect	268	348	269	349
rect	277	348	278	349
rect	280	348	281	349
rect	289	348	290	349
rect	305	348	306	349
rect	308	348	309	349
rect	311	348	312	349
rect	320	348	321	349
rect	323	348	324	349
rect	333	348	334	349
rect	343	348	344	349
rect	346	348	347	349
rect	349	348	350	349
rect	358	348	359	349
rect	361	348	362	349
rect	378	348	379	349
rect	382	348	383	349
rect	395	348	396	349
rect	7	349	8	350
rect	51	349	52	350
rect	54	349	55	350
rect	63	349	64	350
rect	72	349	73	350
rect	75	349	76	350
rect	78	349	79	350
rect	81	349	82	350
rect	84	349	85	350
rect	87	349	88	350
rect	96	349	97	350
rect	99	349	100	350
rect	102	349	103	350
rect	105	349	106	350
rect	114	349	115	350
rect	123	349	124	350
rect	126	349	127	350
rect	129	349	130	350
rect	132	349	133	350
rect	135	349	136	350
rect	138	349	139	350
rect	144	349	145	350
rect	147	349	148	350
rect	150	349	151	350
rect	153	349	154	350
rect	156	349	157	350
rect	165	349	166	350
rect	168	349	169	350
rect	171	349	172	350
rect	174	349	175	350
rect	177	349	178	350
rect	180	349	181	350
rect	183	349	184	350
rect	192	349	193	350
rect	195	349	196	350
rect	198	349	199	350
rect	201	349	202	350
rect	204	349	205	350
rect	207	349	208	350
rect	210	349	211	350
rect	216	349	217	350
rect	226	349	227	350
rect	229	349	230	350
rect	232	349	233	350
rect	235	349	236	350
rect	244	349	245	350
rect	247	349	248	350
rect	256	349	257	350
rect	259	349	260	350
rect	268	349	269	350
rect	277	349	278	350
rect	280	349	281	350
rect	289	349	290	350
rect	305	349	306	350
rect	308	349	309	350
rect	311	349	312	350
rect	320	349	321	350
rect	323	349	324	350
rect	333	349	334	350
rect	343	349	344	350
rect	346	349	347	350
rect	349	349	350	350
rect	358	349	359	350
rect	361	349	362	350
rect	378	349	379	350
rect	382	349	383	350
rect	395	349	396	350
rect	4	356	5	357
rect	7	356	8	357
rect	10	356	11	357
rect	20	356	21	357
rect	51	356	52	357
rect	54	356	55	357
rect	63	356	64	357
rect	72	356	73	357
rect	75	356	76	357
rect	78	356	79	357
rect	81	356	82	357
rect	84	356	85	357
rect	87	356	88	357
rect	96	356	97	357
rect	99	356	100	357
rect	102	356	103	357
rect	105	356	106	357
rect	114	356	115	357
rect	123	356	124	357
rect	132	356	133	357
rect	135	356	136	357
rect	138	356	139	357
rect	147	356	148	357
rect	150	356	151	357
rect	153	356	154	357
rect	156	356	157	357
rect	159	356	160	357
rect	165	356	166	357
rect	168	356	169	357
rect	171	356	172	357
rect	174	356	175	357
rect	177	356	178	357
rect	180	356	181	357
rect	183	356	184	357
rect	186	356	187	357
rect	192	356	193	357
rect	195	356	196	357
rect	204	356	205	357
rect	207	356	208	357
rect	210	356	211	357
rect	213	356	214	357
rect	223	356	224	357
rect	226	356	227	357
rect	229	356	230	357
rect	232	356	233	357
rect	235	356	236	357
rect	244	356	245	357
rect	247	356	248	357
rect	256	356	257	357
rect	259	356	260	357
rect	268	356	269	357
rect	277	356	278	357
rect	280	356	281	357
rect	289	356	290	357
rect	305	356	306	357
rect	308	356	309	357
rect	311	356	312	357
rect	320	356	321	357
rect	323	356	324	357
rect	326	356	327	357
rect	346	356	347	357
rect	349	356	350	357
rect	358	356	359	357
rect	371	356	372	357
rect	375	356	376	357
rect	392	356	393	357
rect	395	356	396	357
rect	4	357	5	358
rect	7	357	8	358
rect	10	357	11	358
rect	20	357	21	358
rect	51	357	52	358
rect	54	357	55	358
rect	63	357	64	358
rect	72	357	73	358
rect	75	357	76	358
rect	78	357	79	358
rect	81	357	82	358
rect	84	357	85	358
rect	87	357	88	358
rect	96	357	97	358
rect	99	357	100	358
rect	102	357	103	358
rect	105	357	106	358
rect	114	357	115	358
rect	123	357	124	358
rect	132	357	133	358
rect	135	357	136	358
rect	138	357	139	358
rect	147	357	148	358
rect	150	357	151	358
rect	153	357	154	358
rect	156	357	157	358
rect	168	357	169	358
rect	171	357	172	358
rect	174	357	175	358
rect	177	357	178	358
rect	180	357	181	358
rect	183	357	184	358
rect	186	357	187	358
rect	192	357	193	358
rect	195	357	196	358
rect	204	357	205	358
rect	207	357	208	358
rect	210	357	211	358
rect	213	357	214	358
rect	223	357	224	358
rect	226	357	227	358
rect	229	357	230	358
rect	232	357	233	358
rect	235	357	236	358
rect	244	357	245	358
rect	247	357	248	358
rect	256	357	257	358
rect	259	357	260	358
rect	268	357	269	358
rect	277	357	278	358
rect	280	357	281	358
rect	289	357	290	358
rect	305	357	306	358
rect	308	357	309	358
rect	311	357	312	358
rect	320	357	321	358
rect	323	357	324	358
rect	326	357	327	358
rect	346	357	347	358
rect	349	357	350	358
rect	358	357	359	358
rect	371	357	372	358
rect	375	357	376	358
rect	392	357	393	358
rect	395	357	396	358
rect	4	358	5	359
rect	7	358	8	359
rect	10	358	11	359
rect	20	358	21	359
rect	51	358	52	359
rect	54	358	55	359
rect	63	358	64	359
rect	72	358	73	359
rect	75	358	76	359
rect	78	358	79	359
rect	81	358	82	359
rect	84	358	85	359
rect	87	358	88	359
rect	96	358	97	359
rect	99	358	100	359
rect	102	358	103	359
rect	105	358	106	359
rect	114	358	115	359
rect	123	358	124	359
rect	132	358	133	359
rect	135	358	136	359
rect	138	358	139	359
rect	147	358	148	359
rect	150	358	151	359
rect	153	358	154	359
rect	156	358	157	359
rect	168	358	169	359
rect	171	358	172	359
rect	174	358	175	359
rect	177	358	178	359
rect	180	358	181	359
rect	183	358	184	359
rect	186	358	187	359
rect	192	358	193	359
rect	195	358	196	359
rect	204	358	205	359
rect	207	358	208	359
rect	210	358	211	359
rect	213	358	214	359
rect	223	358	224	359
rect	226	358	227	359
rect	229	358	230	359
rect	232	358	233	359
rect	235	358	236	359
rect	244	358	245	359
rect	247	358	248	359
rect	256	358	257	359
rect	259	358	260	359
rect	268	358	269	359
rect	277	358	278	359
rect	280	358	281	359
rect	289	358	290	359
rect	305	358	306	359
rect	308	358	309	359
rect	311	358	312	359
rect	320	358	321	359
rect	323	358	324	359
rect	326	358	327	359
rect	346	358	347	359
rect	349	358	350	359
rect	358	358	359	359
rect	371	358	372	359
rect	375	358	376	359
rect	392	358	393	359
rect	395	358	396	359
rect	4	359	5	360
rect	7	359	8	360
rect	10	359	11	360
rect	20	359	21	360
rect	51	359	52	360
rect	54	359	55	360
rect	63	359	64	360
rect	72	359	73	360
rect	75	359	76	360
rect	78	359	79	360
rect	81	359	82	360
rect	84	359	85	360
rect	87	359	88	360
rect	96	359	97	360
rect	99	359	100	360
rect	102	359	103	360
rect	105	359	106	360
rect	114	359	115	360
rect	123	359	124	360
rect	132	359	133	360
rect	135	359	136	360
rect	138	359	139	360
rect	147	359	148	360
rect	150	359	151	360
rect	153	359	154	360
rect	168	359	169	360
rect	171	359	172	360
rect	174	359	175	360
rect	177	359	178	360
rect	180	359	181	360
rect	183	359	184	360
rect	186	359	187	360
rect	192	359	193	360
rect	195	359	196	360
rect	204	359	205	360
rect	207	359	208	360
rect	210	359	211	360
rect	213	359	214	360
rect	223	359	224	360
rect	226	359	227	360
rect	229	359	230	360
rect	232	359	233	360
rect	235	359	236	360
rect	244	359	245	360
rect	247	359	248	360
rect	256	359	257	360
rect	259	359	260	360
rect	268	359	269	360
rect	277	359	278	360
rect	280	359	281	360
rect	289	359	290	360
rect	305	359	306	360
rect	308	359	309	360
rect	311	359	312	360
rect	320	359	321	360
rect	323	359	324	360
rect	326	359	327	360
rect	346	359	347	360
rect	349	359	350	360
rect	358	359	359	360
rect	371	359	372	360
rect	375	359	376	360
rect	392	359	393	360
rect	395	359	396	360
rect	4	360	5	361
rect	7	360	8	361
rect	10	360	11	361
rect	20	360	21	361
rect	51	360	52	361
rect	54	360	55	361
rect	63	360	64	361
rect	72	360	73	361
rect	75	360	76	361
rect	78	360	79	361
rect	81	360	82	361
rect	84	360	85	361
rect	87	360	88	361
rect	96	360	97	361
rect	99	360	100	361
rect	102	360	103	361
rect	105	360	106	361
rect	114	360	115	361
rect	123	360	124	361
rect	132	360	133	361
rect	135	360	136	361
rect	138	360	139	361
rect	147	360	148	361
rect	150	360	151	361
rect	153	360	154	361
rect	168	360	169	361
rect	171	360	172	361
rect	174	360	175	361
rect	177	360	178	361
rect	180	360	181	361
rect	183	360	184	361
rect	186	360	187	361
rect	192	360	193	361
rect	195	360	196	361
rect	204	360	205	361
rect	207	360	208	361
rect	210	360	211	361
rect	213	360	214	361
rect	223	360	224	361
rect	226	360	227	361
rect	229	360	230	361
rect	232	360	233	361
rect	235	360	236	361
rect	244	360	245	361
rect	247	360	248	361
rect	256	360	257	361
rect	259	360	260	361
rect	268	360	269	361
rect	274	360	275	361
rect	277	360	278	361
rect	280	360	281	361
rect	289	360	290	361
rect	305	360	306	361
rect	308	360	309	361
rect	311	360	312	361
rect	320	360	321	361
rect	323	360	324	361
rect	326	360	327	361
rect	346	360	347	361
rect	349	360	350	361
rect	358	360	359	361
rect	371	360	372	361
rect	375	360	376	361
rect	392	360	393	361
rect	395	360	396	361
rect	4	361	5	362
rect	7	361	8	362
rect	10	361	11	362
rect	20	361	21	362
rect	51	361	52	362
rect	54	361	55	362
rect	63	361	64	362
rect	72	361	73	362
rect	75	361	76	362
rect	78	361	79	362
rect	81	361	82	362
rect	84	361	85	362
rect	87	361	88	362
rect	96	361	97	362
rect	102	361	103	362
rect	105	361	106	362
rect	114	361	115	362
rect	123	361	124	362
rect	135	361	136	362
rect	138	361	139	362
rect	147	361	148	362
rect	150	361	151	362
rect	153	361	154	362
rect	168	361	169	362
rect	171	361	172	362
rect	174	361	175	362
rect	177	361	178	362
rect	180	361	181	362
rect	186	361	187	362
rect	192	361	193	362
rect	195	361	196	362
rect	204	361	205	362
rect	207	361	208	362
rect	210	361	211	362
rect	213	361	214	362
rect	223	361	224	362
rect	226	361	227	362
rect	229	361	230	362
rect	232	361	233	362
rect	235	361	236	362
rect	244	361	245	362
rect	247	361	248	362
rect	256	361	257	362
rect	259	361	260	362
rect	268	361	269	362
rect	274	361	275	362
rect	277	361	278	362
rect	280	361	281	362
rect	289	361	290	362
rect	305	361	306	362
rect	308	361	309	362
rect	311	361	312	362
rect	320	361	321	362
rect	323	361	324	362
rect	326	361	327	362
rect	346	361	347	362
rect	349	361	350	362
rect	358	361	359	362
rect	371	361	372	362
rect	375	361	376	362
rect	392	361	393	362
rect	395	361	396	362
rect	4	362	5	363
rect	7	362	8	363
rect	10	362	11	363
rect	20	362	21	363
rect	51	362	52	363
rect	54	362	55	363
rect	63	362	64	363
rect	72	362	73	363
rect	75	362	76	363
rect	78	362	79	363
rect	81	362	82	363
rect	84	362	85	363
rect	87	362	88	363
rect	91	362	92	363
rect	96	362	97	363
rect	102	362	103	363
rect	105	362	106	363
rect	114	362	115	363
rect	118	362	119	363
rect	123	362	124	363
rect	135	362	136	363
rect	138	362	139	363
rect	147	362	148	363
rect	150	362	151	363
rect	153	362	154	363
rect	157	362	158	363
rect	168	362	169	363
rect	171	362	172	363
rect	174	362	175	363
rect	177	362	178	363
rect	180	362	181	363
rect	186	362	187	363
rect	192	362	193	363
rect	195	362	196	363
rect	204	362	205	363
rect	207	362	208	363
rect	210	362	211	363
rect	213	362	214	363
rect	223	362	224	363
rect	226	362	227	363
rect	229	362	230	363
rect	232	362	233	363
rect	235	362	236	363
rect	244	362	245	363
rect	247	362	248	363
rect	256	362	257	363
rect	259	362	260	363
rect	268	362	269	363
rect	274	362	275	363
rect	277	362	278	363
rect	280	362	281	363
rect	289	362	290	363
rect	305	362	306	363
rect	308	362	309	363
rect	311	362	312	363
rect	320	362	321	363
rect	323	362	324	363
rect	326	362	327	363
rect	346	362	347	363
rect	349	362	350	363
rect	358	362	359	363
rect	371	362	372	363
rect	375	362	376	363
rect	392	362	393	363
rect	395	362	396	363
rect	4	363	5	364
rect	7	363	8	364
rect	10	363	11	364
rect	20	363	21	364
rect	51	363	52	364
rect	54	363	55	364
rect	63	363	64	364
rect	72	363	73	364
rect	75	363	76	364
rect	81	363	82	364
rect	84	363	85	364
rect	87	363	88	364
rect	91	363	92	364
rect	96	363	97	364
rect	102	363	103	364
rect	105	363	106	364
rect	114	363	115	364
rect	118	363	119	364
rect	123	363	124	364
rect	135	363	136	364
rect	138	363	139	364
rect	147	363	148	364
rect	150	363	151	364
rect	153	363	154	364
rect	157	363	158	364
rect	168	363	169	364
rect	171	363	172	364
rect	174	363	175	364
rect	177	363	178	364
rect	180	363	181	364
rect	186	363	187	364
rect	192	363	193	364
rect	195	363	196	364
rect	204	363	205	364
rect	207	363	208	364
rect	210	363	211	364
rect	223	363	224	364
rect	226	363	227	364
rect	229	363	230	364
rect	232	363	233	364
rect	235	363	236	364
rect	244	363	245	364
rect	247	363	248	364
rect	256	363	257	364
rect	259	363	260	364
rect	268	363	269	364
rect	274	363	275	364
rect	277	363	278	364
rect	289	363	290	364
rect	305	363	306	364
rect	308	363	309	364
rect	311	363	312	364
rect	320	363	321	364
rect	326	363	327	364
rect	346	363	347	364
rect	349	363	350	364
rect	358	363	359	364
rect	371	363	372	364
rect	375	363	376	364
rect	392	363	393	364
rect	395	363	396	364
rect	4	364	5	365
rect	7	364	8	365
rect	10	364	11	365
rect	20	364	21	365
rect	51	364	52	365
rect	54	364	55	365
rect	63	364	64	365
rect	72	364	73	365
rect	75	364	76	365
rect	81	364	82	365
rect	84	364	85	365
rect	87	364	88	365
rect	91	364	92	365
rect	96	364	97	365
rect	102	364	103	365
rect	105	364	106	365
rect	114	364	115	365
rect	118	364	119	365
rect	123	364	124	365
rect	135	364	136	365
rect	138	364	139	365
rect	147	364	148	365
rect	150	364	151	365
rect	153	364	154	365
rect	157	364	158	365
rect	168	364	169	365
rect	171	364	172	365
rect	174	364	175	365
rect	177	364	178	365
rect	180	364	181	365
rect	186	364	187	365
rect	192	364	193	365
rect	195	364	196	365
rect	204	364	205	365
rect	207	364	208	365
rect	210	364	211	365
rect	223	364	224	365
rect	226	364	227	365
rect	229	364	230	365
rect	232	364	233	365
rect	235	364	236	365
rect	241	364	242	365
rect	244	364	245	365
rect	247	364	248	365
rect	256	364	257	365
rect	259	364	260	365
rect	268	364	269	365
rect	274	364	275	365
rect	277	364	278	365
rect	289	364	290	365
rect	295	364	296	365
rect	305	364	306	365
rect	308	364	309	365
rect	311	364	312	365
rect	320	364	321	365
rect	326	364	327	365
rect	346	364	347	365
rect	349	364	350	365
rect	358	364	359	365
rect	371	364	372	365
rect	375	364	376	365
rect	392	364	393	365
rect	395	364	396	365
rect	4	365	5	366
rect	7	365	8	366
rect	10	365	11	366
rect	20	365	21	366
rect	51	365	52	366
rect	54	365	55	366
rect	63	365	64	366
rect	75	365	76	366
rect	81	365	82	366
rect	87	365	88	366
rect	91	365	92	366
rect	96	365	97	366
rect	102	365	103	366
rect	105	365	106	366
rect	114	365	115	366
rect	118	365	119	366
rect	123	365	124	366
rect	135	365	136	366
rect	138	365	139	366
rect	147	365	148	366
rect	150	365	151	366
rect	153	365	154	366
rect	157	365	158	366
rect	171	365	172	366
rect	174	365	175	366
rect	177	365	178	366
rect	180	365	181	366
rect	186	365	187	366
rect	192	365	193	366
rect	195	365	196	366
rect	204	365	205	366
rect	207	365	208	366
rect	210	365	211	366
rect	223	365	224	366
rect	226	365	227	366
rect	229	365	230	366
rect	232	365	233	366
rect	235	365	236	366
rect	241	365	242	366
rect	247	365	248	366
rect	256	365	257	366
rect	259	365	260	366
rect	268	365	269	366
rect	274	365	275	366
rect	277	365	278	366
rect	289	365	290	366
rect	295	365	296	366
rect	305	365	306	366
rect	308	365	309	366
rect	320	365	321	366
rect	326	365	327	366
rect	346	365	347	366
rect	349	365	350	366
rect	358	365	359	366
rect	371	365	372	366
rect	375	365	376	366
rect	392	365	393	366
rect	395	365	396	366
rect	4	366	5	367
rect	7	366	8	367
rect	10	366	11	367
rect	20	366	21	367
rect	51	366	52	367
rect	54	366	55	367
rect	63	366	64	367
rect	75	366	76	367
rect	79	366	80	367
rect	81	366	82	367
rect	87	366	88	367
rect	91	366	92	367
rect	94	366	95	367
rect	96	366	97	367
rect	102	366	103	367
rect	105	366	106	367
rect	114	366	115	367
rect	118	366	119	367
rect	123	366	124	367
rect	133	366	134	367
rect	135	366	136	367
rect	138	366	139	367
rect	147	366	148	367
rect	150	366	151	367
rect	153	366	154	367
rect	157	366	158	367
rect	171	366	172	367
rect	174	366	175	367
rect	177	366	178	367
rect	180	366	181	367
rect	186	366	187	367
rect	189	366	190	367
rect	192	366	193	367
rect	195	366	196	367
rect	204	366	205	367
rect	207	366	208	367
rect	210	366	211	367
rect	223	366	224	367
rect	226	366	227	367
rect	229	366	230	367
rect	232	366	233	367
rect	235	366	236	367
rect	241	366	242	367
rect	247	366	248	367
rect	256	366	257	367
rect	259	366	260	367
rect	268	366	269	367
rect	274	366	275	367
rect	277	366	278	367
rect	283	366	284	367
rect	289	366	290	367
rect	295	366	296	367
rect	305	366	306	367
rect	308	366	309	367
rect	320	366	321	367
rect	326	366	327	367
rect	346	366	347	367
rect	349	366	350	367
rect	358	366	359	367
rect	371	366	372	367
rect	375	366	376	367
rect	392	366	393	367
rect	395	366	396	367
rect	4	367	5	368
rect	7	367	8	368
rect	10	367	11	368
rect	20	367	21	368
rect	51	367	52	368
rect	54	367	55	368
rect	63	367	64	368
rect	79	367	80	368
rect	87	367	88	368
rect	91	367	92	368
rect	94	367	95	368
rect	96	367	97	368
rect	102	367	103	368
rect	105	367	106	368
rect	114	367	115	368
rect	118	367	119	368
rect	123	367	124	368
rect	133	367	134	368
rect	135	367	136	368
rect	138	367	139	368
rect	147	367	148	368
rect	150	367	151	368
rect	153	367	154	368
rect	157	367	158	368
rect	171	367	172	368
rect	174	367	175	368
rect	177	367	178	368
rect	180	367	181	368
rect	186	367	187	368
rect	189	367	190	368
rect	192	367	193	368
rect	195	367	196	368
rect	204	367	205	368
rect	207	367	208	368
rect	210	367	211	368
rect	223	367	224	368
rect	226	367	227	368
rect	229	367	230	368
rect	232	367	233	368
rect	235	367	236	368
rect	241	367	242	368
rect	247	367	248	368
rect	256	367	257	368
rect	259	367	260	368
rect	268	367	269	368
rect	274	367	275	368
rect	277	367	278	368
rect	283	367	284	368
rect	289	367	290	368
rect	295	367	296	368
rect	305	367	306	368
rect	308	367	309	368
rect	320	367	321	368
rect	346	367	347	368
rect	349	367	350	368
rect	358	367	359	368
rect	371	367	372	368
rect	375	367	376	368
rect	392	367	393	368
rect	395	367	396	368
rect	4	368	5	369
rect	7	368	8	369
rect	10	368	11	369
rect	20	368	21	369
rect	51	368	52	369
rect	54	368	55	369
rect	63	368	64	369
rect	73	368	74	369
rect	79	368	80	369
rect	87	368	88	369
rect	91	368	92	369
rect	94	368	95	369
rect	96	368	97	369
rect	102	368	103	369
rect	105	368	106	369
rect	114	368	115	369
rect	118	368	119	369
rect	123	368	124	369
rect	133	368	134	369
rect	135	368	136	369
rect	138	368	139	369
rect	147	368	148	369
rect	150	368	151	369
rect	153	368	154	369
rect	157	368	158	369
rect	171	368	172	369
rect	174	368	175	369
rect	177	368	178	369
rect	180	368	181	369
rect	186	368	187	369
rect	189	368	190	369
rect	192	368	193	369
rect	195	368	196	369
rect	204	368	205	369
rect	207	368	208	369
rect	210	368	211	369
rect	223	368	224	369
rect	226	368	227	369
rect	229	368	230	369
rect	232	368	233	369
rect	235	368	236	369
rect	241	368	242	369
rect	247	368	248	369
rect	256	368	257	369
rect	259	368	260	369
rect	268	368	269	369
rect	274	368	275	369
rect	277	368	278	369
rect	283	368	284	369
rect	289	368	290	369
rect	295	368	296	369
rect	305	368	306	369
rect	308	368	309	369
rect	320	368	321	369
rect	346	368	347	369
rect	349	368	350	369
rect	358	368	359	369
rect	371	368	372	369
rect	375	368	376	369
rect	392	368	393	369
rect	395	368	396	369
rect	4	369	5	370
rect	7	369	8	370
rect	10	369	11	370
rect	20	369	21	370
rect	51	369	52	370
rect	54	369	55	370
rect	63	369	64	370
rect	73	369	74	370
rect	79	369	80	370
rect	87	369	88	370
rect	91	369	92	370
rect	94	369	95	370
rect	96	369	97	370
rect	102	369	103	370
rect	114	369	115	370
rect	118	369	119	370
rect	123	369	124	370
rect	133	369	134	370
rect	135	369	136	370
rect	138	369	139	370
rect	147	369	148	370
rect	157	369	158	370
rect	171	369	172	370
rect	174	369	175	370
rect	177	369	178	370
rect	180	369	181	370
rect	186	369	187	370
rect	189	369	190	370
rect	192	369	193	370
rect	204	369	205	370
rect	207	369	208	370
rect	210	369	211	370
rect	223	369	224	370
rect	226	369	227	370
rect	229	369	230	370
rect	232	369	233	370
rect	235	369	236	370
rect	241	369	242	370
rect	247	369	248	370
rect	256	369	257	370
rect	259	369	260	370
rect	268	369	269	370
rect	274	369	275	370
rect	277	369	278	370
rect	283	369	284	370
rect	289	369	290	370
rect	295	369	296	370
rect	305	369	306	370
rect	308	369	309	370
rect	346	369	347	370
rect	358	369	359	370
rect	371	369	372	370
rect	375	369	376	370
rect	392	369	393	370
rect	395	369	396	370
rect	4	370	5	371
rect	7	370	8	371
rect	10	370	11	371
rect	20	370	21	371
rect	51	370	52	371
rect	54	370	55	371
rect	63	370	64	371
rect	73	370	74	371
rect	76	370	77	371
rect	79	370	80	371
rect	87	370	88	371
rect	91	370	92	371
rect	94	370	95	371
rect	96	370	97	371
rect	102	370	103	371
rect	114	370	115	371
rect	118	370	119	371
rect	123	370	124	371
rect	130	370	131	371
rect	133	370	134	371
rect	135	370	136	371
rect	138	370	139	371
rect	147	370	148	371
rect	157	370	158	371
rect	164	370	165	371
rect	167	370	168	371
rect	171	370	172	371
rect	174	370	175	371
rect	177	370	178	371
rect	180	370	181	371
rect	186	370	187	371
rect	189	370	190	371
rect	192	370	193	371
rect	204	370	205	371
rect	207	370	208	371
rect	210	370	211	371
rect	223	370	224	371
rect	226	370	227	371
rect	229	370	230	371
rect	232	370	233	371
rect	235	370	236	371
rect	241	370	242	371
rect	247	370	248	371
rect	256	370	257	371
rect	259	370	260	371
rect	268	370	269	371
rect	274	370	275	371
rect	277	370	278	371
rect	280	370	281	371
rect	283	370	284	371
rect	289	370	290	371
rect	295	370	296	371
rect	305	370	306	371
rect	308	370	309	371
rect	323	370	324	371
rect	346	370	347	371
rect	358	370	359	371
rect	371	370	372	371
rect	375	370	376	371
rect	392	370	393	371
rect	395	370	396	371
rect	4	371	5	372
rect	7	371	8	372
rect	10	371	11	372
rect	20	371	21	372
rect	51	371	52	372
rect	54	371	55	372
rect	63	371	64	372
rect	73	371	74	372
rect	76	371	77	372
rect	79	371	80	372
rect	87	371	88	372
rect	91	371	92	372
rect	94	371	95	372
rect	96	371	97	372
rect	114	371	115	372
rect	118	371	119	372
rect	123	371	124	372
rect	130	371	131	372
rect	133	371	134	372
rect	135	371	136	372
rect	138	371	139	372
rect	157	371	158	372
rect	164	371	165	372
rect	167	371	168	372
rect	174	371	175	372
rect	177	371	178	372
rect	180	371	181	372
rect	189	371	190	372
rect	204	371	205	372
rect	207	371	208	372
rect	223	371	224	372
rect	226	371	227	372
rect	229	371	230	372
rect	235	371	236	372
rect	241	371	242	372
rect	247	371	248	372
rect	256	371	257	372
rect	259	371	260	372
rect	274	371	275	372
rect	277	371	278	372
rect	280	371	281	372
rect	283	371	284	372
rect	289	371	290	372
rect	295	371	296	372
rect	305	371	306	372
rect	308	371	309	372
rect	323	371	324	372
rect	346	371	347	372
rect	371	371	372	372
rect	375	371	376	372
rect	392	371	393	372
rect	395	371	396	372
rect	4	372	5	373
rect	7	372	8	373
rect	10	372	11	373
rect	20	372	21	373
rect	51	372	52	373
rect	54	372	55	373
rect	63	372	64	373
rect	70	372	71	373
rect	73	372	74	373
rect	76	372	77	373
rect	79	372	80	373
rect	87	372	88	373
rect	91	372	92	373
rect	94	372	95	373
rect	96	372	97	373
rect	114	372	115	373
rect	118	372	119	373
rect	123	372	124	373
rect	130	372	131	373
rect	133	372	134	373
rect	135	372	136	373
rect	138	372	139	373
rect	145	372	146	373
rect	151	372	152	373
rect	157	372	158	373
rect	164	372	165	373
rect	167	372	168	373
rect	174	372	175	373
rect	177	372	178	373
rect	180	372	181	373
rect	189	372	190	373
rect	201	372	202	373
rect	204	372	205	373
rect	207	372	208	373
rect	220	372	221	373
rect	223	372	224	373
rect	226	372	227	373
rect	229	372	230	373
rect	235	372	236	373
rect	241	372	242	373
rect	244	372	245	373
rect	247	372	248	373
rect	256	372	257	373
rect	259	372	260	373
rect	271	372	272	373
rect	274	372	275	373
rect	277	372	278	373
rect	280	372	281	373
rect	283	372	284	373
rect	289	372	290	373
rect	295	372	296	373
rect	305	372	306	373
rect	308	372	309	373
rect	323	372	324	373
rect	326	372	327	373
rect	346	372	347	373
rect	348	372	349	373
rect	371	372	372	373
rect	375	372	376	373
rect	392	372	393	373
rect	395	372	396	373
rect	7	373	8	374
rect	10	373	11	374
rect	51	373	52	374
rect	54	373	55	374
rect	63	373	64	374
rect	70	373	71	374
rect	73	373	74	374
rect	76	373	77	374
rect	79	373	80	374
rect	87	373	88	374
rect	91	373	92	374
rect	94	373	95	374
rect	118	373	119	374
rect	123	373	124	374
rect	130	373	131	374
rect	133	373	134	374
rect	138	373	139	374
rect	145	373	146	374
rect	151	373	152	374
rect	157	373	158	374
rect	164	373	165	374
rect	167	373	168	374
rect	174	373	175	374
rect	177	373	178	374
rect	189	373	190	374
rect	201	373	202	374
rect	204	373	205	374
rect	220	373	221	374
rect	223	373	224	374
rect	226	373	227	374
rect	235	373	236	374
rect	241	373	242	374
rect	244	373	245	374
rect	259	373	260	374
rect	271	373	272	374
rect	274	373	275	374
rect	277	373	278	374
rect	280	373	281	374
rect	283	373	284	374
rect	289	373	290	374
rect	295	373	296	374
rect	305	373	306	374
rect	323	373	324	374
rect	326	373	327	374
rect	346	373	347	374
rect	348	373	349	374
rect	371	373	372	374
rect	392	373	393	374
rect	395	373	396	374
rect	7	374	8	375
rect	10	374	11	375
rect	51	374	52	375
rect	54	374	55	375
rect	63	374	64	375
rect	67	374	68	375
rect	70	374	71	375
rect	73	374	74	375
rect	76	374	77	375
rect	79	374	80	375
rect	87	374	88	375
rect	91	374	92	375
rect	94	374	95	375
rect	106	374	107	375
rect	118	374	119	375
rect	121	374	122	375
rect	123	374	124	375
rect	130	374	131	375
rect	133	374	134	375
rect	138	374	139	375
rect	145	374	146	375
rect	148	374	149	375
rect	151	374	152	375
rect	157	374	158	375
rect	164	374	165	375
rect	167	374	168	375
rect	174	374	175	375
rect	177	374	178	375
rect	189	374	190	375
rect	192	374	193	375
rect	201	374	202	375
rect	204	374	205	375
rect	217	374	218	375
rect	220	374	221	375
rect	223	374	224	375
rect	226	374	227	375
rect	232	374	233	375
rect	235	374	236	375
rect	241	374	242	375
rect	244	374	245	375
rect	253	374	254	375
rect	259	374	260	375
rect	268	374	269	375
rect	271	374	272	375
rect	274	374	275	375
rect	277	374	278	375
rect	280	374	281	375
rect	283	374	284	375
rect	289	374	290	375
rect	295	374	296	375
rect	305	374	306	375
rect	323	374	324	375
rect	326	374	327	375
rect	332	374	333	375
rect	346	374	347	375
rect	348	374	349	375
rect	371	374	372	375
rect	392	374	393	375
rect	395	374	396	375
rect	10	375	11	376
rect	51	375	52	376
rect	63	375	64	376
rect	67	375	68	376
rect	70	375	71	376
rect	73	375	74	376
rect	76	375	77	376
rect	79	375	80	376
rect	87	375	88	376
rect	91	375	92	376
rect	94	375	95	376
rect	106	375	107	376
rect	118	375	119	376
rect	121	375	122	376
rect	123	375	124	376
rect	130	375	131	376
rect	133	375	134	376
rect	138	375	139	376
rect	145	375	146	376
rect	148	375	149	376
rect	151	375	152	376
rect	157	375	158	376
rect	164	375	165	376
rect	167	375	168	376
rect	174	375	175	376
rect	177	375	178	376
rect	189	375	190	376
rect	192	375	193	376
rect	201	375	202	376
rect	204	375	205	376
rect	217	375	218	376
rect	220	375	221	376
rect	223	375	224	376
rect	226	375	227	376
rect	232	375	233	376
rect	235	375	236	376
rect	241	375	242	376
rect	244	375	245	376
rect	253	375	254	376
rect	259	375	260	376
rect	268	375	269	376
rect	271	375	272	376
rect	274	375	275	376
rect	277	375	278	376
rect	280	375	281	376
rect	283	375	284	376
rect	289	375	290	376
rect	295	375	296	376
rect	305	375	306	376
rect	323	375	324	376
rect	326	375	327	376
rect	332	375	333	376
rect	346	375	347	376
rect	348	375	349	376
rect	371	375	372	376
rect	392	375	393	376
rect	4	376	5	377
rect	10	376	11	377
rect	51	376	52	377
rect	63	376	64	377
rect	67	376	68	377
rect	70	376	71	377
rect	73	376	74	377
rect	76	376	77	377
rect	79	376	80	377
rect	87	376	88	377
rect	91	376	92	377
rect	94	376	95	377
rect	106	376	107	377
rect	118	376	119	377
rect	121	376	122	377
rect	123	376	124	377
rect	130	376	131	377
rect	133	376	134	377
rect	138	376	139	377
rect	145	376	146	377
rect	148	376	149	377
rect	151	376	152	377
rect	157	376	158	377
rect	164	376	165	377
rect	167	376	168	377
rect	174	376	175	377
rect	177	376	178	377
rect	189	376	190	377
rect	192	376	193	377
rect	201	376	202	377
rect	204	376	205	377
rect	217	376	218	377
rect	220	376	221	377
rect	223	376	224	377
rect	226	376	227	377
rect	232	376	233	377
rect	235	376	236	377
rect	241	376	242	377
rect	244	376	245	377
rect	253	376	254	377
rect	259	376	260	377
rect	268	376	269	377
rect	271	376	272	377
rect	274	376	275	377
rect	277	376	278	377
rect	280	376	281	377
rect	283	376	284	377
rect	289	376	290	377
rect	295	376	296	377
rect	305	376	306	377
rect	323	376	324	377
rect	326	376	327	377
rect	332	376	333	377
rect	346	376	347	377
rect	348	376	349	377
rect	351	376	352	377
rect	364	376	365	377
rect	371	376	372	377
rect	392	376	393	377
rect	4	377	5	378
rect	10	377	11	378
rect	51	377	52	378
rect	63	377	64	378
rect	67	377	68	378
rect	70	377	71	378
rect	73	377	74	378
rect	76	377	77	378
rect	79	377	80	378
rect	87	377	88	378
rect	91	377	92	378
rect	94	377	95	378
rect	106	377	107	378
rect	118	377	119	378
rect	121	377	122	378
rect	123	377	124	378
rect	130	377	131	378
rect	133	377	134	378
rect	145	377	146	378
rect	148	377	149	378
rect	151	377	152	378
rect	157	377	158	378
rect	164	377	165	378
rect	167	377	168	378
rect	174	377	175	378
rect	189	377	190	378
rect	192	377	193	378
rect	201	377	202	378
rect	204	377	205	378
rect	217	377	218	378
rect	220	377	221	378
rect	223	377	224	378
rect	226	377	227	378
rect	232	377	233	378
rect	235	377	236	378
rect	241	377	242	378
rect	244	377	245	378
rect	253	377	254	378
rect	268	377	269	378
rect	271	377	272	378
rect	274	377	275	378
rect	277	377	278	378
rect	280	377	281	378
rect	283	377	284	378
rect	289	377	290	378
rect	295	377	296	378
rect	323	377	324	378
rect	326	377	327	378
rect	332	377	333	378
rect	346	377	347	378
rect	348	377	349	378
rect	351	377	352	378
rect	364	377	365	378
rect	392	377	393	378
rect	4	378	5	379
rect	8	378	9	379
rect	10	378	11	379
rect	51	378	52	379
rect	63	378	64	379
rect	67	378	68	379
rect	70	378	71	379
rect	73	378	74	379
rect	76	378	77	379
rect	79	378	80	379
rect	87	378	88	379
rect	91	378	92	379
rect	94	378	95	379
rect	106	378	107	379
rect	118	378	119	379
rect	121	378	122	379
rect	123	378	124	379
rect	130	378	131	379
rect	133	378	134	379
rect	142	378	143	379
rect	145	378	146	379
rect	148	378	149	379
rect	151	378	152	379
rect	157	378	158	379
rect	164	378	165	379
rect	167	378	168	379
rect	174	378	175	379
rect	186	378	187	379
rect	189	378	190	379
rect	192	378	193	379
rect	201	378	202	379
rect	204	378	205	379
rect	217	378	218	379
rect	220	378	221	379
rect	223	378	224	379
rect	226	378	227	379
rect	232	378	233	379
rect	235	378	236	379
rect	241	378	242	379
rect	244	378	245	379
rect	253	378	254	379
rect	265	378	266	379
rect	268	378	269	379
rect	271	378	272	379
rect	274	378	275	379
rect	277	378	278	379
rect	280	378	281	379
rect	283	378	284	379
rect	289	378	290	379
rect	295	378	296	379
rect	311	378	312	379
rect	317	378	318	379
rect	320	378	321	379
rect	323	378	324	379
rect	326	378	327	379
rect	332	378	333	379
rect	346	378	347	379
rect	348	378	349	379
rect	351	378	352	379
rect	364	378	365	379
rect	392	378	393	379
rect	4	379	5	380
rect	8	379	9	380
rect	67	379	68	380
rect	70	379	71	380
rect	73	379	74	380
rect	76	379	77	380
rect	79	379	80	380
rect	91	379	92	380
rect	94	379	95	380
rect	106	379	107	380
rect	118	379	119	380
rect	121	379	122	380
rect	130	379	131	380
rect	133	379	134	380
rect	142	379	143	380
rect	145	379	146	380
rect	148	379	149	380
rect	151	379	152	380
rect	157	379	158	380
rect	164	379	165	380
rect	167	379	168	380
rect	186	379	187	380
rect	189	379	190	380
rect	192	379	193	380
rect	201	379	202	380
rect	217	379	218	380
rect	220	379	221	380
rect	232	379	233	380
rect	241	379	242	380
rect	244	379	245	380
rect	253	379	254	380
rect	265	379	266	380
rect	268	379	269	380
rect	271	379	272	380
rect	274	379	275	380
rect	280	379	281	380
rect	283	379	284	380
rect	295	379	296	380
rect	311	379	312	380
rect	317	379	318	380
rect	320	379	321	380
rect	323	379	324	380
rect	326	379	327	380
rect	332	379	333	380
rect	348	379	349	380
rect	351	379	352	380
rect	364	379	365	380
rect	4	380	5	381
rect	8	380	9	381
rect	14	380	15	381
rect	58	380	59	381
rect	67	380	68	381
rect	70	380	71	381
rect	73	380	74	381
rect	76	380	77	381
rect	79	380	80	381
rect	82	380	83	381
rect	91	380	92	381
rect	94	380	95	381
rect	97	380	98	381
rect	106	380	107	381
rect	115	380	116	381
rect	118	380	119	381
rect	121	380	122	381
rect	130	380	131	381
rect	133	380	134	381
rect	139	380	140	381
rect	142	380	143	381
rect	145	380	146	381
rect	148	380	149	381
rect	151	380	152	381
rect	157	380	158	381
rect	164	380	165	381
rect	167	380	168	381
rect	183	380	184	381
rect	186	380	187	381
rect	189	380	190	381
rect	192	380	193	381
rect	201	380	202	381
rect	217	380	218	381
rect	220	380	221	381
rect	229	380	230	381
rect	232	380	233	381
rect	241	380	242	381
rect	244	380	245	381
rect	253	380	254	381
rect	256	380	257	381
rect	265	380	266	381
rect	268	380	269	381
rect	271	380	272	381
rect	274	380	275	381
rect	280	380	281	381
rect	283	380	284	381
rect	286	380	287	381
rect	295	380	296	381
rect	298	380	299	381
rect	311	380	312	381
rect	317	380	318	381
rect	320	380	321	381
rect	323	380	324	381
rect	326	380	327	381
rect	332	380	333	381
rect	348	380	349	381
rect	351	380	352	381
rect	361	380	362	381
rect	364	380	365	381
rect	4	387	5	388
rect	8	387	9	388
rect	14	387	15	388
rect	20	387	21	388
rect	58	387	59	388
rect	67	387	68	388
rect	70	387	71	388
rect	73	387	74	388
rect	76	387	77	388
rect	79	387	80	388
rect	82	387	83	388
rect	91	387	92	388
rect	94	387	95	388
rect	97	387	98	388
rect	106	387	107	388
rect	115	387	116	388
rect	118	387	119	388
rect	121	387	122	388
rect	124	387	125	388
rect	127	387	128	388
rect	130	387	131	388
rect	139	387	140	388
rect	142	387	143	388
rect	145	387	146	388
rect	148	387	149	388
rect	151	387	152	388
rect	167	387	168	388
rect	173	387	174	388
rect	180	387	181	388
rect	183	387	184	388
rect	192	387	193	388
rect	201	387	202	388
rect	217	387	218	388
rect	220	387	221	388
rect	229	387	230	388
rect	232	387	233	388
rect	241	387	242	388
rect	244	387	245	388
rect	253	387	254	388
rect	256	387	257	388
rect	265	387	266	388
rect	268	387	269	388
rect	271	387	272	388
rect	277	387	278	388
rect	280	387	281	388
rect	283	387	284	388
rect	286	387	287	388
rect	289	387	290	388
rect	295	387	296	388
rect	311	387	312	388
rect	320	387	321	388
rect	323	387	324	388
rect	332	387	333	388
rect	338	387	339	388
rect	345	387	346	388
rect	348	387	349	388
rect	354	387	355	388
rect	364	387	365	388
rect	4	388	5	389
rect	8	388	9	389
rect	14	388	15	389
rect	20	388	21	389
rect	58	388	59	389
rect	67	388	68	389
rect	70	388	71	389
rect	73	388	74	389
rect	76	388	77	389
rect	79	388	80	389
rect	82	388	83	389
rect	91	388	92	389
rect	94	388	95	389
rect	97	388	98	389
rect	106	388	107	389
rect	115	388	116	389
rect	118	388	119	389
rect	121	388	122	389
rect	124	388	125	389
rect	127	388	128	389
rect	130	388	131	389
rect	139	388	140	389
rect	142	388	143	389
rect	145	388	146	389
rect	148	388	149	389
rect	151	388	152	389
rect	167	388	168	389
rect	173	388	174	389
rect	180	388	181	389
rect	183	388	184	389
rect	192	388	193	389
rect	201	388	202	389
rect	217	388	218	389
rect	220	388	221	389
rect	229	388	230	389
rect	232	388	233	389
rect	241	388	242	389
rect	244	388	245	389
rect	253	388	254	389
rect	256	388	257	389
rect	265	388	266	389
rect	268	388	269	389
rect	271	388	272	389
rect	280	388	281	389
rect	283	388	284	389
rect	289	388	290	389
rect	295	388	296	389
rect	311	388	312	389
rect	320	388	321	389
rect	323	388	324	389
rect	332	388	333	389
rect	338	388	339	389
rect	345	388	346	389
rect	348	388	349	389
rect	354	388	355	389
rect	364	388	365	389
rect	4	389	5	390
rect	8	389	9	390
rect	14	389	15	390
rect	20	389	21	390
rect	58	389	59	390
rect	67	389	68	390
rect	70	389	71	390
rect	73	389	74	390
rect	76	389	77	390
rect	79	389	80	390
rect	82	389	83	390
rect	91	389	92	390
rect	94	389	95	390
rect	97	389	98	390
rect	106	389	107	390
rect	115	389	116	390
rect	118	389	119	390
rect	121	389	122	390
rect	124	389	125	390
rect	127	389	128	390
rect	130	389	131	390
rect	139	389	140	390
rect	142	389	143	390
rect	145	389	146	390
rect	148	389	149	390
rect	151	389	152	390
rect	167	389	168	390
rect	173	389	174	390
rect	180	389	181	390
rect	183	389	184	390
rect	192	389	193	390
rect	201	389	202	390
rect	217	389	218	390
rect	220	389	221	390
rect	229	389	230	390
rect	232	389	233	390
rect	241	389	242	390
rect	244	389	245	390
rect	253	389	254	390
rect	256	389	257	390
rect	265	389	266	390
rect	268	389	269	390
rect	271	389	272	390
rect	280	389	281	390
rect	283	389	284	390
rect	289	389	290	390
rect	295	389	296	390
rect	311	389	312	390
rect	320	389	321	390
rect	323	389	324	390
rect	332	389	333	390
rect	338	389	339	390
rect	345	389	346	390
rect	348	389	349	390
rect	354	389	355	390
rect	364	389	365	390
rect	4	390	5	391
rect	8	390	9	391
rect	14	390	15	391
rect	20	390	21	391
rect	58	390	59	391
rect	67	390	68	391
rect	70	390	71	391
rect	73	390	74	391
rect	76	390	77	391
rect	79	390	80	391
rect	82	390	83	391
rect	91	390	92	391
rect	94	390	95	391
rect	97	390	98	391
rect	106	390	107	391
rect	115	390	116	391
rect	118	390	119	391
rect	121	390	122	391
rect	124	390	125	391
rect	127	390	128	391
rect	130	390	131	391
rect	139	390	140	391
rect	142	390	143	391
rect	145	390	146	391
rect	148	390	149	391
rect	151	390	152	391
rect	167	390	168	391
rect	173	390	174	391
rect	180	390	181	391
rect	183	390	184	391
rect	192	390	193	391
rect	201	390	202	391
rect	217	390	218	391
rect	220	390	221	391
rect	229	390	230	391
rect	232	390	233	391
rect	241	390	242	391
rect	244	390	245	391
rect	253	390	254	391
rect	256	390	257	391
rect	265	390	266	391
rect	268	390	269	391
rect	271	390	272	391
rect	280	390	281	391
rect	289	390	290	391
rect	295	390	296	391
rect	311	390	312	391
rect	320	390	321	391
rect	332	390	333	391
rect	338	390	339	391
rect	345	390	346	391
rect	348	390	349	391
rect	354	390	355	391
rect	364	390	365	391
rect	4	391	5	392
rect	8	391	9	392
rect	14	391	15	392
rect	20	391	21	392
rect	58	391	59	392
rect	67	391	68	392
rect	70	391	71	392
rect	73	391	74	392
rect	76	391	77	392
rect	79	391	80	392
rect	82	391	83	392
rect	91	391	92	392
rect	94	391	95	392
rect	97	391	98	392
rect	106	391	107	392
rect	115	391	116	392
rect	118	391	119	392
rect	121	391	122	392
rect	124	391	125	392
rect	127	391	128	392
rect	130	391	131	392
rect	139	391	140	392
rect	142	391	143	392
rect	145	391	146	392
rect	148	391	149	392
rect	151	391	152	392
rect	167	391	168	392
rect	173	391	174	392
rect	180	391	181	392
rect	183	391	184	392
rect	192	391	193	392
rect	201	391	202	392
rect	217	391	218	392
rect	220	391	221	392
rect	229	391	230	392
rect	232	391	233	392
rect	241	391	242	392
rect	244	391	245	392
rect	253	391	254	392
rect	256	391	257	392
rect	263	391	264	392
rect	265	391	266	392
rect	268	391	269	392
rect	271	391	272	392
rect	280	391	281	392
rect	287	391	288	392
rect	289	391	290	392
rect	295	391	296	392
rect	311	391	312	392
rect	320	391	321	392
rect	332	391	333	392
rect	338	391	339	392
rect	345	391	346	392
rect	348	391	349	392
rect	354	391	355	392
rect	364	391	365	392
rect	4	392	5	393
rect	8	392	9	393
rect	14	392	15	393
rect	20	392	21	393
rect	58	392	59	393
rect	67	392	68	393
rect	70	392	71	393
rect	73	392	74	393
rect	76	392	77	393
rect	79	392	80	393
rect	82	392	83	393
rect	91	392	92	393
rect	94	392	95	393
rect	97	392	98	393
rect	106	392	107	393
rect	115	392	116	393
rect	118	392	119	393
rect	124	392	125	393
rect	130	392	131	393
rect	139	392	140	393
rect	142	392	143	393
rect	145	392	146	393
rect	148	392	149	393
rect	151	392	152	393
rect	167	392	168	393
rect	173	392	174	393
rect	180	392	181	393
rect	183	392	184	393
rect	192	392	193	393
rect	201	392	202	393
rect	217	392	218	393
rect	220	392	221	393
rect	229	392	230	393
rect	232	392	233	393
rect	244	392	245	393
rect	253	392	254	393
rect	256	392	257	393
rect	263	392	264	393
rect	265	392	266	393
rect	268	392	269	393
rect	271	392	272	393
rect	280	392	281	393
rect	287	392	288	393
rect	289	392	290	393
rect	295	392	296	393
rect	320	392	321	393
rect	332	392	333	393
rect	338	392	339	393
rect	345	392	346	393
rect	348	392	349	393
rect	354	392	355	393
rect	364	392	365	393
rect	4	393	5	394
rect	8	393	9	394
rect	14	393	15	394
rect	20	393	21	394
rect	58	393	59	394
rect	67	393	68	394
rect	70	393	71	394
rect	73	393	74	394
rect	76	393	77	394
rect	79	393	80	394
rect	82	393	83	394
rect	91	393	92	394
rect	94	393	95	394
rect	97	393	98	394
rect	106	393	107	394
rect	115	393	116	394
rect	118	393	119	394
rect	124	393	125	394
rect	130	393	131	394
rect	139	393	140	394
rect	142	393	143	394
rect	145	393	146	394
rect	148	393	149	394
rect	151	393	152	394
rect	167	393	168	394
rect	173	393	174	394
rect	180	393	181	394
rect	183	393	184	394
rect	192	393	193	394
rect	201	393	202	394
rect	212	393	213	394
rect	217	393	218	394
rect	220	393	221	394
rect	229	393	230	394
rect	232	393	233	394
rect	244	393	245	394
rect	253	393	254	394
rect	256	393	257	394
rect	260	393	261	394
rect	263	393	264	394
rect	265	393	266	394
rect	268	393	269	394
rect	271	393	272	394
rect	280	393	281	394
rect	287	393	288	394
rect	289	393	290	394
rect	295	393	296	394
rect	320	393	321	394
rect	332	393	333	394
rect	338	393	339	394
rect	345	393	346	394
rect	348	393	349	394
rect	354	393	355	394
rect	364	393	365	394
rect	4	394	5	395
rect	8	394	9	395
rect	14	394	15	395
rect	20	394	21	395
rect	58	394	59	395
rect	67	394	68	395
rect	70	394	71	395
rect	73	394	74	395
rect	76	394	77	395
rect	79	394	80	395
rect	82	394	83	395
rect	91	394	92	395
rect	94	394	95	395
rect	97	394	98	395
rect	106	394	107	395
rect	115	394	116	395
rect	118	394	119	395
rect	124	394	125	395
rect	130	394	131	395
rect	142	394	143	395
rect	145	394	146	395
rect	148	394	149	395
rect	151	394	152	395
rect	167	394	168	395
rect	173	394	174	395
rect	180	394	181	395
rect	183	394	184	395
rect	192	394	193	395
rect	201	394	202	395
rect	212	394	213	395
rect	217	394	218	395
rect	220	394	221	395
rect	229	394	230	395
rect	232	394	233	395
rect	244	394	245	395
rect	253	394	254	395
rect	256	394	257	395
rect	260	394	261	395
rect	263	394	264	395
rect	265	394	266	395
rect	268	394	269	395
rect	280	394	281	395
rect	287	394	288	395
rect	289	394	290	395
rect	295	394	296	395
rect	320	394	321	395
rect	338	394	339	395
rect	345	394	346	395
rect	348	394	349	395
rect	354	394	355	395
rect	364	394	365	395
rect	4	395	5	396
rect	8	395	9	396
rect	14	395	15	396
rect	20	395	21	396
rect	58	395	59	396
rect	67	395	68	396
rect	70	395	71	396
rect	73	395	74	396
rect	76	395	77	396
rect	79	395	80	396
rect	82	395	83	396
rect	91	395	92	396
rect	94	395	95	396
rect	97	395	98	396
rect	106	395	107	396
rect	115	395	116	396
rect	118	395	119	396
rect	121	395	122	396
rect	124	395	125	396
rect	130	395	131	396
rect	142	395	143	396
rect	145	395	146	396
rect	148	395	149	396
rect	151	395	152	396
rect	167	395	168	396
rect	173	395	174	396
rect	180	395	181	396
rect	183	395	184	396
rect	192	395	193	396
rect	201	395	202	396
rect	212	395	213	396
rect	217	395	218	396
rect	220	395	221	396
rect	229	395	230	396
rect	232	395	233	396
rect	242	395	243	396
rect	244	395	245	396
rect	253	395	254	396
rect	256	395	257	396
rect	260	395	261	396
rect	263	395	264	396
rect	265	395	266	396
rect	268	395	269	396
rect	280	395	281	396
rect	284	395	285	396
rect	287	395	288	396
rect	289	395	290	396
rect	295	395	296	396
rect	320	395	321	396
rect	338	395	339	396
rect	345	395	346	396
rect	348	395	349	396
rect	354	395	355	396
rect	364	395	365	396
rect	4	396	5	397
rect	8	396	9	397
rect	14	396	15	397
rect	20	396	21	397
rect	58	396	59	397
rect	67	396	68	397
rect	70	396	71	397
rect	73	396	74	397
rect	76	396	77	397
rect	79	396	80	397
rect	82	396	83	397
rect	91	396	92	397
rect	94	396	95	397
rect	97	396	98	397
rect	106	396	107	397
rect	115	396	116	397
rect	118	396	119	397
rect	121	396	122	397
rect	124	396	125	397
rect	142	396	143	397
rect	145	396	146	397
rect	148	396	149	397
rect	151	396	152	397
rect	167	396	168	397
rect	173	396	174	397
rect	180	396	181	397
rect	183	396	184	397
rect	192	396	193	397
rect	201	396	202	397
rect	212	396	213	397
rect	217	396	218	397
rect	220	396	221	397
rect	229	396	230	397
rect	232	396	233	397
rect	242	396	243	397
rect	244	396	245	397
rect	253	396	254	397
rect	256	396	257	397
rect	260	396	261	397
rect	263	396	264	397
rect	268	396	269	397
rect	284	396	285	397
rect	287	396	288	397
rect	295	396	296	397
rect	320	396	321	397
rect	338	396	339	397
rect	345	396	346	397
rect	348	396	349	397
rect	364	396	365	397
rect	4	397	5	398
rect	8	397	9	398
rect	14	397	15	398
rect	20	397	21	398
rect	58	397	59	398
rect	67	397	68	398
rect	70	397	71	398
rect	73	397	74	398
rect	76	397	77	398
rect	79	397	80	398
rect	82	397	83	398
rect	91	397	92	398
rect	94	397	95	398
rect	97	397	98	398
rect	106	397	107	398
rect	112	397	113	398
rect	115	397	116	398
rect	118	397	119	398
rect	121	397	122	398
rect	124	397	125	398
rect	140	397	141	398
rect	142	397	143	398
rect	145	397	146	398
rect	148	397	149	398
rect	151	397	152	398
rect	167	397	168	398
rect	173	397	174	398
rect	180	397	181	398
rect	183	397	184	398
rect	192	397	193	398
rect	201	397	202	398
rect	212	397	213	398
rect	215	397	216	398
rect	217	397	218	398
rect	220	397	221	398
rect	227	397	228	398
rect	229	397	230	398
rect	232	397	233	398
rect	242	397	243	398
rect	244	397	245	398
rect	253	397	254	398
rect	256	397	257	398
rect	260	397	261	398
rect	263	397	264	398
rect	268	397	269	398
rect	284	397	285	398
rect	287	397	288	398
rect	293	397	294	398
rect	295	397	296	398
rect	320	397	321	398
rect	338	397	339	398
rect	345	397	346	398
rect	348	397	349	398
rect	364	397	365	398
rect	4	398	5	399
rect	8	398	9	399
rect	14	398	15	399
rect	20	398	21	399
rect	58	398	59	399
rect	67	398	68	399
rect	70	398	71	399
rect	73	398	74	399
rect	76	398	77	399
rect	79	398	80	399
rect	82	398	83	399
rect	91	398	92	399
rect	94	398	95	399
rect	97	398	98	399
rect	106	398	107	399
rect	112	398	113	399
rect	115	398	116	399
rect	118	398	119	399
rect	121	398	122	399
rect	124	398	125	399
rect	140	398	141	399
rect	142	398	143	399
rect	145	398	146	399
rect	151	398	152	399
rect	167	398	168	399
rect	173	398	174	399
rect	180	398	181	399
rect	183	398	184	399
rect	192	398	193	399
rect	212	398	213	399
rect	215	398	216	399
rect	217	398	218	399
rect	220	398	221	399
rect	227	398	228	399
rect	232	398	233	399
rect	242	398	243	399
rect	244	398	245	399
rect	260	398	261	399
rect	263	398	264	399
rect	268	398	269	399
rect	284	398	285	399
rect	287	398	288	399
rect	293	398	294	399
rect	295	398	296	399
rect	338	398	339	399
rect	345	398	346	399
rect	348	398	349	399
rect	4	399	5	400
rect	8	399	9	400
rect	14	399	15	400
rect	20	399	21	400
rect	58	399	59	400
rect	67	399	68	400
rect	70	399	71	400
rect	73	399	74	400
rect	76	399	77	400
rect	79	399	80	400
rect	82	399	83	400
rect	91	399	92	400
rect	94	399	95	400
rect	97	399	98	400
rect	106	399	107	400
rect	112	399	113	400
rect	115	399	116	400
rect	118	399	119	400
rect	121	399	122	400
rect	124	399	125	400
rect	130	399	131	400
rect	140	399	141	400
rect	142	399	143	400
rect	145	399	146	400
rect	151	399	152	400
rect	167	399	168	400
rect	173	399	174	400
rect	180	399	181	400
rect	183	399	184	400
rect	192	399	193	400
rect	206	399	207	400
rect	209	399	210	400
rect	212	399	213	400
rect	215	399	216	400
rect	217	399	218	400
rect	220	399	221	400
rect	227	399	228	400
rect	232	399	233	400
rect	239	399	240	400
rect	242	399	243	400
rect	244	399	245	400
rect	260	399	261	400
rect	263	399	264	400
rect	266	399	267	400
rect	268	399	269	400
rect	275	399	276	400
rect	284	399	285	400
rect	287	399	288	400
rect	293	399	294	400
rect	295	399	296	400
rect	331	399	332	400
rect	338	399	339	400
rect	345	399	346	400
rect	348	399	349	400
rect	4	400	5	401
rect	8	400	9	401
rect	14	400	15	401
rect	20	400	21	401
rect	58	400	59	401
rect	67	400	68	401
rect	73	400	74	401
rect	76	400	77	401
rect	79	400	80	401
rect	91	400	92	401
rect	94	400	95	401
rect	106	400	107	401
rect	112	400	113	401
rect	115	400	116	401
rect	118	400	119	401
rect	121	400	122	401
rect	124	400	125	401
rect	130	400	131	401
rect	140	400	141	401
rect	142	400	143	401
rect	145	400	146	401
rect	151	400	152	401
rect	167	400	168	401
rect	173	400	174	401
rect	180	400	181	401
rect	183	400	184	401
rect	192	400	193	401
rect	206	400	207	401
rect	209	400	210	401
rect	212	400	213	401
rect	215	400	216	401
rect	217	400	218	401
rect	220	400	221	401
rect	227	400	228	401
rect	232	400	233	401
rect	239	400	240	401
rect	242	400	243	401
rect	244	400	245	401
rect	260	400	261	401
rect	263	400	264	401
rect	266	400	267	401
rect	268	400	269	401
rect	275	400	276	401
rect	284	400	285	401
rect	287	400	288	401
rect	293	400	294	401
rect	295	400	296	401
rect	331	400	332	401
rect	338	400	339	401
rect	345	400	346	401
rect	4	401	5	402
rect	8	401	9	402
rect	14	401	15	402
rect	20	401	21	402
rect	58	401	59	402
rect	63	401	64	402
rect	67	401	68	402
rect	73	401	74	402
rect	76	401	77	402
rect	79	401	80	402
rect	81	401	82	402
rect	91	401	92	402
rect	94	401	95	402
rect	106	401	107	402
rect	112	401	113	402
rect	115	401	116	402
rect	118	401	119	402
rect	121	401	122	402
rect	124	401	125	402
rect	130	401	131	402
rect	140	401	141	402
rect	142	401	143	402
rect	145	401	146	402
rect	151	401	152	402
rect	167	401	168	402
rect	173	401	174	402
rect	180	401	181	402
rect	183	401	184	402
rect	192	401	193	402
rect	206	401	207	402
rect	209	401	210	402
rect	212	401	213	402
rect	215	401	216	402
rect	217	401	218	402
rect	220	401	221	402
rect	227	401	228	402
rect	232	401	233	402
rect	239	401	240	402
rect	242	401	243	402
rect	244	401	245	402
rect	260	401	261	402
rect	263	401	264	402
rect	266	401	267	402
rect	268	401	269	402
rect	275	401	276	402
rect	284	401	285	402
rect	287	401	288	402
rect	293	401	294	402
rect	295	401	296	402
rect	306	401	307	402
rect	312	401	313	402
rect	318	401	319	402
rect	328	401	329	402
rect	331	401	332	402
rect	338	401	339	402
rect	345	401	346	402
rect	4	402	5	403
rect	8	402	9	403
rect	14	402	15	403
rect	20	402	21	403
rect	58	402	59	403
rect	63	402	64	403
rect	73	402	74	403
rect	79	402	80	403
rect	81	402	82	403
rect	91	402	92	403
rect	94	402	95	403
rect	112	402	113	403
rect	115	402	116	403
rect	121	402	122	403
rect	130	402	131	403
rect	140	402	141	403
rect	142	402	143	403
rect	151	402	152	403
rect	167	402	168	403
rect	173	402	174	403
rect	180	402	181	403
rect	183	402	184	403
rect	192	402	193	403
rect	206	402	207	403
rect	209	402	210	403
rect	212	402	213	403
rect	215	402	216	403
rect	227	402	228	403
rect	239	402	240	403
rect	242	402	243	403
rect	244	402	245	403
rect	260	402	261	403
rect	263	402	264	403
rect	266	402	267	403
rect	275	402	276	403
rect	284	402	285	403
rect	287	402	288	403
rect	293	402	294	403
rect	295	402	296	403
rect	306	402	307	403
rect	312	402	313	403
rect	318	402	319	403
rect	328	402	329	403
rect	331	402	332	403
rect	345	402	346	403
rect	4	403	5	404
rect	8	403	9	404
rect	14	403	15	404
rect	20	403	21	404
rect	58	403	59	404
rect	60	403	61	404
rect	63	403	64	404
rect	73	403	74	404
rect	79	403	80	404
rect	81	403	82	404
rect	84	403	85	404
rect	91	403	92	404
rect	94	403	95	404
rect	97	403	98	404
rect	112	403	113	404
rect	115	403	116	404
rect	121	403	122	404
rect	127	403	128	404
rect	130	403	131	404
rect	140	403	141	404
rect	142	403	143	404
rect	151	403	152	404
rect	167	403	168	404
rect	173	403	174	404
rect	180	403	181	404
rect	183	403	184	404
rect	192	403	193	404
rect	197	403	198	404
rect	206	403	207	404
rect	209	403	210	404
rect	212	403	213	404
rect	215	403	216	404
rect	221	403	222	404
rect	227	403	228	404
rect	230	403	231	404
rect	236	403	237	404
rect	239	403	240	404
rect	242	403	243	404
rect	244	403	245	404
rect	260	403	261	404
rect	263	403	264	404
rect	266	403	267	404
rect	272	403	273	404
rect	275	403	276	404
rect	284	403	285	404
rect	287	403	288	404
rect	293	403	294	404
rect	295	403	296	404
rect	306	403	307	404
rect	312	403	313	404
rect	318	403	319	404
rect	328	403	329	404
rect	331	403	332	404
rect	345	403	346	404
rect	60	404	61	405
rect	63	404	64	405
rect	81	404	82	405
rect	84	404	85	405
rect	91	404	92	405
rect	97	404	98	405
rect	112	404	113	405
rect	121	404	122	405
rect	127	404	128	405
rect	130	404	131	405
rect	140	404	141	405
rect	197	404	198	405
rect	206	404	207	405
rect	209	404	210	405
rect	212	404	213	405
rect	215	404	216	405
rect	221	404	222	405
rect	227	404	228	405
rect	230	404	231	405
rect	236	404	237	405
rect	239	404	240	405
rect	242	404	243	405
rect	260	404	261	405
rect	263	404	264	405
rect	266	404	267	405
rect	272	404	273	405
rect	275	404	276	405
rect	284	404	285	405
rect	287	404	288	405
rect	293	404	294	405
rect	306	404	307	405
rect	312	404	313	405
rect	318	404	319	405
rect	328	404	329	405
rect	331	404	332	405
rect	60	405	61	406
rect	63	405	64	406
rect	66	405	67	406
rect	75	405	76	406
rect	78	405	79	406
rect	81	405	82	406
rect	84	405	85	406
rect	91	405	92	406
rect	97	405	98	406
rect	100	405	101	406
rect	109	405	110	406
rect	112	405	113	406
rect	121	405	122	406
rect	124	405	125	406
rect	127	405	128	406
rect	130	405	131	406
rect	140	405	141	406
rect	146	405	147	406
rect	197	405	198	406
rect	200	405	201	406
rect	206	405	207	406
rect	209	405	210	406
rect	212	405	213	406
rect	215	405	216	406
rect	218	405	219	406
rect	221	405	222	406
rect	227	405	228	406
rect	230	405	231	406
rect	236	405	237	406
rect	239	405	240	406
rect	242	405	243	406
rect	251	405	252	406
rect	260	405	261	406
rect	263	405	264	406
rect	266	405	267	406
rect	272	405	273	406
rect	275	405	276	406
rect	284	405	285	406
rect	287	405	288	406
rect	293	405	294	406
rect	303	405	304	406
rect	306	405	307	406
rect	312	405	313	406
rect	318	405	319	406
rect	328	405	329	406
rect	331	405	332	406
rect	57	412	58	413
rect	63	412	64	413
rect	66	412	67	413
rect	72	412	73	413
rect	75	412	76	413
rect	78	412	79	413
rect	81	412	82	413
rect	97	412	98	413
rect	100	412	101	413
rect	103	412	104	413
rect	109	412	110	413
rect	112	412	113	413
rect	118	412	119	413
rect	121	412	122	413
rect	124	412	125	413
rect	127	412	128	413
rect	130	412	131	413
rect	133	412	134	413
rect	143	412	144	413
rect	146	412	147	413
rect	197	412	198	413
rect	200	412	201	413
rect	206	412	207	413
rect	209	412	210	413
rect	212	412	213	413
rect	218	412	219	413
rect	221	412	222	413
rect	230	412	231	413
rect	239	412	240	413
rect	242	412	243	413
rect	251	412	252	413
rect	257	412	258	413
rect	260	412	261	413
rect	263	412	264	413
rect	266	412	267	413
rect	275	412	276	413
rect	278	412	279	413
rect	284	412	285	413
rect	287	412	288	413
rect	293	412	294	413
rect	297	412	298	413
rect	303	412	304	413
rect	306	412	307	413
rect	312	412	313	413
rect	325	412	326	413
rect	328	412	329	413
rect	331	412	332	413
rect	57	413	58	414
rect	63	413	64	414
rect	66	413	67	414
rect	75	413	76	414
rect	81	413	82	414
rect	97	413	98	414
rect	100	413	101	414
rect	103	413	104	414
rect	109	413	110	414
rect	118	413	119	414
rect	121	413	122	414
rect	124	413	125	414
rect	127	413	128	414
rect	130	413	131	414
rect	133	413	134	414
rect	143	413	144	414
rect	146	413	147	414
rect	197	413	198	414
rect	200	413	201	414
rect	206	413	207	414
rect	209	413	210	414
rect	212	413	213	414
rect	218	413	219	414
rect	221	413	222	414
rect	230	413	231	414
rect	239	413	240	414
rect	242	413	243	414
rect	251	413	252	414
rect	257	413	258	414
rect	260	413	261	414
rect	266	413	267	414
rect	275	413	276	414
rect	278	413	279	414
rect	284	413	285	414
rect	287	413	288	414
rect	293	413	294	414
rect	297	413	298	414
rect	303	413	304	414
rect	306	413	307	414
rect	325	413	326	414
rect	328	413	329	414
rect	331	413	332	414
rect	57	414	58	415
rect	63	414	64	415
rect	66	414	67	415
rect	75	414	76	415
rect	81	414	82	415
rect	89	414	90	415
rect	97	414	98	415
rect	100	414	101	415
rect	103	414	104	415
rect	109	414	110	415
rect	118	414	119	415
rect	121	414	122	415
rect	124	414	125	415
rect	127	414	128	415
rect	130	414	131	415
rect	133	414	134	415
rect	143	414	144	415
rect	146	414	147	415
rect	197	414	198	415
rect	200	414	201	415
rect	206	414	207	415
rect	209	414	210	415
rect	212	414	213	415
rect	218	414	219	415
rect	221	414	222	415
rect	230	414	231	415
rect	237	414	238	415
rect	239	414	240	415
rect	242	414	243	415
rect	251	414	252	415
rect	257	414	258	415
rect	260	414	261	415
rect	266	414	267	415
rect	268	414	269	415
rect	275	414	276	415
rect	278	414	279	415
rect	284	414	285	415
rect	287	414	288	415
rect	293	414	294	415
rect	297	414	298	415
rect	303	414	304	415
rect	306	414	307	415
rect	325	414	326	415
rect	328	414	329	415
rect	331	414	332	415
rect	57	415	58	416
rect	63	415	64	416
rect	66	415	67	416
rect	81	415	82	416
rect	89	415	90	416
rect	97	415	98	416
rect	100	415	101	416
rect	103	415	104	416
rect	124	415	125	416
rect	127	415	128	416
rect	130	415	131	416
rect	133	415	134	416
rect	146	415	147	416
rect	197	415	198	416
rect	200	415	201	416
rect	206	415	207	416
rect	209	415	210	416
rect	212	415	213	416
rect	218	415	219	416
rect	221	415	222	416
rect	237	415	238	416
rect	239	415	240	416
rect	242	415	243	416
rect	251	415	252	416
rect	257	415	258	416
rect	260	415	261	416
rect	266	415	267	416
rect	268	415	269	416
rect	275	415	276	416
rect	278	415	279	416
rect	284	415	285	416
rect	287	415	288	416
rect	293	415	294	416
rect	303	415	304	416
rect	306	415	307	416
rect	325	415	326	416
rect	328	415	329	416
rect	331	415	332	416
rect	57	416	58	417
rect	63	416	64	417
rect	66	416	67	417
rect	77	416	78	417
rect	81	416	82	417
rect	89	416	90	417
rect	97	416	98	417
rect	100	416	101	417
rect	103	416	104	417
rect	113	416	114	417
rect	124	416	125	417
rect	127	416	128	417
rect	130	416	131	417
rect	133	416	134	417
rect	146	416	147	417
rect	197	416	198	417
rect	200	416	201	417
rect	206	416	207	417
rect	209	416	210	417
rect	212	416	213	417
rect	218	416	219	417
rect	221	416	222	417
rect	237	416	238	417
rect	239	416	240	417
rect	242	416	243	417
rect	251	416	252	417
rect	257	416	258	417
rect	260	416	261	417
rect	262	416	263	417
rect	266	416	267	417
rect	268	416	269	417
rect	275	416	276	417
rect	278	416	279	417
rect	284	416	285	417
rect	287	416	288	417
rect	293	416	294	417
rect	303	416	304	417
rect	306	416	307	417
rect	325	416	326	417
rect	328	416	329	417
rect	331	416	332	417
rect	57	417	58	418
rect	63	417	64	418
rect	66	417	67	418
rect	77	417	78	418
rect	81	417	82	418
rect	89	417	90	418
rect	97	417	98	418
rect	100	417	101	418
rect	103	417	104	418
rect	113	417	114	418
rect	124	417	125	418
rect	127	417	128	418
rect	130	417	131	418
rect	133	417	134	418
rect	146	417	147	418
rect	197	417	198	418
rect	200	417	201	418
rect	206	417	207	418
rect	209	417	210	418
rect	212	417	213	418
rect	218	417	219	418
rect	237	417	238	418
rect	242	417	243	418
rect	251	417	252	418
rect	257	417	258	418
rect	260	417	261	418
rect	262	417	263	418
rect	266	417	267	418
rect	268	417	269	418
rect	275	417	276	418
rect	278	417	279	418
rect	284	417	285	418
rect	287	417	288	418
rect	293	417	294	418
rect	303	417	304	418
rect	325	417	326	418
rect	328	417	329	418
rect	331	417	332	418
rect	57	418	58	419
rect	63	418	64	419
rect	66	418	67	419
rect	74	418	75	419
rect	77	418	78	419
rect	81	418	82	419
rect	89	418	90	419
rect	97	418	98	419
rect	100	418	101	419
rect	103	418	104	419
rect	113	418	114	419
rect	124	418	125	419
rect	127	418	128	419
rect	130	418	131	419
rect	133	418	134	419
rect	146	418	147	419
rect	197	418	198	419
rect	200	418	201	419
rect	206	418	207	419
rect	209	418	210	419
rect	212	418	213	419
rect	218	418	219	419
rect	231	418	232	419
rect	237	418	238	419
rect	242	418	243	419
rect	251	418	252	419
rect	253	418	254	419
rect	257	418	258	419
rect	260	418	261	419
rect	262	418	263	419
rect	266	418	267	419
rect	268	418	269	419
rect	275	418	276	419
rect	278	418	279	419
rect	284	418	285	419
rect	287	418	288	419
rect	293	418	294	419
rect	303	418	304	419
rect	325	418	326	419
rect	328	418	329	419
rect	331	418	332	419
rect	57	419	58	420
rect	63	419	64	420
rect	74	419	75	420
rect	77	419	78	420
rect	81	419	82	420
rect	89	419	90	420
rect	97	419	98	420
rect	100	419	101	420
rect	103	419	104	420
rect	113	419	114	420
rect	124	419	125	420
rect	127	419	128	420
rect	130	419	131	420
rect	133	419	134	420
rect	146	419	147	420
rect	197	419	198	420
rect	200	419	201	420
rect	209	419	210	420
rect	212	419	213	420
rect	218	419	219	420
rect	231	419	232	420
rect	237	419	238	420
rect	242	419	243	420
rect	251	419	252	420
rect	253	419	254	420
rect	257	419	258	420
rect	260	419	261	420
rect	262	419	263	420
rect	266	419	267	420
rect	268	419	269	420
rect	278	419	279	420
rect	284	419	285	420
rect	287	419	288	420
rect	293	419	294	420
rect	325	419	326	420
rect	328	419	329	420
rect	331	419	332	420
rect	57	420	58	421
rect	63	420	64	421
rect	74	420	75	421
rect	77	420	78	421
rect	81	420	82	421
rect	89	420	90	421
rect	97	420	98	421
rect	100	420	101	421
rect	103	420	104	421
rect	113	420	114	421
rect	124	420	125	421
rect	127	420	128	421
rect	130	420	131	421
rect	133	420	134	421
rect	146	420	147	421
rect	197	420	198	421
rect	200	420	201	421
rect	209	420	210	421
rect	212	420	213	421
rect	218	420	219	421
rect	224	420	225	421
rect	231	420	232	421
rect	237	420	238	421
rect	242	420	243	421
rect	251	420	252	421
rect	253	420	254	421
rect	257	420	258	421
rect	260	420	261	421
rect	262	420	263	421
rect	266	420	267	421
rect	268	420	269	421
rect	278	420	279	421
rect	281	420	282	421
rect	284	420	285	421
rect	287	420	288	421
rect	293	420	294	421
rect	325	420	326	421
rect	328	420	329	421
rect	331	420	332	421
rect	57	421	58	422
rect	63	421	64	422
rect	74	421	75	422
rect	77	421	78	422
rect	81	421	82	422
rect	89	421	90	422
rect	97	421	98	422
rect	100	421	101	422
rect	103	421	104	422
rect	113	421	114	422
rect	124	421	125	422
rect	127	421	128	422
rect	133	421	134	422
rect	146	421	147	422
rect	200	421	201	422
rect	209	421	210	422
rect	212	421	213	422
rect	224	421	225	422
rect	231	421	232	422
rect	237	421	238	422
rect	251	421	252	422
rect	253	421	254	422
rect	257	421	258	422
rect	260	421	261	422
rect	262	421	263	422
rect	266	421	267	422
rect	268	421	269	422
rect	278	421	279	422
rect	281	421	282	422
rect	284	421	285	422
rect	287	421	288	422
rect	293	421	294	422
rect	328	421	329	422
rect	331	421	332	422
rect	57	422	58	423
rect	63	422	64	423
rect	74	422	75	423
rect	77	422	78	423
rect	81	422	82	423
rect	89	422	90	423
rect	97	422	98	423
rect	100	422	101	423
rect	103	422	104	423
rect	107	422	108	423
rect	113	422	114	423
rect	124	422	125	423
rect	127	422	128	423
rect	133	422	134	423
rect	146	422	147	423
rect	186	422	187	423
rect	200	422	201	423
rect	205	422	206	423
rect	209	422	210	423
rect	212	422	213	423
rect	221	422	222	423
rect	224	422	225	423
rect	231	422	232	423
rect	237	422	238	423
rect	247	422	248	423
rect	251	422	252	423
rect	253	422	254	423
rect	257	422	258	423
rect	260	422	261	423
rect	262	422	263	423
rect	266	422	267	423
rect	268	422	269	423
rect	278	422	279	423
rect	281	422	282	423
rect	284	422	285	423
rect	287	422	288	423
rect	293	422	294	423
rect	328	422	329	423
rect	331	422	332	423
rect	57	423	58	424
rect	63	423	64	424
rect	74	423	75	424
rect	77	423	78	424
rect	81	423	82	424
rect	89	423	90	424
rect	97	423	98	424
rect	100	423	101	424
rect	107	423	108	424
rect	113	423	114	424
rect	124	423	125	424
rect	127	423	128	424
rect	133	423	134	424
rect	186	423	187	424
rect	205	423	206	424
rect	221	423	222	424
rect	224	423	225	424
rect	231	423	232	424
rect	237	423	238	424
rect	247	423	248	424
rect	253	423	254	424
rect	262	423	263	424
rect	268	423	269	424
rect	281	423	282	424
rect	328	423	329	424
rect	331	423	332	424
rect	57	424	58	425
rect	63	424	64	425
rect	74	424	75	425
rect	77	424	78	425
rect	81	424	82	425
rect	89	424	90	425
rect	97	424	98	425
rect	100	424	101	425
rect	107	424	108	425
rect	113	424	114	425
rect	124	424	125	425
rect	127	424	128	425
rect	133	424	134	425
rect	186	424	187	425
rect	196	424	197	425
rect	205	424	206	425
rect	218	424	219	425
rect	221	424	222	425
rect	224	424	225	425
rect	231	424	232	425
rect	237	424	238	425
rect	247	424	248	425
rect	253	424	254	425
rect	262	424	263	425
rect	265	424	266	425
rect	268	424	269	425
rect	281	424	282	425
rect	328	424	329	425
rect	331	424	332	425
rect	57	425	58	426
rect	63	425	64	426
rect	74	425	75	426
rect	77	425	78	426
rect	81	425	82	426
rect	89	425	90	426
rect	97	425	98	426
rect	107	425	108	426
rect	113	425	114	426
rect	124	425	125	426
rect	127	425	128	426
rect	133	425	134	426
rect	186	425	187	426
rect	196	425	197	426
rect	205	425	206	426
rect	218	425	219	426
rect	221	425	222	426
rect	224	425	225	426
rect	231	425	232	426
rect	237	425	238	426
rect	247	425	248	426
rect	253	425	254	426
rect	262	425	263	426
rect	265	425	266	426
rect	268	425	269	426
rect	281	425	282	426
rect	331	425	332	426
rect	57	426	58	427
rect	63	426	64	427
rect	74	426	75	427
rect	77	426	78	427
rect	81	426	82	427
rect	89	426	90	427
rect	97	426	98	427
rect	107	426	108	427
rect	110	426	111	427
rect	113	426	114	427
rect	120	426	121	427
rect	124	426	125	427
rect	127	426	128	427
rect	133	426	134	427
rect	186	426	187	427
rect	196	426	197	427
rect	205	426	206	427
rect	218	426	219	427
rect	221	426	222	427
rect	224	426	225	427
rect	231	426	232	427
rect	237	426	238	427
rect	247	426	248	427
rect	253	426	254	427
rect	262	426	263	427
rect	265	426	266	427
rect	268	426	269	427
rect	281	426	282	427
rect	331	426	332	427
rect	74	427	75	428
rect	77	427	78	428
rect	89	427	90	428
rect	107	427	108	428
rect	110	427	111	428
rect	113	427	114	428
rect	120	427	121	428
rect	186	427	187	428
rect	196	427	197	428
rect	205	427	206	428
rect	218	427	219	428
rect	221	427	222	428
rect	224	427	225	428
rect	231	427	232	428
rect	237	427	238	428
rect	247	427	248	428
rect	253	427	254	428
rect	262	427	263	428
rect	265	427	266	428
rect	268	427	269	428
rect	281	427	282	428
rect	74	428	75	429
rect	77	428	78	429
rect	80	428	81	429
rect	89	428	90	429
rect	98	428	99	429
rect	101	428	102	429
rect	107	428	108	429
rect	110	428	111	429
rect	113	428	114	429
rect	120	428	121	429
rect	186	428	187	429
rect	190	428	191	429
rect	196	428	197	429
rect	205	428	206	429
rect	218	428	219	429
rect	221	428	222	429
rect	224	428	225	429
rect	231	428	232	429
rect	237	428	238	429
rect	247	428	248	429
rect	253	428	254	429
rect	262	428	263	429
rect	265	428	266	429
rect	268	428	269	429
rect	281	428	282	429
rect	71	435	72	436
rect	77	435	78	436
rect	80	435	81	436
rect	86	435	87	436
rect	89	435	90	436
rect	95	435	96	436
rect	98	435	99	436
rect	107	435	108	436
rect	110	435	111	436
rect	116	435	117	436
rect	196	435	197	436
rect	202	435	203	436
rect	205	435	206	436
rect	218	435	219	436
rect	221	435	222	436
rect	224	435	225	436
rect	227	435	228	436
rect	231	435	232	436
rect	237	435	238	436
rect	247	435	248	436
rect	250	435	251	436
rect	253	435	254	436
rect	259	435	260	436
rect	262	435	263	436
rect	265	435	266	436
rect	281	435	282	436
rect	77	436	78	437
rect	86	436	87	437
rect	89	436	90	437
rect	95	436	96	437
rect	98	436	99	437
rect	107	436	108	437
rect	110	436	111	437
rect	116	436	117	437
rect	196	436	197	437
rect	202	436	203	437
rect	205	436	206	437
rect	218	436	219	437
rect	221	436	222	437
rect	224	436	225	437
rect	227	436	228	437
rect	231	436	232	437
rect	237	436	238	437
rect	247	436	248	437
rect	250	436	251	437
rect	253	436	254	437
rect	259	436	260	437
rect	262	436	263	437
rect	265	436	266	437
rect	281	436	282	437
rect	77	437	78	438
rect	86	437	87	438
rect	89	437	90	438
rect	95	437	96	438
rect	98	437	99	438
rect	107	437	108	438
rect	110	437	111	438
rect	116	437	117	438
rect	196	437	197	438
rect	202	437	203	438
rect	205	437	206	438
rect	218	437	219	438
rect	221	437	222	438
rect	224	437	225	438
rect	227	437	228	438
rect	231	437	232	438
rect	237	437	238	438
rect	247	437	248	438
rect	250	437	251	438
rect	253	437	254	438
rect	259	437	260	438
rect	262	437	263	438
rect	265	437	266	438
rect	281	437	282	438
rect	77	438	78	439
rect	86	438	87	439
rect	89	438	90	439
rect	95	438	96	439
rect	98	438	99	439
rect	107	438	108	439
rect	110	438	111	439
rect	116	438	117	439
rect	196	438	197	439
rect	202	438	203	439
rect	205	438	206	439
rect	218	438	219	439
rect	221	438	222	439
rect	224	438	225	439
rect	227	438	228	439
rect	231	438	232	439
rect	237	438	238	439
rect	247	438	248	439
rect	250	438	251	439
rect	253	438	254	439
rect	259	438	260	439
rect	262	438	263	439
rect	265	438	266	439
rect	281	438	282	439
rect	77	439	78	440
rect	81	439	82	440
rect	86	439	87	440
rect	89	439	90	440
rect	95	439	96	440
rect	98	439	99	440
rect	107	439	108	440
rect	110	439	111	440
rect	116	439	117	440
rect	167	439	168	440
rect	196	439	197	440
rect	202	439	203	440
rect	205	439	206	440
rect	218	439	219	440
rect	221	439	222	440
rect	224	439	225	440
rect	227	439	228	440
rect	231	439	232	440
rect	237	439	238	440
rect	247	439	248	440
rect	250	439	251	440
rect	253	439	254	440
rect	259	439	260	440
rect	262	439	263	440
rect	265	439	266	440
rect	281	439	282	440
rect	81	440	82	441
rect	89	440	90	441
rect	95	440	96	441
rect	107	440	108	441
rect	116	440	117	441
rect	167	440	168	441
rect	196	440	197	441
rect	202	440	203	441
rect	205	440	206	441
rect	218	440	219	441
rect	221	440	222	441
rect	227	440	228	441
rect	231	440	232	441
rect	237	440	238	441
rect	247	440	248	441
rect	253	440	254	441
rect	259	440	260	441
rect	262	440	263	441
rect	281	440	282	441
rect	81	441	82	442
rect	89	441	90	442
rect	95	441	96	442
rect	101	441	102	442
rect	107	441	108	442
rect	116	441	117	442
rect	167	441	168	442
rect	196	441	197	442
rect	202	441	203	442
rect	205	441	206	442
rect	218	441	219	442
rect	221	441	222	442
rect	227	441	228	442
rect	231	441	232	442
rect	237	441	238	442
rect	247	441	248	442
rect	253	441	254	442
rect	259	441	260	442
rect	262	441	263	442
rect	281	441	282	442
rect	81	442	82	443
rect	101	442	102	443
rect	107	442	108	443
rect	116	442	117	443
rect	167	442	168	443
rect	202	442	203	443
rect	205	442	206	443
rect	218	442	219	443
rect	221	442	222	443
rect	227	442	228	443
rect	281	442	282	443
rect	78	443	79	444
rect	81	443	82	444
rect	101	443	102	444
rect	107	443	108	444
rect	116	443	117	444
rect	167	443	168	444
rect	202	443	203	444
rect	205	443	206	444
rect	218	443	219	444
rect	221	443	222	444
rect	227	443	228	444
rect	281	443	282	444
rect	78	444	79	445
rect	81	444	82	445
rect	101	444	102	445
rect	167	444	168	445
rect	32	445	33	446
rect	78	445	79	446
rect	81	445	82	446
rect	98	445	99	446
rect	101	445	102	446
rect	167	445	168	446
rect	98	452	99	453
rect	101	452	102	453
rect	104	452	105	453
rect	107	452	108	453
rect	98	453	99	454
rect	104	453	105	454
rect	98	454	99	455
rect	104	454	105	455
<< via >>
rect	69	0	70	1
rect	72	0	73	1
rect	56	2	57	3
rect	131	2	132	3
rect	190	2	191	3
rect	193	2	194	3
rect	43	4	44	5
rect	109	4	110	5
rect	118	4	119	5
rect	124	4	125	5
rect	173	4	174	5
rect	220	4	221	5
rect	237	4	238	5
rect	243	4	244	5
rect	246	4	247	5
rect	252	4	253	5
rect	262	4	263	5
rect	265	4	266	5
rect	32	13	33	14
rect	252	13	253	14
rect	180	15	181	16
rect	182	15	183	16
rect	190	15	191	16
rect	191	15	192	16
rect	246	15	247	16
rect	253	15	254	16
rect	108	17	109	18
rect	109	17	110	18
rect	179	17	180	18
rect	200	17	201	18
rect	220	17	221	18
rect	221	17	222	18
rect	243	17	244	18
rect	265	17	266	18
rect	95	19	96	20
rect	118	19	119	20
rect	167	19	168	20
rect	170	19	171	20
rect	177	19	178	20
rect	200	19	201	20
rect	209	19	210	20
rect	278	19	279	20
rect	53	21	54	22
rect	56	21	57	22
rect	71	21	72	22
rect	72	21	73	22
rect	85	21	86	22
rect	131	21	132	22
rect	163	21	164	22
rect	256	21	257	22
rect	285	21	286	22
rect	302	21	303	22
rect	11	23	12	24
rect	14	23	15	24
rect	29	23	30	24
rect	30	23	31	24
rect	50	23	51	24
rect	53	23	54	24
rect	62	23	63	24
rect	125	23	126	24
rect	142	23	143	24
rect	152	23	153	24
rect	161	23	162	24
rect	214	23	215	24
rect	218	23	219	24
rect	227	23	228	24
rect	244	23	245	24
rect	247	23	248	24
rect	262	23	263	24
rect	296	23	297	24
rect	11	25	12	26
rect	164	25	165	26
rect	170	25	171	26
rect	176	25	177	26
rect	188	25	189	26
rect	305	25	306	26
rect	215	34	216	35
rect	218	34	219	35
rect	203	36	204	37
rect	218	36	219	37
rect	200	38	201	39
rect	203	38	204	39
rect	197	40	198	41
rect	309	40	310	41
rect	176	42	177	43
rect	200	42	201	43
rect	265	42	266	43
rect	276	42	277	43
rect	173	44	174	45
rect	197	44	198	45
rect	261	44	262	45
rect	273	44	274	45
rect	167	46	168	47
rect	176	46	177	47
rect	231	46	232	47
rect	246	46	247	47
rect	258	46	259	47
rect	270	46	271	47
rect	164	48	165	49
rect	173	48	174	49
rect	227	48	228	49
rect	233	48	234	49
rect	250	48	251	49
rect	300	48	301	49
rect	119	50	120	51
rect	122	50	123	51
rect	152	50	153	51
rect	167	50	168	51
rect	170	50	171	51
rect	182	50	183	51
rect	206	50	207	51
rect	209	50	210	51
rect	221	50	222	51
rect	230	50	231	51
rect	240	50	241	51
rect	288	50	289	51
rect	305	50	306	51
rect	330	50	331	51
rect	56	52	57	53
rect	62	52	63	53
rect	77	52	78	53
rect	267	52	268	53
rect	302	52	303	53
rect	339	52	340	53
rect	53	54	54	55
rect	62	54	63	55
rect	71	54	72	55
rect	80	54	81	55
rect	108	54	109	55
rect	110	54	111	55
rect	114	54	115	55
rect	128	54	129	55
rect	149	54	150	55
rect	158	54	159	55
rect	164	54	165	55
rect	179	54	180	55
rect	188	54	189	55
rect	191	54	192	55
rect	194	54	195	55
rect	357	54	358	55
rect	34	56	35	57
rect	179	56	180	57
rect	191	56	192	57
rect	244	56	245	57
rect	249	56	250	57
rect	253	56	254	57
rect	256	56	257	57
rect	264	56	265	57
rect	278	56	279	57
rect	279	56	280	57
rect	297	56	298	57
rect	306	56	307	57
rect	14	58	15	59
rect	21	58	22	59
rect	30	58	31	59
rect	37	58	38	59
rect	47	58	48	59
rect	53	58	54	59
rect	71	58	72	59
rect	141	58	142	59
rect	146	58	147	59
rect	318	58	319	59
rect	321	58	322	59
rect	333	58	334	59
rect	348	58	349	59
rect	354	58	355	59
rect	357	67	358	68
rect	396	67	397	68
rect	339	69	340	70
rect	357	69	358	70
rect	330	71	331	72
rect	339	71	340	72
rect	294	73	295	74
rect	330	73	331	74
rect	288	75	289	76
rect	315	75	316	76
rect	200	77	201	78
rect	324	77	325	78
rect	167	79	168	80
rect	200	79	201	80
rect	249	79	250	80
rect	252	79	253	80
rect	264	79	265	80
rect	294	79	295	80
rect	148	81	149	82
rect	188	81	189	82
rect	227	81	228	82
rect	249	81	250	82
rect	261	81	262	82
rect	291	81	292	82
rect	164	83	165	84
rect	188	83	189	84
rect	218	83	219	84
rect	228	83	229	84
rect	258	83	259	84
rect	288	83	289	84
rect	161	85	162	86
rect	164	85	165	86
rect	167	85	168	86
rect	170	85	171	86
rect	194	85	195	86
rect	270	85	271	86
rect	297	85	298	86
rect	333	85	334	86
rect	348	85	349	86
rect	369	85	370	86
rect	53	87	54	88
rect	59	87	60	88
rect	68	87	69	88
rect	71	87	72	88
rect	77	87	78	88
rect	112	87	113	88
rect	138	87	139	88
rect	148	87	149	88
rect	158	87	159	88
rect	194	87	195	88
rect	203	87	204	88
rect	225	87	226	88
rect	255	87	256	88
rect	306	87	307	88
rect	318	87	319	88
rect	348	87	349	88
rect	37	89	38	90
rect	40	89	41	90
rect	50	89	51	90
rect	203	89	204	90
rect	215	89	216	90
rect	219	89	220	90
rect	230	89	231	90
rect	264	89	265	90
rect	276	89	277	90
rect	297	89	298	90
rect	318	89	319	90
rect	321	89	322	90
rect	34	91	35	92
rect	37	91	38	92
rect	50	91	51	92
rect	56	91	57	92
rect	62	91	63	92
rect	77	91	78	92
rect	80	91	81	92
rect	86	91	87	92
rect	119	91	120	92
rect	130	91	131	92
rect	136	91	137	92
rect	139	91	140	92
rect	142	91	143	92
rect	360	91	361	92
rect	21	93	22	94
rect	28	93	29	94
rect	31	93	32	94
rect	89	93	90	94
rect	110	93	111	94
rect	121	93	122	94
rect	128	93	129	94
rect	151	93	152	94
rect	155	93	156	94
rect	191	93	192	94
rect	197	93	198	94
rect	222	93	223	94
rect	231	93	232	94
rect	255	93	256	94
rect	258	93	259	94
rect	261	93	262	94
rect	267	93	268	94
rect	273	93	274	94
rect	276	93	277	94
rect	279	93	280	94
rect	309	93	310	94
rect	321	93	322	94
rect	11	95	12	96
rect	170	95	171	96
rect	197	95	198	96
rect	206	95	207	96
rect	209	95	210	96
rect	240	95	241	96
rect	246	95	247	96
rect	267	95	268	96
rect	279	95	280	96
rect	285	95	286	96
rect	300	95	301	96
rect	336	95	337	96
rect	378	95	379	96
rect	381	95	382	96
rect	384	95	385	96
rect	387	95	388	96
rect	213	104	214	105
rect	219	104	220	105
rect	339	104	340	105
rect	342	104	343	105
rect	378	104	379	105
rect	419	104	420	105
rect	203	106	204	107
rect	219	106	220	107
rect	267	106	268	107
rect	279	106	280	107
rect	297	106	298	107
rect	303	106	304	107
rect	330	106	331	107
rect	402	106	403	107
rect	185	108	186	109
rect	204	108	205	109
rect	261	108	262	109
rect	297	108	298	109
rect	300	108	301	109
rect	306	108	307	109
rect	336	108	337	109
rect	378	108	379	109
rect	387	108	388	109
rect	402	108	403	109
rect	183	110	184	111
rect	188	110	189	111
rect	191	110	192	111
rect	213	110	214	111
rect	249	110	250	111
rect	261	110	262	111
rect	264	110	265	111
rect	312	110	313	111
rect	321	110	322	111
rect	339	110	340	111
rect	351	110	352	111
rect	387	110	388	111
rect	173	112	174	113
rect	189	112	190	113
rect	194	112	195	113
rect	216	112	217	113
rect	222	112	223	113
rect	243	112	244	113
rect	246	112	247	113
rect	252	112	253	113
rect	264	112	265	113
rect	276	112	277	113
rect	294	112	295	113
rect	351	112	352	113
rect	357	112	358	113
rect	372	112	373	113
rect	151	114	152	115
rect	174	114	175	115
rect	179	114	180	115
rect	195	114	196	115
rect	200	114	201	115
rect	222	114	223	115
rect	228	114	229	115
rect	234	114	235	115
rect	240	114	241	115
rect	276	114	277	115
rect	285	114	286	115
rect	336	114	337	115
rect	345	114	346	115
rect	369	114	370	115
rect	89	116	90	117
rect	92	116	93	117
rect	112	116	113	117
rect	118	116	119	117
rect	148	116	149	117
rect	155	116	156	117
rect	176	116	177	117
rect	192	116	193	117
rect	197	116	198	117
rect	207	116	208	117
rect	225	116	226	117
rect	267	116	268	117
rect	273	116	274	117
rect	285	116	286	117
rect	294	116	295	117
rect	309	116	310	117
rect	315	116	316	117
rect	363	116	364	117
rect	40	118	41	119
rect	42	118	43	119
rect	59	118	60	119
rect	70	118	71	119
rect	86	118	87	119
rect	89	118	90	119
rect	109	118	110	119
rect	115	118	116	119
rect	121	118	122	119
rect	127	118	128	119
rect	130	118	131	119
rect	136	118	137	119
rect	139	118	140	119
rect	152	118	153	119
rect	170	118	171	119
rect	177	118	178	119
rect	186	118	187	119
rect	357	118	358	119
rect	37	120	38	121
rect	39	120	40	121
rect	56	120	57	121
rect	58	120	59	121
rect	61	120	62	121
rect	68	120	69	121
rect	77	120	78	121
rect	86	120	87	121
rect	95	120	96	121
rect	321	120	322	121
rect	333	120	334	121
rect	366	120	367	121
rect	31	122	32	123
rect	158	122	159	123
rect	167	122	168	123
rect	210	122	211	123
rect	225	122	226	123
rect	231	122	232	123
rect	237	122	238	123
rect	315	122	316	123
rect	318	122	319	123
rect	333	122	334	123
rect	360	122	361	123
rect	369	122	370	123
rect	18	124	19	125
rect	21	124	22	125
rect	28	124	29	125
rect	30	124	31	125
rect	34	124	35	125
rect	249	124	250	125
rect	270	124	271	125
rect	282	124	283	125
rect	291	124	292	125
rect	318	124	319	125
rect	354	124	355	125
rect	360	124	361	125
rect	396	124	397	125
rect	416	124	417	125
rect	11	126	12	127
rect	252	126	253	127
rect	258	126	259	127
rect	273	126	274	127
rect	288	126	289	127
rect	300	126	301	127
rect	327	126	328	127
rect	330	126	331	127
rect	348	126	349	127
rect	396	126	397	127
rect	216	135	217	136
rect	231	135	232	136
rect	201	137	202	138
rect	210	137	211	138
rect	216	137	217	138
rect	225	137	226	138
rect	237	137	238	138
rect	261	137	262	138
rect	306	137	307	138
rect	315	137	316	138
rect	149	139	150	140
rect	267	139	268	140
rect	276	139	277	140
rect	288	139	289	140
rect	297	139	298	140
rect	315	139	316	140
rect	183	141	184	142
rect	207	141	208	142
rect	225	141	226	142
rect	228	141	229	142
rect	234	141	235	142
rect	255	141	256	142
rect	267	141	268	142
rect	273	141	274	142
rect	276	141	277	142
rect	279	141	280	142
rect	291	141	292	142
rect	300	141	301	142
rect	318	141	319	142
rect	327	141	328	142
rect	189	143	190	144
rect	207	143	208	144
rect	222	143	223	144
rect	234	143	235	144
rect	243	143	244	144
rect	261	143	262	144
rect	264	143	265	144
rect	279	143	280	144
rect	285	143	286	144
rect	297	143	298	144
rect	312	143	313	144
rect	324	143	325	144
rect	351	143	352	144
rect	352	143	353	144
rect	369	143	370	144
rect	382	143	383	144
rect	92	145	93	146
rect	98	145	99	146
rect	158	145	159	146
rect	167	145	168	146
rect	180	145	181	146
rect	410	145	411	146
rect	89	147	90	148
rect	95	147	96	148
rect	136	147	137	148
rect	140	147	141	148
rect	158	147	159	148
rect	300	147	301	148
rect	312	147	313	148
rect	330	147	331	148
rect	346	147	347	148
rect	357	147	358	148
rect	366	147	367	148
rect	373	147	374	148
rect	42	149	43	150
rect	47	149	48	150
rect	86	149	87	150
rect	107	149	108	150
rect	118	149	119	150
rect	119	149	120	150
rect	127	149	128	150
rect	137	149	138	150
rect	155	149	156	150
rect	164	149	165	150
rect	177	149	178	150
rect	189	149	190	150
rect	192	149	193	150
rect	210	149	211	150
rect	213	149	214	150
rect	228	149	229	150
rect	237	149	238	150
rect	246	149	247	150
rect	252	149	253	150
rect	264	149	265	150
rect	273	149	274	150
rect	294	149	295	150
rect	309	149	310	150
rect	333	149	334	150
rect	342	149	343	150
rect	349	149	350	150
rect	354	149	355	150
rect	370	149	371	150
rect	36	151	37	152
rect	112	151	113	152
rect	115	151	116	152
rect	116	151	117	152
rect	128	151	129	152
rect	130	151	131	152
rect	152	151	153	152
rect	161	151	162	152
rect	174	151	175	152
rect	192	151	193	152
rect	195	151	196	152
rect	213	151	214	152
rect	219	151	220	152
rect	246	151	247	152
rect	249	151	250	152
rect	258	151	259	152
rect	282	151	283	152
rect	294	151	295	152
rect	303	151	304	152
rect	318	151	319	152
rect	321	151	322	152
rect	330	151	331	152
rect	339	151	340	152
rect	367	151	368	152
rect	21	153	22	154
rect	55	153	56	154
rect	58	153	59	154
rect	65	153	66	154
rect	75	153	76	154
rect	358	153	359	154
rect	387	153	388	154
rect	391	153	392	154
rect	396	153	397	154
rect	402	153	403	154
rect	30	155	31	156
rect	35	155	36	156
rect	39	155	40	156
rect	44	155	45	156
rect	56	155	57	156
rect	61	155	62	156
rect	70	155	71	156
rect	324	155	325	156
rect	336	155	337	156
rect	355	155	356	156
rect	363	155	364	156
rect	375	155	376	156
rect	378	155	379	156
rect	394	155	395	156
rect	413	155	414	156
rect	419	155	420	156
rect	248	164	249	165
rect	273	164	274	165
rect	276	164	277	165
rect	281	164	282	165
rect	330	164	331	165
rect	332	164	333	165
rect	242	166	243	167
rect	246	166	247	167
rect	275	166	276	167
rect	309	166	310	167
rect	318	166	319	167
rect	329	166	330	167
rect	245	168	246	169
rect	255	168	256	169
rect	269	168	270	169
rect	279	168	280	169
rect	306	168	307	169
rect	321	168	322	169
rect	231	170	232	171
rect	251	170	252	171
rect	264	170	265	171
rect	278	170	279	171
rect	297	170	298	171
rect	305	170	306	171
rect	315	170	316	171
rect	317	170	318	171
rect	207	172	208	173
rect	230	172	231	173
rect	234	172	235	173
rect	254	172	255	173
rect	258	172	259	173
rect	266	172	267	173
rect	272	172	273	173
rect	373	172	374	173
rect	50	174	51	175
rect	291	174	292	175
rect	294	174	295	175
rect	314	174	315	175
rect	149	176	150	177
rect	152	176	153	177
rect	192	176	193	177
rect	208	176	209	177
rect	219	176	220	177
rect	290	176	291	177
rect	293	176	294	177
rect	312	176	313	177
rect	353	176	354	177
rect	367	176	368	177
rect	137	178	138	179
rect	149	178	150	179
rect	177	178	178	179
rect	183	178	184	179
rect	192	178	193	179
rect	201	178	202	179
rect	204	178	205	179
rect	205	178	206	179
rect	213	178	214	179
rect	233	178	234	179
rect	237	178	238	179
rect	257	178	258	179
rect	263	178	264	179
rect	327	178	328	179
rect	344	178	345	179
rect	349	178	350	179
rect	358	178	359	179
rect	359	178	360	179
rect	368	178	369	179
rect	382	178	383	179
rect	42	180	43	181
rect	44	180	45	181
rect	128	180	129	181
rect	137	180	138	181
rect	167	180	168	181
rect	168	180	169	181
rect	173	180	174	181
rect	284	180	285	181
rect	288	180	289	181
rect	296	180	297	181
rect	341	180	342	181
rect	346	180	347	181
rect	356	180	357	181
rect	370	180	371	181
rect	394	180	395	181
rect	397	180	398	181
rect	35	182	36	183
rect	45	182	46	183
rect	98	182	99	183
rect	100	182	101	183
rect	119	182	120	183
rect	128	182	129	183
rect	164	182	165	183
rect	174	182	175	183
rect	183	182	184	183
rect	186	182	187	183
rect	189	182	190	183
rect	202	182	203	183
rect	210	182	211	183
rect	211	182	212	183
rect	214	182	215	183
rect	216	182	217	183
rect	220	182	221	183
rect	225	182	226	183
rect	228	182	229	183
rect	240	182	241	183
rect	261	182	262	183
rect	371	182	372	183
rect	388	182	389	183
rect	391	182	392	183
rect	394	182	395	183
rect	413	182	414	183
rect	8	184	9	185
rect	14	184	15	185
rect	29	184	30	185
rect	30	184	31	185
rect	36	184	37	185
rect	39	184	40	185
rect	47	184	48	185
rect	48	184	49	185
rect	51	184	52	185
rect	56	184	57	185
rect	65	184	66	185
rect	67	184	68	185
rect	95	184	96	185
rect	97	184	98	185
rect	107	184	108	185
rect	119	184	120	185
rect	161	184	162	185
rect	171	184	172	185
rect	186	184	187	185
rect	303	184	304	185
rect	326	184	327	185
rect	388	184	389	185
rect	391	184	392	185
rect	410	184	411	185
rect	312	193	313	194
rect	332	193	333	194
rect	310	195	311	196
rect	326	195	327	196
rect	205	197	206	198
rect	227	197	228	198
rect	317	197	318	198
rect	325	197	326	198
rect	206	199	207	200
rect	214	199	215	200
rect	316	199	317	200
rect	320	199	321	200
rect	211	201	212	202
rect	215	201	216	202
rect	242	201	243	202
rect	260	201	261	202
rect	319	201	320	202
rect	344	201	345	202
rect	48	203	49	204
rect	56	203	57	204
rect	212	203	213	204
rect	248	203	249	204
rect	329	203	330	204
rect	331	203	332	204
rect	343	203	344	204
rect	368	203	369	204
rect	45	205	46	206
rect	53	205	54	206
rect	149	205	150	206
rect	159	205	160	206
rect	249	205	250	206
rect	257	205	258	206
rect	261	205	262	206
rect	266	205	267	206
rect	269	205	270	206
rect	273	205	274	206
rect	281	205	282	206
rect	285	205	286	206
rect	307	205	308	206
rect	341	205	342	206
rect	39	207	40	208
rect	47	207	48	208
rect	100	207	101	208
rect	101	207	102	208
rect	119	207	120	208
rect	126	207	127	208
rect	137	207	138	208
rect	150	207	151	208
rect	180	207	181	208
rect	183	207	184	208
rect	224	207	225	208
rect	245	207	246	208
rect	258	207	259	208
rect	290	207	291	208
rect	304	207	305	208
rect	305	207	306	208
rect	312	207	313	208
rect	328	207	329	208
rect	340	207	341	208
rect	353	207	354	208
rect	27	209	28	210
rect	264	209	265	210
rect	267	209	268	210
rect	293	209	294	210
rect	301	209	302	210
rect	314	209	315	210
rect	322	209	323	210
rect	356	209	357	210
rect	388	209	389	210
rect	397	209	398	210
rect	14	211	15	212
rect	17	211	18	212
rect	26	211	27	212
rect	30	211	31	212
rect	38	211	39	212
rect	51	211	52	212
rect	67	211	68	212
rect	75	211	76	212
rect	97	211	98	212
rect	98	211	99	212
rect	116	211	117	212
rect	117	211	118	212
rect	128	211	129	212
rect	135	211	136	212
rect	138	211	139	212
rect	140	211	141	212
rect	147	211	148	212
rect	152	211	153	212
rect	174	211	175	212
rect	180	211	181	212
rect	233	211	234	212
rect	246	211	247	212
rect	254	211	255	212
rect	338	211	339	212
rect	368	211	369	212
rect	391	211	392	212
rect	8	213	9	214
rect	352	213	353	214
rect	359	213	360	214
rect	371	213	372	214
rect	387	213	388	214
rect	394	213	395	214
rect	8	215	9	216
rect	14	215	15	216
rect	24	215	25	216
rect	35	215	36	216
rect	42	215	43	216
rect	50	215	51	216
rect	61	215	62	216
rect	72	215	73	216
rect	81	215	82	216
rect	162	215	163	216
rect	171	215	172	216
rect	177	215	178	216
rect	202	215	203	216
rect	203	215	204	216
rect	208	215	209	216
rect	227	215	228	216
rect	230	215	231	216
rect	243	215	244	216
rect	251	215	252	216
rect	270	215	271	216
rect	278	215	279	216
rect	282	215	283	216
rect	296	215	297	216
rect	385	215	386	216
rect	240	224	241	225
rect	267	224	268	225
rect	261	226	262	227
rect	266	226	267	227
rect	180	228	181	229
rect	188	228	189	229
rect	249	228	250	229
rect	252	228	253	229
rect	258	228	259	229
rect	276	228	277	229
rect	137	230	138	231
rect	138	230	139	231
rect	150	230	151	231
rect	161	230	162	231
rect	177	230	178	231
rect	185	230	186	231
rect	221	230	222	231
rect	224	230	225	231
rect	248	230	249	231
rect	260	230	261	231
rect	273	230	274	231
rect	275	230	276	231
rect	56	232	57	233
rect	60	232	61	233
rect	135	232	136	233
rect	149	232	150	233
rect	170	232	171	233
rect	179	232	180	233
rect	203	232	204	233
rect	210	232	211	233
rect	215	232	216	233
rect	232	232	233	233
rect	246	232	247	233
rect	272	232	273	233
rect	53	234	54	235
rect	57	234	58	235
rect	101	234	102	235
rect	106	234	107	235
rect	134	234	135	235
rect	147	234	148	235
rect	168	234	169	235
rect	176	234	177	235
rect	197	234	198	235
rect	206	234	207	235
rect	214	234	215	235
rect	220	234	221	235
rect	243	234	244	235
rect	251	234	252	235
rect	325	234	326	235
rect	336	234	337	235
rect	50	236	51	237
rect	54	236	55	237
rect	98	236	99	237
rect	109	236	110	237
rect	117	236	118	237
rect	118	236	119	237
rect	126	236	127	237
rect	140	236	141	237
rect	159	236	160	237
rect	173	236	174	237
rect	193	236	194	237
rect	285	236	286	237
rect	319	236	320	237
rect	334	236	335	237
rect	340	236	341	237
rect	346	236	347	237
rect	47	238	48	239
rect	51	238	52	239
rect	80	238	81	239
rect	158	238	159	239
rect	165	238	166	239
rect	324	238	325	239
rect	328	238	329	239
rect	339	238	340	239
rect	24	240	25	241
rect	26	240	27	241
rect	35	240	36	241
rect	48	240	49	241
rect	75	240	76	241
rect	327	240	328	241
rect	331	240	332	241
rect	362	240	363	241
rect	17	242	18	243
rect	27	242	28	243
rect	30	242	31	243
rect	38	242	39	243
rect	72	242	73	243
rect	83	242	84	243
rect	92	242	93	243
rect	333	242	334	243
rect	343	242	344	243
rect	349	242	350	243
rect	360	242	361	243
rect	368	242	369	243
rect	371	242	372	243
rect	376	242	377	243
rect	14	244	15	245
rect	21	244	22	245
rect	36	244	37	245
rect	39	244	40	245
rect	66	244	67	245
rect	223	244	224	245
rect	227	244	228	245
rect	254	244	255	245
rect	270	244	271	245
rect	287	244	288	245
rect	307	244	308	245
rect	308	244	309	245
rect	316	244	317	245
rect	381	244	382	245
rect	4	246	5	247
rect	257	246	258	247
rect	264	246	265	247
rect	269	246	270	247
rect	282	246	283	247
rect	284	246	285	247
rect	296	246	297	247
rect	301	246	302	247
rect	304	246	305	247
rect	305	246	306	247
rect	310	246	311	247
rect	322	246	323	247
rect	348	246	349	247
rect	352	246	353	247
rect	357	246	358	247
rect	363	246	364	247
rect	370	246	371	247
rect	373	246	374	247
rect	379	246	380	247
rect	387	246	388	247
rect	281	255	282	256
rect	366	255	367	256
rect	179	257	180	258
rect	185	257	186	258
rect	275	257	276	258
rect	280	257	281	258
rect	57	259	58	260
rect	63	259	64	260
rect	158	259	159	260
rect	164	259	165	260
rect	173	259	174	260
rect	200	259	201	260
rect	257	259	258	260
rect	262	259	263	260
rect	266	259	267	260
rect	289	259	290	260
rect	379	259	380	260
rect	381	259	382	260
rect	21	261	22	262
rect	33	261	34	262
rect	54	261	55	262
rect	57	261	58	262
rect	140	261	141	262
rect	151	261	152	262
rect	163	261	164	262
rect	172	261	173	262
rect	176	261	177	262
rect	185	261	186	262
rect	254	261	255	262
rect	265	261	266	262
rect	272	261	273	262
rect	277	261	278	262
rect	284	261	285	262
rect	298	261	299	262
rect	333	261	334	262
rect	341	261	342	262
rect	357	261	358	262
rect	378	261	379	262
rect	21	263	22	264
rect	24	263	25	264
rect	27	263	28	264
rect	36	263	37	264
rect	51	263	52	264
rect	54	263	55	264
rect	60	263	61	264
rect	66	263	67	264
rect	112	263	113	264
rect	124	263	125	264
rect	134	263	135	264
rect	139	263	140	264
rect	161	263	162	264
rect	175	263	176	264
rect	194	263	195	264
rect	320	263	321	264
rect	326	263	327	264
rect	336	263	337	264
rect	339	263	340	264
rect	344	263	345	264
rect	348	263	349	264
rect	360	263	361	264
rect	24	265	25	266
rect	30	265	31	266
rect	39	265	40	266
rect	45	265	46	266
rect	48	265	49	266
rect	75	265	76	266
rect	89	265	90	266
rect	91	265	92	266
rect	103	265	104	266
rect	112	265	113	266
rect	133	265	134	266
rect	142	265	143	266
rect	160	265	161	266
rect	170	265	171	266
rect	191	265	192	266
rect	197	265	198	266
rect	223	265	224	266
rect	227	265	228	266
rect	251	265	252	266
rect	274	265	275	266
rect	283	265	284	266
rect	287	265	288	266
rect	314	265	315	266
rect	363	265	364	266
rect	373	265	374	266
rect	387	265	388	266
rect	4	267	5	268
rect	60	267	61	268
rect	83	267	84	268
rect	100	267	101	268
rect	103	267	104	268
rect	106	267	107	268
rect	109	267	110	268
rect	115	267	116	268
rect	118	267	119	268
rect	127	267	128	268
rect	130	267	131	268
rect	137	267	138	268
rect	149	267	150	268
rect	169	267	170	268
rect	188	267	189	268
rect	194	267	195	268
rect	220	267	221	268
rect	224	267	225	268
rect	232	267	233	268
rect	236	267	237	268
rect	248	267	249	268
rect	259	267	260	268
rect	269	267	270	268
rect	292	267	293	268
rect	296	267	297	268
rect	302	267	303	268
rect	305	267	306	268
rect	317	267	318	268
rect	323	267	324	268
rect	324	267	325	268
rect	329	267	330	268
rect	335	267	336	268
rect	338	267	339	268
rect	357	267	358	268
rect	369	267	370	268
rect	376	267	377	268
rect	292	276	293	277
rect	311	276	312	277
rect	381	276	382	277
rect	387	276	388	277
rect	289	278	290	279
rect	308	278	309	279
rect	338	278	339	279
rect	357	278	358	279
rect	360	278	361	279
rect	381	278	382	279
rect	178	280	179	281
rect	179	280	180	281
rect	188	280	189	281
rect	191	280	192	281
rect	274	280	275	281
rect	308	280	309	281
rect	335	280	336	281
rect	360	280	361	281
rect	63	282	64	283
rect	69	282	70	283
rect	107	282	108	283
rect	115	282	116	283
rect	130	282	131	283
rect	133	282	134	283
rect	145	282	146	283
rect	167	282	168	283
rect	172	282	173	283
rect	182	282	183	283
rect	185	282	186	283
rect	200	282	201	283
rect	274	282	275	283
rect	277	282	278	283
rect	280	282	281	283
rect	292	282	293	283
rect	326	282	327	283
rect	330	282	331	283
rect	336	282	337	283
rect	344	282	345	283
rect	372	282	373	283
rect	393	282	394	283
rect	60	284	61	285
rect	63	284	64	285
rect	66	284	67	285
rect	72	284	73	285
rect	109	284	110	285
rect	112	284	113	285
rect	127	284	128	285
rect	130	284	131	285
rect	142	284	143	285
rect	148	284	149	285
rect	160	284	161	285
rect	164	284	165	285
rect	169	284	170	285
rect	203	284	204	285
rect	206	284	207	285
rect	215	284	216	285
rect	227	284	228	285
rect	230	284	231	285
rect	236	284	237	285
rect	246	284	247	285
rect	259	284	260	285
rect	271	284	272	285
rect	277	284	278	285
rect	283	284	284	285
rect	320	284	321	285
rect	345	284	346	285
rect	366	284	367	285
rect	375	284	376	285
rect	23	286	24	287
rect	24	286	25	287
rect	36	286	37	287
rect	42	286	43	287
rect	57	286	58	287
rect	66	286	67	287
rect	100	286	101	287
rect	112	286	113	287
rect	115	286	116	287
rect	118	286	119	287
rect	124	286	125	287
rect	145	286	146	287
rect	151	286	152	287
rect	170	286	171	287
rect	175	286	176	287
rect	191	286	192	287
rect	197	286	198	287
rect	218	286	219	287
rect	227	286	228	287
rect	236	286	237	287
rect	255	286	256	287
rect	262	286	263	287
rect	265	286	266	287
rect	280	286	281	287
rect	317	286	318	287
rect	318	286	319	287
rect	323	286	324	287
rect	324	286	325	287
rect	333	286	334	287
rect	341	286	342	287
rect	350	286	351	287
rect	354	286	355	287
rect	363	286	364	287
rect	372	286	373	287
rect	1	288	2	289
rect	11	288	12	289
rect	14	288	15	289
rect	21	288	22	289
rect	33	288	34	289
rect	39	288	40	289
rect	45	288	46	289
rect	51	288	52	289
rect	54	288	55	289
rect	60	288	61	289
rect	75	288	76	289
rect	81	288	82	289
rect	91	288	92	289
rect	97	288	98	289
rect	100	288	101	289
rect	103	288	104	289
rect	107	288	108	289
rect	118	288	119	289
rect	121	288	122	289
rect	127	288	128	289
rect	142	288	143	289
rect	151	288	152	289
rect	154	288	155	289
rect	185	288	186	289
rect	194	288	195	289
rect	209	288	210	289
rect	224	288	225	289
rect	351	288	352	289
rect	363	288	364	289
rect	369	288	370	289
rect	133	297	134	298
rect	137	297	138	298
rect	203	297	204	298
rect	242	297	243	298
rect	246	297	247	298
rect	251	297	252	298
rect	130	299	131	300
rect	134	299	135	300
rect	185	299	186	300
rect	203	299	204	300
rect	218	299	219	300
rect	245	299	246	300
rect	112	301	113	302
rect	131	301	132	302
rect	176	301	177	302
rect	185	301	186	302
rect	206	301	207	302
rect	221	301	222	302
rect	287	301	288	302
rect	292	301	293	302
rect	387	301	388	302
rect	394	301	395	302
rect	113	303	114	304
rect	124	303	125	304
rect	176	303	177	304
rect	188	303	189	304
rect	200	303	201	304
rect	218	303	219	304
rect	269	303	270	304
rect	271	303	272	304
rect	280	303	281	304
rect	293	303	294	304
rect	357	303	358	304
rect	388	303	389	304
rect	125	305	126	306
rect	127	305	128	306
rect	139	305	140	306
rect	152	305	153	306
rect	170	305	171	306
rect	188	305	189	306
rect	197	305	198	306
rect	215	305	216	306
rect	233	305	234	306
rect	281	305	282	306
rect	358	305	359	306
rect	363	305	364	306
rect	72	307	73	308
rect	83	307	84	308
rect	95	307	96	308
rect	100	307	101	308
rect	128	307	129	308
rect	148	307	149	308
rect	164	307	165	308
rect	170	307	171	308
rect	191	307	192	308
rect	206	307	207	308
rect	233	307	234	308
rect	239	307	240	308
rect	272	307	273	308
rect	289	307	290	308
rect	348	307	349	308
rect	360	307	361	308
rect	66	309	67	310
rect	77	309	78	310
rect	101	309	102	310
rect	109	309	110	310
rect	121	309	122	310
rect	413	309	414	310
rect	1	311	2	312
rect	14	311	15	312
rect	42	311	43	312
rect	47	311	48	312
rect	63	311	64	312
rect	74	311	75	312
rect	81	311	82	312
rect	92	311	93	312
rect	95	311	96	312
rect	110	311	111	312
rect	122	311	123	312
rect	142	311	143	312
rect	145	311	146	312
rect	155	311	156	312
rect	161	311	162	312
rect	164	311	165	312
rect	182	311	183	312
rect	200	311	201	312
rect	224	311	225	312
rect	361	311	362	312
rect	378	311	379	312
rect	379	311	380	312
rect	4	313	5	314
rect	8	313	9	314
rect	14	313	15	314
rect	23	313	24	314
rect	39	313	40	314
rect	44	313	45	314
rect	51	313	52	314
rect	56	313	57	314
rect	60	313	61	314
rect	65	313	66	314
rect	69	313	70	314
rect	80	313	81	314
rect	97	313	98	314
rect	104	313	105	314
rect	107	313	108	314
rect	115	313	116	314
rect	118	313	119	314
rect	140	313	141	314
rect	146	313	147	314
rect	149	313	150	314
rect	158	313	159	314
rect	173	313	174	314
rect	179	313	180	314
rect	197	313	198	314
rect	209	313	210	314
rect	224	313	225	314
rect	230	313	231	314
rect	236	313	237	314
rect	277	313	278	314
rect	290	313	291	314
rect	335	313	336	314
rect	336	313	337	314
rect	354	313	355	314
rect	366	313	367	314
rect	372	313	373	314
rect	384	313	385	314
rect	390	313	391	314
rect	410	313	411	314
rect	4	315	5	316
rect	212	315	213	316
rect	227	315	228	316
rect	248	315	249	316
rect	255	315	256	316
rect	260	315	261	316
rect	274	315	275	316
rect	284	315	285	316
rect	308	315	309	316
rect	311	315	312	316
rect	323	315	324	316
rect	324	315	325	316
rect	332	315	333	316
rect	333	315	334	316
rect	345	315	346	316
rect	370	315	371	316
rect	375	315	376	316
rect	391	315	392	316
rect	400	315	401	316
rect	419	315	420	316
rect	213	324	214	325
rect	230	324	231	325
rect	229	326	230	327
rect	236	326	237	327
rect	147	328	148	329
rect	173	328	174	329
rect	213	328	214	329
rect	235	328	236	329
rect	293	328	294	329
rect	348	328	349	329
rect	174	330	175	331
rect	191	330	192	331
rect	226	330	227	331
rect	233	330	234	331
rect	305	330	306	331
rect	323	330	324	331
rect	349	330	350	331
rect	361	330	362	331
rect	192	332	193	333
rect	200	332	201	333
rect	232	332	233	333
rect	248	332	249	333
rect	256	332	257	333
rect	260	332	261	333
rect	323	332	324	333
rect	361	332	362	333
rect	201	334	202	335
rect	215	334	216	335
rect	245	334	246	335
rect	247	334	248	335
rect	259	334	260	335
rect	269	334	270	335
rect	277	334	278	335
rect	281	334	282	335
rect	320	334	321	335
rect	332	334	333	335
rect	346	334	347	335
rect	358	334	359	335
rect	131	336	132	337
rect	333	336	334	337
rect	358	336	359	337
rect	379	336	380	337
rect	382	336	383	337
rect	388	336	389	337
rect	83	338	84	339
rect	87	338	88	339
rect	132	338	133	339
rect	152	338	153	339
rect	170	338	171	339
rect	183	338	184	339
rect	195	338	196	339
rect	203	338	204	339
rect	206	338	207	339
rect	210	338	211	339
rect	216	338	217	339
rect	410	338	411	339
rect	80	340	81	341
rect	84	340	85	341
rect	99	340	100	341
rect	104	340	105	341
rect	113	340	114	341
rect	114	340	115	341
rect	144	340	145	341
rect	149	340	150	341
rect	153	340	154	341
rect	155	340	156	341
rect	171	340	172	341
rect	197	340	198	341
rect	207	340	208	341
rect	221	340	222	341
rect	244	340	245	341
rect	251	340	252	341
rect	268	340	269	341
rect	287	340	288	341
rect	311	340	312	341
rect	382	340	383	341
rect	72	342	73	343
rect	101	342	102	343
rect	105	342	106	343
rect	122	342	123	343
rect	134	342	135	343
rect	378	342	379	343
rect	77	344	78	345
rect	81	344	82	345
rect	102	344	103	345
rect	107	344	108	345
rect	110	344	111	345
rect	123	344	124	345
rect	128	344	129	345
rect	135	344	136	345
rect	150	344	151	345
rect	176	344	177	345
rect	204	344	205	345
rect	218	344	219	345
rect	224	344	225	345
rect	343	344	344	345
rect	47	346	48	347
rect	54	346	55	347
rect	65	346	66	347
rect	78	346	79	347
rect	96	346	97	347
rect	116	346	117	347
rect	125	346	126	347
rect	126	346	127	347
rect	140	346	141	347
rect	156	346	157	347
rect	167	346	168	347
rect	168	346	169	347
rect	179	346	180	347
rect	180	346	181	347
rect	198	346	199	347
rect	272	346	273	347
rect	280	346	281	347
rect	284	346	285	347
rect	289	346	290	347
rect	290	346	291	347
rect	308	346	309	347
rect	335	346	336	347
rect	394	346	395	347
rect	395	346	396	347
rect	7	348	8	349
rect	14	348	15	349
rect	44	348	45	349
rect	51	348	52	349
rect	56	348	57	349
rect	63	348	64	349
rect	74	348	75	349
rect	75	348	76	349
rect	92	348	93	349
rect	129	348	130	349
rect	137	348	138	349
rect	138	348	139	349
rect	164	348	165	349
rect	165	348	166	349
rect	177	348	178	349
rect	185	348	186	349
rect	188	348	189	349
rect	338	348	339	349
rect	370	348	371	349
rect	376	348	377	349
rect	391	348	392	349
rect	400	348	401	349
rect	416	348	417	349
rect	419	348	420	349
rect	159	357	160	358
rect	165	357	166	358
rect	156	359	157	360
rect	274	359	275	360
rect	91	361	92	362
rect	99	361	100	362
rect	118	361	119	362
rect	132	361	133	362
rect	157	361	158	362
rect	183	361	184	362
rect	78	363	79	364
rect	213	363	214	364
rect	241	363	242	364
rect	280	363	281	364
rect	295	363	296	364
rect	323	363	324	364
rect	72	365	73	366
rect	79	365	80	366
rect	84	365	85	366
rect	94	365	95	366
rect	133	365	134	366
rect	168	365	169	366
rect	189	365	190	366
rect	244	365	245	366
rect	283	365	284	366
rect	311	365	312	366
rect	73	367	74	368
rect	75	367	76	368
rect	81	367	82	368
rect	326	367	327	368
rect	76	369	77	370
rect	105	369	106	370
rect	130	369	131	370
rect	150	369	151	370
rect	153	369	154	370
rect	164	369	165	370
rect	167	369	168	370
rect	195	369	196	370
rect	280	369	281	370
rect	320	369	321	370
rect	323	369	324	370
rect	349	369	350	370
rect	70	371	71	372
rect	102	371	103	372
rect	145	371	146	372
rect	147	371	148	372
rect	151	371	152	372
rect	171	371	172	372
rect	186	371	187	372
rect	192	371	193	372
rect	201	371	202	372
rect	210	371	211	372
rect	220	371	221	372
rect	232	371	233	372
rect	244	371	245	372
rect	268	371	269	372
rect	271	371	272	372
rect	326	371	327	372
rect	348	371	349	372
rect	358	371	359	372
rect	4	373	5	374
rect	20	373	21	374
rect	67	373	68	374
rect	96	373	97	374
rect	106	373	107	374
rect	114	373	115	374
rect	121	373	122	374
rect	135	373	136	374
rect	148	373	149	374
rect	180	373	181	374
rect	192	373	193	374
rect	207	373	208	374
rect	217	373	218	374
rect	229	373	230	374
rect	232	373	233	374
rect	247	373	248	374
rect	253	373	254	374
rect	256	373	257	374
rect	268	373	269	374
rect	308	373	309	374
rect	332	373	333	374
rect	375	373	376	374
rect	4	375	5	376
rect	7	375	8	376
rect	54	375	55	376
rect	351	375	352	376
rect	364	375	365	376
rect	395	375	396	376
rect	8	377	9	378
rect	138	377	139	378
rect	142	377	143	378
rect	177	377	178	378
rect	186	377	187	378
rect	259	377	260	378
rect	265	377	266	378
rect	305	377	306	378
rect	311	377	312	378
rect	317	377	318	378
rect	320	377	321	378
rect	371	377	372	378
rect	10	379	11	380
rect	14	379	15	380
rect	51	379	52	380
rect	58	379	59	380
rect	63	379	64	380
rect	82	379	83	380
rect	87	379	88	380
rect	97	379	98	380
rect	115	379	116	380
rect	123	379	124	380
rect	139	379	140	380
rect	174	379	175	380
rect	183	379	184	380
rect	204	379	205	380
rect	223	379	224	380
rect	226	379	227	380
rect	229	379	230	380
rect	235	379	236	380
rect	256	379	257	380
rect	277	379	278	380
rect	286	379	287	380
rect	289	379	290	380
rect	298	379	299	380
rect	346	379	347	380
rect	361	379	362	380
rect	392	379	393	380
rect	277	388	278	389
rect	286	388	287	389
rect	263	390	264	391
rect	283	390	284	391
rect	287	390	288	391
rect	323	390	324	391
rect	121	392	122	393
rect	127	392	128	393
rect	212	392	213	393
rect	241	392	242	393
rect	260	392	261	393
rect	311	392	312	393
rect	121	394	122	395
rect	139	394	140	395
rect	242	394	243	395
rect	271	394	272	395
rect	284	394	285	395
rect	332	394	333	395
rect	112	396	113	397
rect	130	396	131	397
rect	140	396	141	397
rect	215	396	216	397
rect	227	396	228	397
rect	265	396	266	397
rect	280	396	281	397
rect	289	396	290	397
rect	293	396	294	397
rect	354	396	355	397
rect	130	398	131	399
rect	148	398	149	399
rect	201	398	202	399
rect	206	398	207	399
rect	209	398	210	399
rect	229	398	230	399
rect	239	398	240	399
rect	253	398	254	399
rect	256	398	257	399
rect	266	398	267	399
rect	275	398	276	399
rect	320	398	321	399
rect	331	398	332	399
rect	364	398	365	399
rect	63	400	64	401
rect	70	400	71	401
rect	81	400	82	401
rect	82	400	83	401
rect	97	400	98	401
rect	306	400	307	401
rect	312	400	313	401
rect	318	400	319	401
rect	328	400	329	401
rect	348	400	349	401
rect	60	402	61	403
rect	67	402	68	403
rect	76	402	77	403
rect	84	402	85	403
rect	97	402	98	403
rect	106	402	107	403
rect	118	402	119	403
rect	124	402	125	403
rect	127	402	128	403
rect	145	402	146	403
rect	197	402	198	403
rect	217	402	218	403
rect	220	402	221	403
rect	221	402	222	403
rect	230	402	231	403
rect	232	402	233	403
rect	236	402	237	403
rect	268	402	269	403
rect	272	402	273	403
rect	338	402	339	403
rect	4	404	5	405
rect	8	404	9	405
rect	14	404	15	405
rect	20	404	21	405
rect	58	404	59	405
rect	66	404	67	405
rect	73	404	74	405
rect	75	404	76	405
rect	78	404	79	405
rect	79	404	80	405
rect	94	404	95	405
rect	100	404	101	405
rect	109	404	110	405
rect	115	404	116	405
rect	124	404	125	405
rect	142	404	143	405
rect	146	404	147	405
rect	151	404	152	405
rect	167	404	168	405
rect	173	404	174	405
rect	180	404	181	405
rect	183	404	184	405
rect	192	404	193	405
rect	200	404	201	405
rect	218	404	219	405
rect	244	404	245	405
rect	251	404	252	405
rect	295	404	296	405
rect	303	404	304	405
rect	345	404	346	405
rect	72	413	73	414
rect	78	413	79	414
rect	89	413	90	414
rect	112	413	113	414
rect	237	413	238	414
rect	263	413	264	414
rect	268	413	269	414
rect	312	413	313	414
rect	75	415	76	416
rect	77	415	78	416
rect	109	415	110	416
rect	113	415	114	416
rect	118	415	119	416
rect	121	415	122	416
rect	143	415	144	416
rect	230	415	231	416
rect	262	415	263	416
rect	297	415	298	416
rect	74	417	75	418
rect	221	417	222	418
rect	231	417	232	418
rect	239	417	240	418
rect	253	417	254	418
rect	306	417	307	418
rect	66	419	67	420
rect	206	419	207	420
rect	224	419	225	420
rect	275	419	276	420
rect	281	419	282	420
rect	303	419	304	420
rect	107	421	108	422
rect	130	421	131	422
rect	186	421	187	422
rect	197	421	198	422
rect	205	421	206	422
rect	218	421	219	422
rect	221	421	222	422
rect	242	421	243	422
rect	247	421	248	422
rect	325	421	326	422
rect	103	423	104	424
rect	146	423	147	424
rect	196	423	197	424
rect	200	423	201	424
rect	209	423	210	424
rect	212	423	213	424
rect	218	423	219	424
rect	251	423	252	424
rect	257	423	258	424
rect	260	423	261	424
rect	265	423	266	424
rect	266	423	267	424
rect	278	423	279	424
rect	284	423	285	424
rect	287	423	288	424
rect	293	423	294	424
rect	100	425	101	426
rect	110	425	111	426
rect	120	425	121	426
rect	328	425	329	426
rect	57	427	58	428
rect	63	427	64	428
rect	80	427	81	428
rect	81	427	82	428
rect	97	427	98	428
rect	98	427	99	428
rect	101	427	102	428
rect	124	427	125	428
rect	127	427	128	428
rect	133	427	134	428
rect	190	427	191	428
rect	331	427	332	428
rect	71	436	72	437
rect	80	436	81	437
rect	81	438	82	439
rect	167	438	168	439
rect	77	440	78	441
rect	86	440	87	441
rect	98	440	99	441
rect	101	440	102	441
rect	110	440	111	441
rect	224	440	225	441
rect	250	440	251	441
rect	265	440	266	441
rect	78	442	79	443
rect	89	442	90	443
rect	95	442	96	443
rect	196	442	197	443
rect	231	442	232	443
rect	237	442	238	443
rect	247	442	248	443
rect	253	442	254	443
rect	259	442	260	443
rect	262	442	263	443
rect	32	444	33	445
rect	98	444	99	445
rect	107	444	108	445
rect	116	444	117	445
rect	202	444	203	445
rect	205	444	206	445
rect	218	444	219	445
rect	221	444	222	445
rect	227	444	228	445
rect	281	444	282	445
rect	101	453	102	454
rect	107	453	108	454
rect	98	455	99	456
rect	104	455	105	456
