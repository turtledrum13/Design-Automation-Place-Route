magic
tech scmos
timestamp
<< pdiffusion >>
rect	0	9	6	15
rect	0	69	6	75
rect	17	9	23	15
rect	56	69	62	75
rect	0	35	6	41
rect	0	97	6	103
rect	29	35	35	41
rect	20	97	26	103
rect	10	9	16	15
rect	31	69	37	75
rect	27	9	33	15
rect	78	69	84	75
rect	13	35	19	41
rect	10	97	16	103
rect	54	35	60	41
rect	27	97	33	103
rect	0	22	6	28
rect	0	84	6	90
rect	17	22	23	28
rect	35	84	41	90
rect	0	52	6	58
rect	3	110	9	116
rect	35	52	41	58
rect	37	9	43	15
rect	94	69	100	75
rect	60	9	66	15
rect	123	69	129	75
rect	82	35	88	41
rect	37	97	43	103
rect	105	35	111	41
rect	51	97	57	103
rect	47	9	53	15
rect	107	69	113	75
rect	73	9	79	15
rect	130	69	136	75
rect	95	35	101	41
rect	44	97	50	103
rect	112	35	118	41
rect	67	97	73	103
rect	46	22	52	28
rect	82	84	88	90
rect	75	22	81	28
rect	105	84	111	90
rect	67	52	73	58
rect	31	110	37	116
rect	65	22	68	28
rect	6	35	9	41
rect	23	22	26	28
rect	111	84	114	90
rect	6	9	9	15
rect	9	35	12	41
rect	55	84	58	90
rect	41	84	44	90
rect	66	9	69	15
rect	57	97	60	103
rect	53	9	56	15
rect	113	69	116	75
rect	101	84	104	90
rect	31	22	34	28
rect	41	52	44	58
rect	60	35	63	41
rect	116	69	119	75
rect	6	69	9	75
rect	19	35	22	41
rect	23	9	26	15
rect	44	52	47	58
rect	16	97	19	103
rect	88	35	91	41
rect	127	52	130	58
rect	26	22	29	28
rect	14	84	17	90
rect	34	22	37	28
rect	37	69	40	75
rect	33	9	36	15
rect	59	84	62	90
rect	28	84	31	90
rect	100	69	103	75
rect	40	69	43	75
rect	0	110	3	116
rect	69	84	72	90
rect	62	84	65	90
rect	9	69	12	75
rect	33	97	36	103
rect	31	84	34	90
rect	56	9	59	15
rect	6	97	9	103
rect	91	35	94	41
rect	63	35	66	41
rect	66	35	69	41
rect	10	52	13	58
rect	22	35	25	41
rect	136	69	139	75
rect	7	22	10	28
rect	13	52	16	58
rect	62	69	65	75
rect	65	69	68	75
rect	68	22	71	28
rect	88	84	91	90
rect	93	84	96	90
rect	119	69	122	75
rect	35	35	38	41
rect	73	52	76	58
rect	117	52	120	58
rect	7	84	10	90
rect	38	35	41	41
rect	23	84	26	90
rect	107	52	110	58
rect	41	35	44	41
rect	12	69	15	75
rect	44	35	47	41
rect	84	69	87	75
rect	15	69	18	75
rect	72	84	75	90
rect	87	69	90	75
rect	16	52	19	58
rect	44	84	47	90
rect	43	69	46	75
rect	60	22	63	28
rect	10	84	13	90
rect	113	52	116	58
rect	88	52	91	58
rect	91	52	94	58
rect	18	69	21	75
rect	47	52	50	58
rect	140	52	143	58
rect	21	69	24	75
rect	76	52	79	58
rect	69	35	72	41
rect	90	69	93	75
rect	91	97	94	103
rect	123	52	126	58
rect	101	35	104	41
rect	24	69	27	75
rect	57	52	60	58
rect	19	52	22	58
rect	79	52	82	58
rect	6	52	9	58
rect	60	97	63	103
rect	46	69	49	75
rect	50	52	53	58
rect	72	35	75	41
rect	27	69	30	75
rect	103	69	106	75
rect	68	69	71	75
rect	71	69	74	75
rect	19	84	22	90
rect	49	69	52	75
rect	75	35	78	41
rect	82	52	85	58
rect	94	52	97	58
rect	127	35	130	41
rect	102	22	105	28
rect	25	52	28	58
rect	52	69	55	75
rect	25	35	28	41
rect	53	52	56	58
rect	78	35	81	41
rect	28	52	31	58
rect	75	84	78	90
rect	78	84	81	90
rect	50	84	53	90
rect	71	22	74	28
rect	74	69	77	75
rect	131	22	134	28
rect	47	35	50	41
rect	82	22	85	28
rect	50	35	53	41
rect	76	97	79	103
rect	79	97	82	103
rect	69	9	72	15
rect	65	84	68	90
rect	52	22	55	28
rect	42	22	45	28
rect	77	110	80	116
rect	63	97	66	103
rect	43	9	46	15
