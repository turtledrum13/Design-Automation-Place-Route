magic
tech scmos
timestamp
<< pdiffusion >>
rect	0	5	6	11
rect	0	35	6	41
rect	17	5	23	11
rect	56	35	62	41
rect	0	21	6	27
rect	0	49	6	55
rect	29	21	35	27
rect	20	49	26	55
rect	10	5	16	11
rect	31	35	37	41
rect	27	5	33	11
rect	78	35	84	41
rect	13	21	19	27
rect	10	49	16	55
rect	54	21	60	27
rect	27	49	33	55
rect	0	12	6	18
rect	0	42	6	48
rect	17	12	23	18
rect	35	42	41	48
rect	0	28	6	34
rect	3	56	9	62
rect	35	28	41	34
rect	37	5	43	11
rect	94	35	100	41
rect	60	5	66	11
rect	123	35	129	41
rect	82	21	88	27
rect	37	49	43	55
rect	105	21	111	27
rect	51	49	57	55
rect	47	5	53	11
rect	107	35	113	41
rect	73	5	79	11
rect	130	35	136	41
rect	95	21	101	27
rect	44	49	50	55
rect	112	21	118	27
rect	67	49	73	55
rect	46	12	52	18
rect	82	42	88	48
rect	75	12	81	18
rect	105	42	111	48
rect	67	28	73	34
rect	31	56	37	62
rect	65	12	68	18
rect	6	21	9	27
rect	23	12	26	18
rect	111	42	114	48
rect	6	5	9	11
rect	9	21	12	27
rect	55	42	58	48
rect	41	42	44	48
rect	66	5	69	11
rect	57	49	60	55
rect	53	5	56	11
rect	113	35	116	41
rect	101	42	104	48
rect	31	12	34	18
rect	41	28	44	34
rect	60	21	63	27
rect	116	35	119	41
rect	6	35	9	41
rect	19	21	22	27
rect	23	5	26	11
rect	44	28	47	34
rect	16	49	19	55
rect	88	21	91	27
rect	127	28	130	34
rect	26	12	29	18
rect	14	42	17	48
rect	34	12	37	18
rect	37	35	40	41
rect	33	5	36	11
rect	59	42	62	48
rect	28	42	31	48
rect	100	35	103	41
rect	40	35	43	41
rect	0	56	3	62
rect	69	42	72	48
rect	62	42	65	48
rect	9	35	12	41
rect	33	49	36	55
rect	31	42	34	48
rect	56	5	59	11
rect	6	49	9	55
rect	91	21	94	27
rect	63	21	66	27
rect	66	21	69	27
rect	10	28	13	34
rect	22	21	25	27
rect	136	35	139	41
rect	7	12	10	18
rect	13	28	16	34
rect	62	35	65	41
rect	65	35	68	41
rect	68	12	71	18
rect	88	42	91	48
rect	93	42	96	48
rect	119	35	122	41
rect	35	21	38	27
rect	73	28	76	34
rect	117	28	120	34
rect	7	42	10	48
rect	38	21	41	27
rect	23	42	26	48
rect	107	28	110	34
rect	41	21	44	27
rect	12	35	15	41
rect	44	21	47	27
rect	84	35	87	41
rect	15	35	18	41
rect	72	42	75	48
rect	87	35	90	41
rect	16	28	19	34
rect	44	42	47	48
rect	43	35	46	41
rect	60	12	63	18
rect	10	42	13	48
rect	113	28	116	34
rect	88	28	91	34
rect	91	28	94	34
rect	18	35	21	41
rect	47	28	50	34
rect	140	28	143	34
rect	21	35	24	41
rect	76	28	79	34
rect	69	21	72	27
rect	90	35	93	41
rect	91	49	94	55
rect	123	28	126	34
rect	101	21	104	27
rect	24	35	27	41
rect	57	28	60	34
rect	19	28	22	34
rect	79	28	82	34
rect	6	28	9	34
rect	60	49	63	55
rect	46	35	49	41
rect	50	28	53	34
rect	72	21	75	27
rect	27	35	30	41
rect	103	35	106	41
rect	68	35	71	41
rect	71	35	74	41
rect	19	42	22	48
rect	49	35	52	41
rect	75	21	78	27
rect	82	28	85	34
rect	94	28	97	34
rect	127	21	130	27
rect	102	12	105	18
rect	25	28	28	34
rect	52	35	55	41
rect	25	21	28	27
rect	53	28	56	34
rect	78	21	81	27
rect	28	28	31	34
rect	75	42	78	48
rect	78	42	81	48
rect	50	42	53	48
rect	71	12	74	18
rect	74	35	77	41
rect	131	12	134	18
rect	47	21	50	27
rect	82	12	85	18
rect	50	21	53	27
rect	76	49	79	55
rect	79	49	82	55
rect	69	5	72	11
rect	65	42	68	48
rect	52	12	55	18
rect	42	12	45	18
rect	77	56	80	62
rect	63	49	66	55
rect	43	5	46	11
