magic
tech scmos
timestamp
<< pdiffusion >>
rect	4	0	5	1
rect	4	1	5	2
rect	4	2	5	3
rect	4	3	5	4
rect	4	4	5	5
rect	4	5	5	6
rect	4	6	5	7
rect	4	7	5	8
rect	4	8	5	9
rect	4	9	5	10
rect	4	10	5	11
rect	4	11	5	12
rect	4	12	5	13
rect	4	13	5	14
rect	4	14	5	15
rect	4	15	5	16
rect	4	16	5	17
rect	4	17	5	18
rect	4	18	5	19
rect	4	19	5	20
rect	4	20	5	21
rect	4	21	5	22
rect	4	22	5	23
rect	4	23	5	24
rect	4	24	5	25
rect	4	25	5	26
rect	4	26	5	27
rect	4	27	5	28
rect	4	28	5	29
rect	4	29	5	30
rect	4	30	5	31
rect	4	31	5	32
rect	4	32	5	33
rect	4	33	5	34
rect	4	34	5	35
rect	4	35	5	36
rect	4	36	5	37
rect	4	37	5	38
rect	4	38	5	39
rect	4	39	5	40
rect	4	40	5	41
rect	4	41	5	42
rect	4	42	5	43
rect	4	43	5	44
rect	4	44	5	45
rect	4	45	5	46
rect	4	46	5	47
rect	4	47	5	48
rect	4	48	5	49
rect	4	49	5	50
rect	4	50	5	51
rect	4	51	5	52
rect	4	52	5	53
rect	4	53	5	54
rect	4	54	5	55
rect	4	55	5	56
rect	4	56	5	57
rect	5	0	6	1
rect	5	1	6	2
rect	5	2	6	3
rect	5	3	6	4
rect	5	4	6	5
rect	5	5	6	6
rect	5	6	6	7
rect	5	7	6	8
rect	5	8	6	9
rect	5	9	6	10
rect	5	10	6	11
rect	5	11	6	12
rect	5	12	6	13
rect	5	13	6	14
rect	5	14	6	15
rect	5	15	6	16
rect	5	16	6	17
rect	5	17	6	18
rect	5	18	6	19
rect	5	19	6	20
rect	5	20	6	21
rect	5	21	6	22
rect	5	22	6	23
rect	5	23	6	24
rect	5	24	6	25
rect	5	25	6	26
rect	5	26	6	27
rect	5	27	6	28
rect	5	28	6	29
rect	5	29	6	30
rect	5	30	6	31
rect	5	31	6	32
rect	5	32	6	33
rect	5	33	6	34
rect	5	34	6	35
rect	5	35	6	36
rect	5	36	6	37
rect	5	37	6	38
rect	5	38	6	39
rect	5	39	6	40
rect	5	40	6	41
rect	5	41	6	42
rect	5	42	6	43
rect	5	43	6	44
rect	5	44	6	45
rect	5	45	6	46
rect	5	46	6	47
rect	5	47	6	48
rect	5	48	6	49
rect	5	49	6	50
rect	5	50	6	51
rect	5	51	6	52
rect	5	52	6	53
rect	5	53	6	54
rect	5	54	6	55
rect	5	55	6	56
rect	5	56	6	57
rect	6	0	7	1
rect	6	1	7	2
rect	6	2	7	3
rect	6	3	7	4
rect	6	4	7	5
rect	6	5	7	6
rect	6	6	7	7
rect	6	7	7	8
rect	6	8	7	9
rect	6	9	7	10
rect	6	10	7	11
rect	6	11	7	12
rect	6	12	7	13
rect	6	13	7	14
rect	6	14	7	15
rect	6	15	7	16
rect	6	16	7	17
rect	6	17	7	18
rect	6	18	7	19
rect	6	19	7	20
rect	6	20	7	21
rect	6	21	7	22
rect	6	22	7	23
rect	6	23	7	24
rect	6	24	7	25
rect	6	25	7	26
rect	6	26	7	27
rect	6	27	7	28
rect	6	28	7	29
rect	6	29	7	30
rect	6	30	7	31
rect	6	31	7	32
rect	6	32	7	33
rect	6	33	7	34
rect	6	34	7	35
rect	6	35	7	36
rect	6	36	7	37
rect	6	37	7	38
rect	6	38	7	39
rect	6	39	7	40
rect	6	40	7	41
rect	6	41	7	42
rect	6	42	7	43
rect	6	43	7	44
rect	6	44	7	45
rect	6	45	7	46
rect	6	46	7	47
rect	6	47	7	48
rect	6	48	7	49
rect	6	49	7	50
rect	6	50	7	51
rect	6	51	7	52
rect	6	52	7	53
rect	6	53	7	54
rect	6	54	7	55
rect	6	55	7	56
rect	6	56	7	57
rect	7	0	8	1
rect	7	1	8	2
rect	7	2	8	3
rect	7	3	8	4
rect	7	4	8	5
rect	7	5	8	6
rect	7	6	8	7
rect	7	7	8	8
rect	7	8	8	9
rect	7	9	8	10
rect	7	10	8	11
rect	7	11	8	12
rect	7	12	8	13
rect	7	13	8	14
rect	7	14	8	15
rect	7	15	8	16
rect	7	16	8	17
rect	7	17	8	18
rect	7	18	8	19
rect	7	19	8	20
rect	7	20	8	21
rect	7	21	8	22
rect	7	22	8	23
rect	7	23	8	24
rect	7	24	8	25
rect	7	25	8	26
rect	7	26	8	27
rect	7	27	8	28
rect	7	28	8	29
rect	7	29	8	30
rect	7	30	8	31
rect	7	31	8	32
rect	7	32	8	33
rect	7	33	8	34
rect	7	34	8	35
rect	7	35	8	36
rect	7	36	8	37
rect	7	37	8	38
rect	7	38	8	39
rect	7	39	8	40
rect	7	40	8	41
rect	7	41	8	42
rect	7	42	8	43
rect	7	43	8	44
rect	7	44	8	45
rect	7	45	8	46
rect	7	46	8	47
rect	7	47	8	48
rect	7	48	8	49
rect	7	49	8	50
rect	7	50	8	51
rect	7	51	8	52
rect	7	52	8	53
rect	7	53	8	54
rect	7	54	8	55
rect	7	55	8	56
rect	7	56	8	57
rect	8	0	9	1
rect	8	1	9	2
rect	8	2	9	3
rect	8	3	9	4
rect	8	4	9	5
rect	8	5	9	6
rect	8	6	9	7
rect	8	7	9	8
rect	8	8	9	9
rect	8	9	9	10
rect	8	10	9	11
rect	8	11	9	12
rect	8	12	9	13
rect	8	13	9	14
rect	8	14	9	15
rect	8	15	9	16
rect	8	16	9	17
rect	8	17	9	18
rect	8	18	9	19
rect	8	19	9	20
rect	8	20	9	21
rect	8	21	9	22
rect	8	22	9	23
rect	8	23	9	24
rect	8	24	9	25
rect	8	25	9	26
rect	8	26	9	27
rect	8	27	9	28
rect	8	28	9	29
rect	8	29	9	30
rect	8	30	9	31
rect	8	31	9	32
rect	8	32	9	33
rect	8	33	9	34
rect	8	34	9	35
rect	8	35	9	36
rect	8	36	9	37
rect	8	37	9	38
rect	8	38	9	39
rect	8	39	9	40
rect	8	40	9	41
rect	8	41	9	42
rect	8	42	9	43
rect	8	43	9	44
rect	8	44	9	45
rect	8	45	9	46
rect	8	46	9	47
rect	8	47	9	48
rect	8	48	9	49
rect	8	49	9	50
rect	8	50	9	51
rect	8	51	9	52
rect	8	52	9	53
rect	8	53	9	54
rect	8	54	9	55
rect	8	55	9	56
rect	8	56	9	57
rect	9	0	10	1
rect	9	1	10	2
rect	9	2	10	3
rect	9	3	10	4
rect	9	4	10	5
rect	9	5	10	6
rect	9	6	10	7
rect	9	7	10	8
rect	9	8	10	9
rect	9	9	10	10
rect	9	10	10	11
rect	9	11	10	12
rect	9	12	10	13
rect	9	13	10	14
rect	9	14	10	15
rect	9	15	10	16
rect	9	16	10	17
rect	9	17	10	18
rect	9	18	10	19
rect	9	19	10	20
rect	9	20	10	21
rect	9	21	10	22
rect	9	22	10	23
rect	9	23	10	24
rect	9	24	10	25
rect	9	25	10	26
rect	9	26	10	27
rect	9	27	10	28
rect	9	28	10	29
rect	9	29	10	30
rect	9	30	10	31
rect	9	31	10	32
rect	9	32	10	33
rect	9	33	10	34
rect	9	34	10	35
rect	9	35	10	36
rect	9	36	10	37
rect	9	37	10	38
rect	9	38	10	39
rect	9	39	10	40
rect	9	40	10	41
rect	9	41	10	42
rect	9	42	10	43
rect	9	43	10	44
rect	9	44	10	45
rect	9	45	10	46
rect	9	46	10	47
rect	9	47	10	48
rect	9	48	10	49
rect	9	49	10	50
rect	9	50	10	51
rect	9	51	10	52
rect	9	52	10	53
rect	9	53	10	54
rect	9	54	10	55
rect	9	55	10	56
rect	9	56	10	57
rect	21	0	22	1
rect	21	1	22	2
rect	21	2	22	3
rect	21	3	22	4
rect	21	4	22	5
rect	21	5	22	6
rect	21	6	22	7
rect	21	7	22	8
rect	21	8	22	9
rect	21	9	22	10
rect	21	10	22	11
rect	21	11	22	12
rect	21	12	22	13
rect	21	13	22	14
rect	21	14	22	15
rect	21	15	22	16
rect	21	16	22	17
rect	21	17	22	18
rect	21	18	22	19
rect	21	19	22	20
rect	21	20	22	21
rect	21	21	22	22
rect	21	22	22	23
rect	21	23	22	24
rect	21	24	22	25
rect	21	25	22	26
rect	21	26	22	27
rect	21	27	22	28
rect	21	28	22	29
rect	21	29	22	30
rect	21	30	22	31
rect	21	31	22	32
rect	21	32	22	33
rect	21	33	22	34
rect	21	34	22	35
rect	21	35	22	36
rect	21	36	22	37
rect	21	37	22	38
rect	21	38	22	39
rect	21	39	22	40
rect	21	40	22	41
rect	21	41	22	42
rect	21	42	22	43
rect	21	43	22	44
rect	21	44	22	45
rect	21	45	22	46
rect	21	46	22	47
rect	21	47	22	48
rect	21	48	22	49
rect	21	49	22	50
rect	21	50	22	51
rect	21	51	22	52
rect	21	52	22	53
rect	21	53	22	54
rect	21	54	22	55
rect	21	55	22	56
rect	21	56	22	57
rect	21	57	22	58
rect	21	58	22	59
rect	21	59	22	60
rect	21	60	22	61
rect	21	61	22	62
rect	21	62	22	63
rect	21	63	22	64
rect	21	64	22	65
rect	21	65	22	66
rect	21	66	22	67
rect	21	67	22	68
rect	21	68	22	69
rect	21	69	22	70
rect	21	70	22	71
rect	21	71	22	72
rect	21	72	22	73
rect	21	73	22	74
rect	21	74	22	75
rect	22	0	23	1
rect	22	1	23	2
rect	22	2	23	3
rect	22	3	23	4
rect	22	4	23	5
rect	22	5	23	6
rect	22	6	23	7
rect	22	7	23	8
rect	22	8	23	9
rect	22	9	23	10
rect	22	10	23	11
rect	22	11	23	12
rect	22	12	23	13
rect	22	13	23	14
rect	22	14	23	15
rect	22	15	23	16
rect	22	16	23	17
rect	22	17	23	18
rect	22	18	23	19
rect	22	19	23	20
rect	22	20	23	21
rect	22	21	23	22
rect	22	22	23	23
rect	22	23	23	24
rect	22	24	23	25
rect	22	25	23	26
rect	22	26	23	27
rect	22	27	23	28
rect	22	28	23	29
rect	22	29	23	30
rect	22	30	23	31
rect	22	31	23	32
rect	22	32	23	33
rect	22	33	23	34
rect	22	34	23	35
rect	22	35	23	36
rect	22	36	23	37
rect	22	37	23	38
rect	22	38	23	39
rect	22	39	23	40
rect	22	40	23	41
rect	22	41	23	42
rect	22	42	23	43
rect	22	43	23	44
rect	22	44	23	45
rect	22	45	23	46
rect	22	46	23	47
rect	22	47	23	48
rect	22	48	23	49
rect	22	49	23	50
rect	22	50	23	51
rect	22	51	23	52
rect	22	52	23	53
rect	22	53	23	54
rect	22	54	23	55
rect	22	55	23	56
rect	22	56	23	57
rect	22	57	23	58
rect	22	58	23	59
rect	22	59	23	60
rect	22	60	23	61
rect	22	61	23	62
rect	22	62	23	63
rect	22	63	23	64
rect	22	64	23	65
rect	22	65	23	66
rect	22	66	23	67
rect	22	67	23	68
rect	22	68	23	69
rect	22	69	23	70
rect	22	70	23	71
rect	22	71	23	72
rect	22	72	23	73
rect	22	73	23	74
rect	22	74	23	75
rect	23	0	24	1
rect	23	1	24	2
rect	23	2	24	3
rect	23	3	24	4
rect	23	4	24	5
rect	23	5	24	6
rect	23	6	24	7
rect	23	7	24	8
rect	23	8	24	9
rect	23	9	24	10
rect	23	10	24	11
rect	23	11	24	12
rect	23	12	24	13
rect	23	13	24	14
rect	23	14	24	15
rect	23	15	24	16
rect	23	16	24	17
rect	23	17	24	18
rect	23	18	24	19
rect	23	19	24	20
rect	23	20	24	21
rect	23	21	24	22
rect	23	22	24	23
rect	23	23	24	24
rect	23	24	24	25
rect	23	25	24	26
rect	23	26	24	27
rect	23	27	24	28
rect	23	28	24	29
rect	23	29	24	30
rect	23	30	24	31
rect	23	31	24	32
rect	23	32	24	33
rect	23	33	24	34
rect	23	34	24	35
rect	23	35	24	36
rect	23	36	24	37
rect	23	37	24	38
rect	23	38	24	39
rect	23	39	24	40
rect	23	40	24	41
rect	23	41	24	42
rect	23	42	24	43
rect	23	43	24	44
rect	23	44	24	45
rect	23	45	24	46
rect	23	46	24	47
rect	23	47	24	48
rect	23	48	24	49
rect	23	49	24	50
rect	23	50	24	51
rect	23	51	24	52
rect	23	52	24	53
rect	23	53	24	54
rect	23	54	24	55
rect	23	55	24	56
rect	23	56	24	57
rect	23	57	24	58
rect	23	58	24	59
rect	23	59	24	60
rect	23	60	24	61
rect	23	61	24	62
rect	23	62	24	63
rect	23	63	24	64
rect	23	64	24	65
rect	23	65	24	66
rect	23	66	24	67
rect	23	67	24	68
rect	23	68	24	69
rect	23	69	24	70
rect	23	70	24	71
rect	23	71	24	72
rect	23	72	24	73
rect	23	73	24	74
rect	23	74	24	75
rect	24	0	25	1
rect	24	1	25	2
rect	24	2	25	3
rect	24	3	25	4
rect	24	4	25	5
rect	24	5	25	6
rect	24	6	25	7
rect	24	7	25	8
rect	24	8	25	9
rect	24	9	25	10
rect	24	10	25	11
rect	24	11	25	12
rect	24	12	25	13
rect	24	13	25	14
rect	24	14	25	15
rect	24	15	25	16
rect	24	16	25	17
rect	24	17	25	18
rect	24	18	25	19
rect	24	19	25	20
rect	24	20	25	21
rect	24	21	25	22
rect	24	22	25	23
rect	24	23	25	24
rect	24	24	25	25
rect	24	25	25	26
rect	24	26	25	27
rect	24	27	25	28
rect	24	28	25	29
rect	24	29	25	30
rect	24	30	25	31
rect	24	31	25	32
rect	24	32	25	33
rect	24	33	25	34
rect	24	34	25	35
rect	24	35	25	36
rect	24	36	25	37
rect	24	37	25	38
rect	24	38	25	39
rect	24	39	25	40
rect	24	40	25	41
rect	24	41	25	42
rect	24	42	25	43
rect	24	43	25	44
rect	24	44	25	45
rect	24	45	25	46
rect	24	46	25	47
rect	24	47	25	48
rect	24	48	25	49
rect	24	49	25	50
rect	24	50	25	51
rect	24	51	25	52
rect	24	52	25	53
rect	24	53	25	54
rect	24	54	25	55
rect	24	55	25	56
rect	24	56	25	57
rect	24	57	25	58
rect	24	58	25	59
rect	24	59	25	60
rect	24	60	25	61
rect	24	61	25	62
rect	24	62	25	63
rect	24	63	25	64
rect	24	64	25	65
rect	24	65	25	66
rect	24	66	25	67
rect	24	67	25	68
rect	24	68	25	69
rect	24	69	25	70
rect	24	70	25	71
rect	24	71	25	72
rect	24	72	25	73
rect	24	73	25	74
rect	24	74	25	75
rect	25	0	26	1
rect	25	1	26	2
rect	25	2	26	3
rect	25	3	26	4
rect	25	4	26	5
rect	25	5	26	6
rect	25	6	26	7
rect	25	7	26	8
rect	25	8	26	9
rect	25	9	26	10
rect	25	10	26	11
rect	25	11	26	12
rect	25	12	26	13
rect	25	13	26	14
rect	25	14	26	15
rect	25	15	26	16
rect	25	16	26	17
rect	25	17	26	18
rect	25	18	26	19
rect	25	19	26	20
rect	25	20	26	21
rect	25	21	26	22
rect	25	22	26	23
rect	25	23	26	24
rect	25	24	26	25
rect	25	25	26	26
rect	25	26	26	27
rect	25	27	26	28
rect	25	28	26	29
rect	25	29	26	30
rect	25	30	26	31
rect	25	31	26	32
rect	25	32	26	33
rect	25	33	26	34
rect	25	34	26	35
rect	25	35	26	36
rect	25	36	26	37
rect	25	37	26	38
rect	25	38	26	39
rect	25	39	26	40
rect	25	40	26	41
rect	25	41	26	42
rect	25	42	26	43
rect	25	43	26	44
rect	25	44	26	45
rect	25	45	26	46
rect	25	46	26	47
rect	25	47	26	48
rect	25	48	26	49
rect	25	49	26	50
rect	25	50	26	51
rect	25	51	26	52
rect	25	52	26	53
rect	25	53	26	54
rect	25	54	26	55
rect	25	55	26	56
rect	25	56	26	57
rect	25	57	26	58
rect	25	58	26	59
rect	25	59	26	60
rect	25	60	26	61
rect	25	61	26	62
rect	25	62	26	63
rect	25	63	26	64
rect	25	64	26	65
rect	25	65	26	66
rect	25	66	26	67
rect	25	67	26	68
rect	25	68	26	69
rect	25	69	26	70
rect	25	70	26	71
rect	25	71	26	72
rect	25	72	26	73
rect	25	73	26	74
rect	25	74	26	75
rect	26	0	27	1
rect	26	1	27	2
rect	26	2	27	3
rect	26	3	27	4
rect	26	4	27	5
rect	26	5	27	6
rect	26	6	27	7
rect	26	7	27	8
rect	26	8	27	9
rect	26	9	27	10
rect	26	10	27	11
rect	26	11	27	12
rect	26	12	27	13
rect	26	13	27	14
rect	26	14	27	15
rect	26	15	27	16
rect	26	16	27	17
rect	26	17	27	18
rect	26	18	27	19
rect	26	19	27	20
rect	26	20	27	21
rect	26	21	27	22
rect	26	22	27	23
rect	26	23	27	24
rect	26	24	27	25
rect	26	25	27	26
rect	26	26	27	27
rect	26	27	27	28
rect	26	28	27	29
rect	26	29	27	30
rect	26	30	27	31
rect	26	31	27	32
rect	26	32	27	33
rect	26	33	27	34
rect	26	34	27	35
rect	26	35	27	36
rect	26	36	27	37
rect	26	37	27	38
rect	26	38	27	39
rect	26	39	27	40
rect	26	40	27	41
rect	26	41	27	42
rect	26	42	27	43
rect	26	43	27	44
rect	26	44	27	45
rect	26	45	27	46
rect	26	46	27	47
rect	26	47	27	48
rect	26	48	27	49
rect	26	49	27	50
rect	26	50	27	51
rect	26	51	27	52
rect	26	52	27	53
rect	26	53	27	54
rect	26	54	27	55
rect	26	55	27	56
rect	26	56	27	57
rect	26	57	27	58
rect	26	58	27	59
rect	26	59	27	60
rect	26	60	27	61
rect	26	61	27	62
rect	26	62	27	63
rect	26	63	27	64
rect	26	64	27	65
rect	26	65	27	66
rect	26	66	27	67
rect	26	67	27	68
rect	26	68	27	69
rect	26	69	27	70
rect	26	70	27	71
rect	26	71	27	72
rect	26	72	27	73
rect	26	73	27	74
rect	26	74	27	75
rect	38	0	39	1
rect	38	1	39	2
rect	38	2	39	3
rect	38	3	39	4
rect	38	4	39	5
rect	38	5	39	6
rect	38	6	39	7
rect	38	7	39	8
rect	38	8	39	9
rect	38	9	39	10
rect	38	10	39	11
rect	38	11	39	12
rect	38	12	39	13
rect	38	13	39	14
rect	38	14	39	15
rect	38	15	39	16
rect	38	16	39	17
rect	38	17	39	18
rect	38	18	39	19
rect	38	19	39	20
rect	38	20	39	21
rect	38	21	39	22
rect	38	22	39	23
rect	38	23	39	24
rect	38	24	39	25
rect	38	25	39	26
rect	38	26	39	27
rect	38	27	39	28
rect	38	28	39	29
rect	38	29	39	30
rect	38	30	39	31
rect	38	31	39	32
rect	38	32	39	33
rect	38	33	39	34
rect	38	34	39	35
rect	38	35	39	36
rect	38	36	39	37
rect	38	37	39	38
rect	38	38	39	39
rect	38	39	39	40
rect	38	40	39	41
rect	38	41	39	42
rect	38	42	39	43
rect	38	43	39	44
rect	38	44	39	45
rect	38	45	39	46
rect	38	46	39	47
rect	38	47	39	48
rect	38	48	39	49
rect	38	49	39	50
rect	38	50	39	51
rect	38	51	39	52
rect	38	52	39	53
rect	38	53	39	54
rect	38	54	39	55
rect	38	55	39	56
rect	38	56	39	57
rect	38	57	39	58
rect	38	58	39	59
rect	38	59	39	60
rect	38	60	39	61
rect	38	61	39	62
rect	38	62	39	63
rect	38	63	39	64
rect	38	64	39	65
rect	38	65	39	66
rect	38	66	39	67
rect	38	67	39	68
rect	38	68	39	69
rect	38	69	39	70
rect	38	70	39	71
rect	38	71	39	72
rect	38	72	39	73
rect	38	73	39	74
rect	38	74	39	75
rect	38	75	39	76
rect	38	76	39	77
rect	38	77	39	78
rect	38	78	39	79
rect	38	79	39	80
rect	38	80	39	81
rect	38	81	39	82
rect	38	82	39	83
rect	38	83	39	84
rect	38	84	39	85
rect	38	85	39	86
rect	38	86	39	87
rect	39	0	40	1
rect	39	1	40	2
rect	39	2	40	3
rect	39	3	40	4
rect	39	4	40	5
rect	39	5	40	6
rect	39	6	40	7
rect	39	7	40	8
rect	39	8	40	9
rect	39	9	40	10
rect	39	10	40	11
rect	39	11	40	12
rect	39	12	40	13
rect	39	13	40	14
rect	39	14	40	15
rect	39	15	40	16
rect	39	16	40	17
rect	39	17	40	18
rect	39	18	40	19
rect	39	19	40	20
rect	39	20	40	21
rect	39	21	40	22
rect	39	22	40	23
rect	39	23	40	24
rect	39	24	40	25
rect	39	25	40	26
rect	39	26	40	27
rect	39	27	40	28
rect	39	28	40	29
rect	39	29	40	30
rect	39	30	40	31
rect	39	31	40	32
rect	39	32	40	33
rect	39	33	40	34
rect	39	34	40	35
rect	39	35	40	36
rect	39	36	40	37
rect	39	37	40	38
rect	39	38	40	39
rect	39	39	40	40
rect	39	40	40	41
rect	39	41	40	42
rect	39	42	40	43
rect	39	43	40	44
rect	39	44	40	45
rect	39	45	40	46
rect	39	46	40	47
rect	39	47	40	48
rect	39	48	40	49
rect	39	49	40	50
rect	39	50	40	51
rect	39	51	40	52
rect	39	52	40	53
rect	39	53	40	54
rect	39	54	40	55
rect	39	55	40	56
rect	39	56	40	57
rect	39	57	40	58
rect	39	58	40	59
rect	39	59	40	60
rect	39	60	40	61
rect	39	61	40	62
rect	39	62	40	63
rect	39	63	40	64
rect	39	64	40	65
rect	39	65	40	66
rect	39	66	40	67
rect	39	67	40	68
rect	39	68	40	69
rect	39	69	40	70
rect	39	70	40	71
rect	39	71	40	72
rect	39	72	40	73
rect	39	73	40	74
rect	39	74	40	75
rect	39	75	40	76
rect	39	76	40	77
rect	39	77	40	78
rect	39	78	40	79
rect	39	79	40	80
rect	39	80	40	81
rect	39	81	40	82
rect	39	82	40	83
rect	39	83	40	84
rect	39	84	40	85
rect	39	85	40	86
rect	39	86	40	87
rect	40	0	41	1
rect	40	1	41	2
rect	40	2	41	3
rect	40	3	41	4
rect	40	4	41	5
rect	40	5	41	6
rect	40	6	41	7
rect	40	7	41	8
rect	40	8	41	9
rect	40	9	41	10
rect	40	10	41	11
rect	40	11	41	12
rect	40	12	41	13
rect	40	13	41	14
rect	40	14	41	15
rect	40	15	41	16
rect	40	16	41	17
rect	40	17	41	18
rect	40	18	41	19
rect	40	19	41	20
rect	40	20	41	21
rect	40	21	41	22
rect	40	22	41	23
rect	40	23	41	24
rect	40	24	41	25
rect	40	25	41	26
rect	40	26	41	27
rect	40	27	41	28
rect	40	28	41	29
rect	40	29	41	30
rect	40	30	41	31
rect	40	31	41	32
rect	40	32	41	33
rect	40	33	41	34
rect	40	34	41	35
rect	40	35	41	36
rect	40	36	41	37
rect	40	37	41	38
rect	40	38	41	39
rect	40	39	41	40
rect	40	40	41	41
rect	40	41	41	42
rect	40	42	41	43
rect	40	43	41	44
rect	40	44	41	45
rect	40	45	41	46
rect	40	46	41	47
rect	40	47	41	48
rect	40	48	41	49
rect	40	49	41	50
rect	40	50	41	51
rect	40	51	41	52
rect	40	52	41	53
rect	40	53	41	54
rect	40	54	41	55
rect	40	55	41	56
rect	40	56	41	57
rect	40	57	41	58
rect	40	58	41	59
rect	40	59	41	60
rect	40	60	41	61
rect	40	61	41	62
rect	40	62	41	63
rect	40	63	41	64
rect	40	64	41	65
rect	40	65	41	66
rect	40	66	41	67
rect	40	67	41	68
rect	40	68	41	69
rect	40	69	41	70
rect	40	70	41	71
rect	40	71	41	72
rect	40	72	41	73
rect	40	73	41	74
rect	40	74	41	75
rect	40	75	41	76
rect	40	76	41	77
rect	40	77	41	78
rect	40	78	41	79
rect	40	79	41	80
rect	40	80	41	81
rect	40	81	41	82
rect	40	82	41	83
rect	40	83	41	84
rect	40	84	41	85
rect	40	85	41	86
rect	40	86	41	87
rect	41	0	42	1
rect	41	1	42	2
rect	41	2	42	3
rect	41	3	42	4
rect	41	4	42	5
rect	41	5	42	6
rect	41	6	42	7
rect	41	7	42	8
rect	41	8	42	9
rect	41	9	42	10
rect	41	10	42	11
rect	41	11	42	12
rect	41	12	42	13
rect	41	13	42	14
rect	41	14	42	15
rect	41	15	42	16
rect	41	16	42	17
rect	41	17	42	18
rect	41	18	42	19
rect	41	19	42	20
rect	41	20	42	21
rect	41	21	42	22
rect	41	22	42	23
rect	41	23	42	24
rect	41	24	42	25
rect	41	25	42	26
rect	41	26	42	27
rect	41	27	42	28
rect	41	28	42	29
rect	41	29	42	30
rect	41	30	42	31
rect	41	31	42	32
rect	41	32	42	33
rect	41	33	42	34
rect	41	34	42	35
rect	41	35	42	36
rect	41	36	42	37
rect	41	37	42	38
rect	41	38	42	39
rect	41	39	42	40
rect	41	40	42	41
rect	41	41	42	42
rect	41	42	42	43
rect	41	43	42	44
rect	41	44	42	45
rect	41	45	42	46
rect	41	46	42	47
rect	41	47	42	48
rect	41	48	42	49
rect	41	49	42	50
rect	41	50	42	51
rect	41	51	42	52
rect	41	52	42	53
rect	41	53	42	54
rect	41	54	42	55
rect	41	55	42	56
rect	41	56	42	57
rect	41	57	42	58
rect	41	58	42	59
rect	41	59	42	60
rect	41	60	42	61
rect	41	61	42	62
rect	41	62	42	63
rect	41	63	42	64
rect	41	64	42	65
rect	41	65	42	66
rect	41	66	42	67
rect	41	67	42	68
rect	41	68	42	69
rect	41	69	42	70
rect	41	70	42	71
rect	41	71	42	72
rect	41	72	42	73
rect	41	73	42	74
rect	41	74	42	75
rect	41	75	42	76
rect	41	76	42	77
rect	41	77	42	78
rect	41	78	42	79
rect	41	79	42	80
rect	41	80	42	81
rect	41	81	42	82
rect	41	82	42	83
rect	41	83	42	84
rect	41	84	42	85
rect	41	85	42	86
rect	41	86	42	87
rect	42	0	43	1
rect	42	1	43	2
rect	42	2	43	3
rect	42	3	43	4
rect	42	4	43	5
rect	42	5	43	6
rect	42	6	43	7
rect	42	7	43	8
rect	42	8	43	9
rect	42	9	43	10
rect	42	10	43	11
rect	42	11	43	12
rect	42	12	43	13
rect	42	13	43	14
rect	42	14	43	15
rect	42	15	43	16
rect	42	16	43	17
rect	42	17	43	18
rect	42	18	43	19
rect	42	19	43	20
rect	42	20	43	21
rect	42	21	43	22
rect	42	22	43	23
rect	42	23	43	24
rect	42	24	43	25
rect	42	25	43	26
rect	42	26	43	27
rect	42	27	43	28
rect	42	28	43	29
rect	42	29	43	30
rect	42	30	43	31
rect	42	31	43	32
rect	42	32	43	33
rect	42	33	43	34
rect	42	34	43	35
rect	42	35	43	36
rect	42	36	43	37
rect	42	37	43	38
rect	42	38	43	39
rect	42	39	43	40
rect	42	40	43	41
rect	42	41	43	42
rect	42	42	43	43
rect	42	43	43	44
rect	42	44	43	45
rect	42	45	43	46
rect	42	46	43	47
rect	42	47	43	48
rect	42	48	43	49
rect	42	49	43	50
rect	42	50	43	51
rect	42	51	43	52
rect	42	52	43	53
rect	42	53	43	54
rect	42	54	43	55
rect	42	55	43	56
rect	42	56	43	57
rect	42	57	43	58
rect	42	58	43	59
rect	42	59	43	60
rect	42	60	43	61
rect	42	61	43	62
rect	42	62	43	63
rect	42	63	43	64
rect	42	64	43	65
rect	42	65	43	66
rect	42	66	43	67
rect	42	67	43	68
rect	42	68	43	69
rect	42	69	43	70
rect	42	70	43	71
rect	42	71	43	72
rect	42	72	43	73
rect	42	73	43	74
rect	42	74	43	75
rect	42	75	43	76
rect	42	76	43	77
rect	42	77	43	78
rect	42	78	43	79
rect	42	79	43	80
rect	42	80	43	81
rect	42	81	43	82
rect	42	82	43	83
rect	42	83	43	84
rect	42	84	43	85
rect	42	85	43	86
rect	42	86	43	87
rect	43	0	44	1
rect	43	1	44	2
rect	43	2	44	3
rect	43	3	44	4
rect	43	4	44	5
rect	43	5	44	6
rect	43	6	44	7
rect	43	7	44	8
rect	43	8	44	9
rect	43	9	44	10
rect	43	10	44	11
rect	43	11	44	12
rect	43	12	44	13
rect	43	13	44	14
rect	43	14	44	15
rect	43	15	44	16
rect	43	16	44	17
rect	43	17	44	18
rect	43	18	44	19
rect	43	19	44	20
rect	43	20	44	21
rect	43	21	44	22
rect	43	22	44	23
rect	43	23	44	24
rect	43	24	44	25
rect	43	25	44	26
rect	43	26	44	27
rect	43	27	44	28
rect	43	28	44	29
rect	43	29	44	30
rect	43	30	44	31
rect	43	31	44	32
rect	43	32	44	33
rect	43	33	44	34
rect	43	34	44	35
rect	43	35	44	36
rect	43	36	44	37
rect	43	37	44	38
rect	43	38	44	39
rect	43	39	44	40
rect	43	40	44	41
rect	43	41	44	42
rect	43	42	44	43
rect	43	43	44	44
rect	43	44	44	45
rect	43	45	44	46
rect	43	46	44	47
rect	43	47	44	48
rect	43	48	44	49
rect	43	49	44	50
rect	43	50	44	51
rect	43	51	44	52
rect	43	52	44	53
rect	43	53	44	54
rect	43	54	44	55
rect	43	55	44	56
rect	43	56	44	57
rect	43	57	44	58
rect	43	58	44	59
rect	43	59	44	60
rect	43	60	44	61
rect	43	61	44	62
rect	43	62	44	63
rect	43	63	44	64
rect	43	64	44	65
rect	43	65	44	66
rect	43	66	44	67
rect	43	67	44	68
rect	43	68	44	69
rect	43	69	44	70
rect	43	70	44	71
rect	43	71	44	72
rect	43	72	44	73
rect	43	73	44	74
rect	43	74	44	75
rect	43	75	44	76
rect	43	76	44	77
rect	43	77	44	78
rect	43	78	44	79
rect	43	79	44	80
rect	43	80	44	81
rect	43	81	44	82
rect	43	82	44	83
rect	43	83	44	84
rect	43	84	44	85
rect	43	85	44	86
rect	43	86	44	87
rect	59	0	60	1
rect	59	1	60	2
rect	59	2	60	3
rect	59	3	60	4
rect	59	4	60	5
rect	59	5	60	6
rect	59	6	60	7
rect	59	7	60	8
rect	59	8	60	9
rect	59	9	60	10
rect	59	10	60	11
rect	59	11	60	12
rect	59	12	60	13
rect	59	13	60	14
rect	59	14	60	15
rect	59	15	60	16
rect	59	16	60	17
rect	59	17	60	18
rect	59	18	60	19
rect	59	19	60	20
rect	59	20	60	21
rect	59	21	60	22
rect	59	22	60	23
rect	59	23	60	24
rect	59	24	60	25
rect	59	25	60	26
rect	59	26	60	27
rect	59	27	60	28
rect	59	28	60	29
rect	59	29	60	30
rect	59	30	60	31
rect	59	31	60	32
rect	59	32	60	33
rect	59	33	60	34
rect	59	34	60	35
rect	59	35	60	36
rect	59	36	60	37
rect	59	37	60	38
rect	59	38	60	39
rect	59	39	60	40
rect	59	40	60	41
rect	59	41	60	42
rect	59	42	60	43
rect	59	43	60	44
rect	59	44	60	45
rect	59	45	60	46
rect	59	46	60	47
rect	59	47	60	48
rect	59	48	60	49
rect	59	49	60	50
rect	59	50	60	51
rect	59	51	60	52
rect	59	52	60	53
rect	59	53	60	54
rect	59	54	60	55
rect	59	55	60	56
rect	59	56	60	57
rect	59	57	60	58
rect	59	58	60	59
rect	59	59	60	60
rect	59	60	60	61
rect	59	61	60	62
rect	59	62	60	63
rect	59	63	60	64
rect	59	64	60	65
rect	59	65	60	66
rect	59	66	60	67
rect	59	67	60	68
rect	59	68	60	69
rect	59	69	60	70
rect	59	70	60	71
rect	59	71	60	72
rect	59	72	60	73
rect	59	73	60	74
rect	59	74	60	75
rect	59	75	60	76
rect	59	76	60	77
rect	59	77	60	78
rect	59	78	60	79
rect	59	79	60	80
rect	59	80	60	81
rect	59	81	60	82
rect	59	82	60	83
rect	59	83	60	84
rect	59	84	60	85
rect	59	85	60	86
rect	59	86	60	87
rect	59	87	60	88
rect	59	88	60	89
rect	59	89	60	90
rect	59	90	60	91
rect	59	91	60	92
rect	59	92	60	93
rect	60	0	61	1
rect	60	1	61	2
rect	60	2	61	3
rect	60	3	61	4
rect	60	4	61	5
rect	60	5	61	6
rect	60	6	61	7
rect	60	7	61	8
rect	60	8	61	9
rect	60	9	61	10
rect	60	10	61	11
rect	60	11	61	12
rect	60	12	61	13
rect	60	13	61	14
rect	60	14	61	15
rect	60	15	61	16
rect	60	16	61	17
rect	60	17	61	18
rect	60	18	61	19
rect	60	19	61	20
rect	60	20	61	21
rect	60	21	61	22
rect	60	22	61	23
rect	60	23	61	24
rect	60	24	61	25
rect	60	25	61	26
rect	60	26	61	27
rect	60	27	61	28
rect	60	28	61	29
rect	60	29	61	30
rect	60	30	61	31
rect	60	31	61	32
rect	60	32	61	33
rect	60	33	61	34
rect	60	34	61	35
rect	60	35	61	36
rect	60	36	61	37
rect	60	37	61	38
rect	60	38	61	39
rect	60	39	61	40
rect	60	40	61	41
rect	60	41	61	42
rect	60	42	61	43
rect	60	43	61	44
rect	60	44	61	45
rect	60	45	61	46
rect	60	46	61	47
rect	60	47	61	48
rect	60	48	61	49
rect	60	49	61	50
rect	60	50	61	51
rect	60	51	61	52
rect	60	52	61	53
rect	60	53	61	54
rect	60	54	61	55
rect	60	55	61	56
rect	60	56	61	57
rect	60	57	61	58
rect	60	58	61	59
rect	60	59	61	60
rect	60	60	61	61
rect	60	61	61	62
rect	60	62	61	63
rect	60	63	61	64
rect	60	64	61	65
rect	60	65	61	66
rect	60	66	61	67
rect	60	67	61	68
rect	60	68	61	69
rect	60	69	61	70
rect	60	70	61	71
rect	60	71	61	72
rect	60	72	61	73
rect	60	73	61	74
rect	60	74	61	75
rect	60	75	61	76
rect	60	76	61	77
rect	60	77	61	78
rect	60	78	61	79
rect	60	79	61	80
rect	60	80	61	81
rect	60	81	61	82
rect	60	82	61	83
rect	60	83	61	84
rect	60	84	61	85
rect	60	85	61	86
rect	60	86	61	87
rect	60	87	61	88
rect	60	88	61	89
rect	60	89	61	90
rect	60	90	61	91
rect	60	91	61	92
rect	60	92	61	93
rect	61	0	62	1
rect	61	1	62	2
rect	61	2	62	3
rect	61	3	62	4
rect	61	4	62	5
rect	61	5	62	6
rect	61	6	62	7
rect	61	7	62	8
rect	61	8	62	9
rect	61	9	62	10
rect	61	10	62	11
rect	61	11	62	12
rect	61	12	62	13
rect	61	13	62	14
rect	61	14	62	15
rect	61	15	62	16
rect	61	16	62	17
rect	61	17	62	18
rect	61	18	62	19
rect	61	19	62	20
rect	61	20	62	21
rect	61	21	62	22
rect	61	22	62	23
rect	61	23	62	24
rect	61	24	62	25
rect	61	25	62	26
rect	61	26	62	27
rect	61	27	62	28
rect	61	28	62	29
rect	61	29	62	30
rect	61	30	62	31
rect	61	31	62	32
rect	61	32	62	33
rect	61	33	62	34
rect	61	34	62	35
rect	61	35	62	36
rect	61	36	62	37
rect	61	37	62	38
rect	61	38	62	39
rect	61	39	62	40
rect	61	40	62	41
rect	61	41	62	42
rect	61	42	62	43
rect	61	43	62	44
rect	61	44	62	45
rect	61	45	62	46
rect	61	46	62	47
rect	61	47	62	48
rect	61	48	62	49
rect	61	49	62	50
rect	61	50	62	51
rect	61	51	62	52
rect	61	52	62	53
rect	61	53	62	54
rect	61	54	62	55
rect	61	55	62	56
rect	61	56	62	57
rect	61	57	62	58
rect	61	58	62	59
rect	61	59	62	60
rect	61	60	62	61
rect	61	61	62	62
rect	61	62	62	63
rect	61	63	62	64
rect	61	64	62	65
rect	61	65	62	66
rect	61	66	62	67
rect	61	67	62	68
rect	61	68	62	69
rect	61	69	62	70
rect	61	70	62	71
rect	61	71	62	72
rect	61	72	62	73
rect	61	73	62	74
rect	61	74	62	75
rect	61	75	62	76
rect	61	76	62	77
rect	61	77	62	78
rect	61	78	62	79
rect	61	79	62	80
rect	61	80	62	81
rect	61	81	62	82
rect	61	82	62	83
rect	61	83	62	84
rect	61	84	62	85
rect	61	85	62	86
rect	61	86	62	87
rect	61	87	62	88
rect	61	88	62	89
rect	61	89	62	90
rect	61	90	62	91
rect	61	91	62	92
rect	61	92	62	93
rect	62	0	63	1
rect	62	1	63	2
rect	62	2	63	3
rect	62	3	63	4
rect	62	4	63	5
rect	62	5	63	6
rect	62	6	63	7
rect	62	7	63	8
rect	62	8	63	9
rect	62	9	63	10
rect	62	10	63	11
rect	62	11	63	12
rect	62	12	63	13
rect	62	13	63	14
rect	62	14	63	15
rect	62	15	63	16
rect	62	16	63	17
rect	62	17	63	18
rect	62	18	63	19
rect	62	19	63	20
rect	62	20	63	21
rect	62	21	63	22
rect	62	22	63	23
rect	62	23	63	24
rect	62	24	63	25
rect	62	25	63	26
rect	62	26	63	27
rect	62	27	63	28
rect	62	28	63	29
rect	62	29	63	30
rect	62	30	63	31
rect	62	31	63	32
rect	62	32	63	33
rect	62	33	63	34
rect	62	34	63	35
rect	62	35	63	36
rect	62	36	63	37
rect	62	37	63	38
rect	62	38	63	39
rect	62	39	63	40
rect	62	40	63	41
rect	62	41	63	42
rect	62	42	63	43
rect	62	43	63	44
rect	62	44	63	45
rect	62	45	63	46
rect	62	46	63	47
rect	62	47	63	48
rect	62	48	63	49
rect	62	49	63	50
rect	62	50	63	51
rect	62	51	63	52
rect	62	52	63	53
rect	62	53	63	54
rect	62	54	63	55
rect	62	55	63	56
rect	62	56	63	57
rect	62	57	63	58
rect	62	58	63	59
rect	62	59	63	60
rect	62	60	63	61
rect	62	61	63	62
rect	62	62	63	63
rect	62	63	63	64
rect	62	64	63	65
rect	62	65	63	66
rect	62	66	63	67
rect	62	67	63	68
rect	62	68	63	69
rect	62	69	63	70
rect	62	70	63	71
rect	62	71	63	72
rect	62	72	63	73
rect	62	73	63	74
rect	62	74	63	75
rect	62	75	63	76
rect	62	76	63	77
rect	62	77	63	78
rect	62	78	63	79
rect	62	79	63	80
rect	62	80	63	81
rect	62	81	63	82
rect	62	82	63	83
rect	62	83	63	84
rect	62	84	63	85
rect	62	85	63	86
rect	62	86	63	87
rect	62	87	63	88
rect	62	88	63	89
rect	62	89	63	90
rect	62	90	63	91
rect	62	91	63	92
rect	62	92	63	93
rect	63	0	64	1
rect	63	1	64	2
rect	63	2	64	3
rect	63	3	64	4
rect	63	4	64	5
rect	63	5	64	6
rect	63	6	64	7
rect	63	7	64	8
rect	63	8	64	9
rect	63	9	64	10
rect	63	10	64	11
rect	63	11	64	12
rect	63	12	64	13
rect	63	13	64	14
rect	63	14	64	15
rect	63	15	64	16
rect	63	16	64	17
rect	63	17	64	18
rect	63	18	64	19
rect	63	19	64	20
rect	63	20	64	21
rect	63	21	64	22
rect	63	22	64	23
rect	63	23	64	24
rect	63	24	64	25
rect	63	25	64	26
rect	63	26	64	27
rect	63	27	64	28
rect	63	28	64	29
rect	63	29	64	30
rect	63	30	64	31
rect	63	31	64	32
rect	63	32	64	33
rect	63	33	64	34
rect	63	34	64	35
rect	63	35	64	36
rect	63	36	64	37
rect	63	37	64	38
rect	63	38	64	39
rect	63	39	64	40
rect	63	40	64	41
rect	63	41	64	42
rect	63	42	64	43
rect	63	43	64	44
rect	63	44	64	45
rect	63	45	64	46
rect	63	46	64	47
rect	63	47	64	48
rect	63	48	64	49
rect	63	49	64	50
rect	63	50	64	51
rect	63	51	64	52
rect	63	52	64	53
rect	63	53	64	54
rect	63	54	64	55
rect	63	55	64	56
rect	63	56	64	57
rect	63	57	64	58
rect	63	58	64	59
rect	63	59	64	60
rect	63	60	64	61
rect	63	61	64	62
rect	63	62	64	63
rect	63	63	64	64
rect	63	64	64	65
rect	63	65	64	66
rect	63	66	64	67
rect	63	67	64	68
rect	63	68	64	69
rect	63	69	64	70
rect	63	70	64	71
rect	63	71	64	72
rect	63	72	64	73
rect	63	73	64	74
rect	63	74	64	75
rect	63	75	64	76
rect	63	76	64	77
rect	63	77	64	78
rect	63	78	64	79
rect	63	79	64	80
rect	63	80	64	81
rect	63	81	64	82
rect	63	82	64	83
rect	63	83	64	84
rect	63	84	64	85
rect	63	85	64	86
rect	63	86	64	87
rect	63	87	64	88
rect	63	88	64	89
rect	63	89	64	90
rect	63	90	64	91
rect	63	91	64	92
rect	63	92	64	93
rect	64	0	65	1
rect	64	1	65	2
rect	64	2	65	3
rect	64	3	65	4
rect	64	4	65	5
rect	64	5	65	6
rect	64	6	65	7
rect	64	7	65	8
rect	64	8	65	9
rect	64	9	65	10
rect	64	10	65	11
rect	64	11	65	12
rect	64	12	65	13
rect	64	13	65	14
rect	64	14	65	15
rect	64	15	65	16
rect	64	16	65	17
rect	64	17	65	18
rect	64	18	65	19
rect	64	19	65	20
rect	64	20	65	21
rect	64	21	65	22
rect	64	22	65	23
rect	64	23	65	24
rect	64	24	65	25
rect	64	25	65	26
rect	64	26	65	27
rect	64	27	65	28
rect	64	28	65	29
rect	64	29	65	30
rect	64	30	65	31
rect	64	31	65	32
rect	64	32	65	33
rect	64	33	65	34
rect	64	34	65	35
rect	64	35	65	36
rect	64	36	65	37
rect	64	37	65	38
rect	64	38	65	39
rect	64	39	65	40
rect	64	40	65	41
rect	64	41	65	42
rect	64	42	65	43
rect	64	43	65	44
rect	64	44	65	45
rect	64	45	65	46
rect	64	46	65	47
rect	64	47	65	48
rect	64	48	65	49
rect	64	49	65	50
rect	64	50	65	51
rect	64	51	65	52
rect	64	52	65	53
rect	64	53	65	54
rect	64	54	65	55
rect	64	55	65	56
rect	64	56	65	57
rect	64	57	65	58
rect	64	58	65	59
rect	64	59	65	60
rect	64	60	65	61
rect	64	61	65	62
rect	64	62	65	63
rect	64	63	65	64
rect	64	64	65	65
rect	64	65	65	66
rect	64	66	65	67
rect	64	67	65	68
rect	64	68	65	69
rect	64	69	65	70
rect	64	70	65	71
rect	64	71	65	72
rect	64	72	65	73
rect	64	73	65	74
rect	64	74	65	75
rect	64	75	65	76
rect	64	76	65	77
rect	64	77	65	78
rect	64	78	65	79
rect	64	79	65	80
rect	64	80	65	81
rect	64	81	65	82
rect	64	82	65	83
rect	64	83	65	84
rect	64	84	65	85
rect	64	85	65	86
rect	64	86	65	87
rect	64	87	65	88
rect	64	88	65	89
rect	64	89	65	90
rect	64	90	65	91
rect	64	91	65	92
rect	64	92	65	93
rect	86	0	87	1
rect	86	1	87	2
rect	86	2	87	3
rect	86	3	87	4
rect	86	4	87	5
rect	86	5	87	6
rect	86	6	87	7
rect	86	7	87	8
rect	86	8	87	9
rect	86	9	87	10
rect	86	10	87	11
rect	86	11	87	12
rect	86	12	87	13
rect	86	13	87	14
rect	86	14	87	15
rect	86	15	87	16
rect	86	16	87	17
rect	86	17	87	18
rect	86	18	87	19
rect	86	19	87	20
rect	86	20	87	21
rect	86	21	87	22
rect	86	22	87	23
rect	86	23	87	24
rect	86	24	87	25
rect	86	25	87	26
rect	86	26	87	27
rect	86	27	87	28
rect	86	28	87	29
rect	86	29	87	30
rect	86	30	87	31
rect	86	31	87	32
rect	86	32	87	33
rect	86	33	87	34
rect	86	34	87	35
rect	86	35	87	36
rect	86	36	87	37
rect	86	37	87	38
rect	86	38	87	39
rect	86	39	87	40
rect	86	40	87	41
rect	86	41	87	42
rect	86	42	87	43
rect	86	43	87	44
rect	86	44	87	45
rect	86	45	87	46
rect	86	46	87	47
rect	86	47	87	48
rect	86	48	87	49
rect	86	49	87	50
rect	86	50	87	51
rect	86	51	87	52
rect	86	52	87	53
rect	86	53	87	54
rect	86	54	87	55
rect	86	55	87	56
rect	86	56	87	57
rect	86	57	87	58
rect	86	58	87	59
rect	86	59	87	60
rect	86	60	87	61
rect	86	61	87	62
rect	86	62	87	63
rect	86	63	87	64
rect	86	64	87	65
rect	86	65	87	66
rect	86	66	87	67
rect	86	67	87	68
rect	86	68	87	69
rect	86	69	87	70
rect	86	70	87	71
rect	86	71	87	72
rect	86	72	87	73
rect	86	73	87	74
rect	86	74	87	75
rect	86	75	87	76
rect	86	76	87	77
rect	86	77	87	78
rect	86	78	87	79
rect	86	79	87	80
rect	86	80	87	81
rect	86	81	87	82
rect	86	82	87	83
rect	86	83	87	84
rect	86	84	87	85
rect	86	85	87	86
rect	86	86	87	87
rect	86	87	87	88
rect	86	88	87	89
rect	86	89	87	90
rect	86	90	87	91
rect	86	91	87	92
rect	86	92	87	93
rect	86	93	87	94
rect	86	94	87	95
rect	86	95	87	96
rect	86	96	87	97
rect	86	97	87	98
rect	86	98	87	99
rect	86	99	87	100
rect	86	100	87	101
rect	86	101	87	102
rect	86	102	87	103
rect	86	103	87	104
rect	86	104	87	105
rect	87	0	88	1
rect	87	1	88	2
rect	87	2	88	3
rect	87	3	88	4
rect	87	4	88	5
rect	87	5	88	6
rect	87	6	88	7
rect	87	7	88	8
rect	87	8	88	9
rect	87	9	88	10
rect	87	10	88	11
rect	87	11	88	12
rect	87	12	88	13
rect	87	13	88	14
rect	87	14	88	15
rect	87	15	88	16
rect	87	16	88	17
rect	87	17	88	18
rect	87	18	88	19
rect	87	19	88	20
rect	87	20	88	21
rect	87	21	88	22
rect	87	22	88	23
rect	87	23	88	24
rect	87	24	88	25
rect	87	25	88	26
rect	87	26	88	27
rect	87	27	88	28
rect	87	28	88	29
rect	87	29	88	30
rect	87	30	88	31
rect	87	31	88	32
rect	87	32	88	33
rect	87	33	88	34
rect	87	34	88	35
rect	87	35	88	36
rect	87	36	88	37
rect	87	37	88	38
rect	87	38	88	39
rect	87	39	88	40
rect	87	40	88	41
rect	87	41	88	42
rect	87	42	88	43
rect	87	43	88	44
rect	87	44	88	45
rect	87	45	88	46
rect	87	46	88	47
rect	87	47	88	48
rect	87	48	88	49
rect	87	49	88	50
rect	87	50	88	51
rect	87	51	88	52
rect	87	52	88	53
rect	87	53	88	54
rect	87	54	88	55
rect	87	55	88	56
rect	87	56	88	57
rect	87	57	88	58
rect	87	58	88	59
rect	87	59	88	60
rect	87	60	88	61
rect	87	61	88	62
rect	87	62	88	63
rect	87	63	88	64
rect	87	64	88	65
rect	87	65	88	66
rect	87	66	88	67
rect	87	67	88	68
rect	87	68	88	69
rect	87	69	88	70
rect	87	70	88	71
rect	87	71	88	72
rect	87	72	88	73
rect	87	73	88	74
rect	87	74	88	75
rect	87	75	88	76
rect	87	76	88	77
rect	87	77	88	78
rect	87	78	88	79
rect	87	79	88	80
rect	87	80	88	81
rect	87	81	88	82
rect	87	82	88	83
rect	87	83	88	84
rect	87	84	88	85
rect	87	85	88	86
rect	87	86	88	87
rect	87	87	88	88
rect	87	88	88	89
rect	87	89	88	90
rect	87	90	88	91
rect	87	91	88	92
rect	87	92	88	93
rect	87	93	88	94
rect	87	94	88	95
rect	87	95	88	96
rect	87	96	88	97
rect	87	97	88	98
rect	87	98	88	99
rect	87	99	88	100
rect	87	100	88	101
rect	87	101	88	102
rect	87	102	88	103
rect	87	103	88	104
rect	87	104	88	105
rect	88	0	89	1
rect	88	1	89	2
rect	88	2	89	3
rect	88	3	89	4
rect	88	4	89	5
rect	88	5	89	6
rect	88	6	89	7
rect	88	7	89	8
rect	88	8	89	9
rect	88	9	89	10
rect	88	10	89	11
rect	88	11	89	12
rect	88	12	89	13
rect	88	13	89	14
rect	88	14	89	15
rect	88	15	89	16
rect	88	16	89	17
rect	88	17	89	18
rect	88	18	89	19
rect	88	19	89	20
rect	88	20	89	21
rect	88	21	89	22
rect	88	22	89	23
rect	88	23	89	24
rect	88	24	89	25
rect	88	25	89	26
rect	88	26	89	27
rect	88	27	89	28
rect	88	28	89	29
rect	88	29	89	30
rect	88	30	89	31
rect	88	31	89	32
rect	88	32	89	33
rect	88	33	89	34
rect	88	34	89	35
rect	88	35	89	36
rect	88	36	89	37
rect	88	37	89	38
rect	88	38	89	39
rect	88	39	89	40
rect	88	40	89	41
rect	88	41	89	42
rect	88	42	89	43
rect	88	43	89	44
rect	88	44	89	45
rect	88	45	89	46
rect	88	46	89	47
rect	88	47	89	48
rect	88	48	89	49
rect	88	49	89	50
rect	88	50	89	51
rect	88	51	89	52
rect	88	52	89	53
rect	88	53	89	54
rect	88	54	89	55
rect	88	55	89	56
rect	88	56	89	57
rect	88	57	89	58
rect	88	58	89	59
rect	88	59	89	60
rect	88	60	89	61
rect	88	61	89	62
rect	88	62	89	63
rect	88	63	89	64
rect	88	64	89	65
rect	88	65	89	66
rect	88	66	89	67
rect	88	67	89	68
rect	88	68	89	69
rect	88	69	89	70
rect	88	70	89	71
rect	88	71	89	72
rect	88	72	89	73
rect	88	73	89	74
rect	88	74	89	75
rect	88	75	89	76
rect	88	76	89	77
rect	88	77	89	78
rect	88	78	89	79
rect	88	79	89	80
rect	88	80	89	81
rect	88	81	89	82
rect	88	82	89	83
rect	88	83	89	84
rect	88	84	89	85
rect	88	85	89	86
rect	88	86	89	87
rect	88	87	89	88
rect	88	88	89	89
rect	88	89	89	90
rect	88	90	89	91
rect	88	91	89	92
rect	88	92	89	93
rect	88	93	89	94
rect	88	94	89	95
rect	88	95	89	96
rect	88	96	89	97
rect	88	97	89	98
rect	88	98	89	99
rect	88	99	89	100
rect	88	100	89	101
rect	88	101	89	102
rect	88	102	89	103
rect	88	103	89	104
rect	88	104	89	105
rect	89	0	90	1
rect	89	1	90	2
rect	89	2	90	3
rect	89	3	90	4
rect	89	4	90	5
rect	89	5	90	6
rect	89	6	90	7
rect	89	7	90	8
rect	89	8	90	9
rect	89	9	90	10
rect	89	10	90	11
rect	89	11	90	12
rect	89	12	90	13
rect	89	13	90	14
rect	89	14	90	15
rect	89	15	90	16
rect	89	16	90	17
rect	89	17	90	18
rect	89	18	90	19
rect	89	19	90	20
rect	89	20	90	21
rect	89	21	90	22
rect	89	22	90	23
rect	89	23	90	24
rect	89	24	90	25
rect	89	25	90	26
rect	89	26	90	27
rect	89	27	90	28
rect	89	28	90	29
rect	89	29	90	30
rect	89	30	90	31
rect	89	31	90	32
rect	89	32	90	33
rect	89	33	90	34
rect	89	34	90	35
rect	89	35	90	36
rect	89	36	90	37
rect	89	37	90	38
rect	89	38	90	39
rect	89	39	90	40
rect	89	40	90	41
rect	89	41	90	42
rect	89	42	90	43
rect	89	43	90	44
rect	89	44	90	45
rect	89	45	90	46
rect	89	46	90	47
rect	89	47	90	48
rect	89	48	90	49
rect	89	49	90	50
rect	89	50	90	51
rect	89	51	90	52
rect	89	52	90	53
rect	89	53	90	54
rect	89	54	90	55
rect	89	55	90	56
rect	89	56	90	57
rect	89	57	90	58
rect	89	58	90	59
rect	89	59	90	60
rect	89	60	90	61
rect	89	61	90	62
rect	89	62	90	63
rect	89	63	90	64
rect	89	64	90	65
rect	89	65	90	66
rect	89	66	90	67
rect	89	67	90	68
rect	89	68	90	69
rect	89	69	90	70
rect	89	70	90	71
rect	89	71	90	72
rect	89	72	90	73
rect	89	73	90	74
rect	89	74	90	75
rect	89	75	90	76
rect	89	76	90	77
rect	89	77	90	78
rect	89	78	90	79
rect	89	79	90	80
rect	89	80	90	81
rect	89	81	90	82
rect	89	82	90	83
rect	89	83	90	84
rect	89	84	90	85
rect	89	85	90	86
rect	89	86	90	87
rect	89	87	90	88
rect	89	88	90	89
rect	89	89	90	90
rect	89	90	90	91
rect	89	91	90	92
rect	89	92	90	93
rect	89	93	90	94
rect	89	94	90	95
rect	89	95	90	96
rect	89	96	90	97
rect	89	97	90	98
rect	89	98	90	99
rect	89	99	90	100
rect	89	100	90	101
rect	89	101	90	102
rect	89	102	90	103
rect	89	103	90	104
rect	89	104	90	105
rect	90	0	91	1
rect	90	1	91	2
rect	90	2	91	3
rect	90	3	91	4
rect	90	4	91	5
rect	90	5	91	6
rect	90	6	91	7
rect	90	7	91	8
rect	90	8	91	9
rect	90	9	91	10
rect	90	10	91	11
rect	90	11	91	12
rect	90	12	91	13
rect	90	13	91	14
rect	90	14	91	15
rect	90	15	91	16
rect	90	16	91	17
rect	90	17	91	18
rect	90	18	91	19
rect	90	19	91	20
rect	90	20	91	21
rect	90	21	91	22
rect	90	22	91	23
rect	90	23	91	24
rect	90	24	91	25
rect	90	25	91	26
rect	90	26	91	27
rect	90	27	91	28
rect	90	28	91	29
rect	90	29	91	30
rect	90	30	91	31
rect	90	31	91	32
rect	90	32	91	33
rect	90	33	91	34
rect	90	34	91	35
rect	90	35	91	36
rect	90	36	91	37
rect	90	37	91	38
rect	90	38	91	39
rect	90	39	91	40
rect	90	40	91	41
rect	90	41	91	42
rect	90	42	91	43
rect	90	43	91	44
rect	90	44	91	45
rect	90	45	91	46
rect	90	46	91	47
rect	90	47	91	48
rect	90	48	91	49
rect	90	49	91	50
rect	90	50	91	51
rect	90	51	91	52
rect	90	52	91	53
rect	90	53	91	54
rect	90	54	91	55
rect	90	55	91	56
rect	90	56	91	57
rect	90	57	91	58
rect	90	58	91	59
rect	90	59	91	60
rect	90	60	91	61
rect	90	61	91	62
rect	90	62	91	63
rect	90	63	91	64
rect	90	64	91	65
rect	90	65	91	66
rect	90	66	91	67
rect	90	67	91	68
rect	90	68	91	69
rect	90	69	91	70
rect	90	70	91	71
rect	90	71	91	72
rect	90	72	91	73
rect	90	73	91	74
rect	90	74	91	75
rect	90	75	91	76
rect	90	76	91	77
rect	90	77	91	78
rect	90	78	91	79
rect	90	79	91	80
rect	90	80	91	81
rect	90	81	91	82
rect	90	82	91	83
rect	90	83	91	84
rect	90	84	91	85
rect	90	85	91	86
rect	90	86	91	87
rect	90	87	91	88
rect	90	88	91	89
rect	90	89	91	90
rect	90	90	91	91
rect	90	91	91	92
rect	90	92	91	93
rect	90	93	91	94
rect	90	94	91	95
rect	90	95	91	96
rect	90	96	91	97
rect	90	97	91	98
rect	90	98	91	99
rect	90	99	91	100
rect	90	100	91	101
rect	90	101	91	102
rect	90	102	91	103
rect	90	103	91	104
rect	90	104	91	105
rect	91	0	92	1
rect	91	1	92	2
rect	91	2	92	3
rect	91	3	92	4
rect	91	4	92	5
rect	91	5	92	6
rect	91	6	92	7
rect	91	7	92	8
rect	91	8	92	9
rect	91	9	92	10
rect	91	10	92	11
rect	91	11	92	12
rect	91	12	92	13
rect	91	13	92	14
rect	91	14	92	15
rect	91	15	92	16
rect	91	16	92	17
rect	91	17	92	18
rect	91	18	92	19
rect	91	19	92	20
rect	91	20	92	21
rect	91	21	92	22
rect	91	22	92	23
rect	91	23	92	24
rect	91	24	92	25
rect	91	25	92	26
rect	91	26	92	27
rect	91	27	92	28
rect	91	28	92	29
rect	91	29	92	30
rect	91	30	92	31
rect	91	31	92	32
rect	91	32	92	33
rect	91	33	92	34
rect	91	34	92	35
rect	91	35	92	36
rect	91	36	92	37
rect	91	37	92	38
rect	91	38	92	39
rect	91	39	92	40
rect	91	40	92	41
rect	91	41	92	42
rect	91	42	92	43
rect	91	43	92	44
rect	91	44	92	45
rect	91	45	92	46
rect	91	46	92	47
rect	91	47	92	48
rect	91	48	92	49
rect	91	49	92	50
rect	91	50	92	51
rect	91	51	92	52
rect	91	52	92	53
rect	91	53	92	54
rect	91	54	92	55
rect	91	55	92	56
rect	91	56	92	57
rect	91	57	92	58
rect	91	58	92	59
rect	91	59	92	60
rect	91	60	92	61
rect	91	61	92	62
rect	91	62	92	63
rect	91	63	92	64
rect	91	64	92	65
rect	91	65	92	66
rect	91	66	92	67
rect	91	67	92	68
rect	91	68	92	69
rect	91	69	92	70
rect	91	70	92	71
rect	91	71	92	72
rect	91	72	92	73
rect	91	73	92	74
rect	91	74	92	75
rect	91	75	92	76
rect	91	76	92	77
rect	91	77	92	78
rect	91	78	92	79
rect	91	79	92	80
rect	91	80	92	81
rect	91	81	92	82
rect	91	82	92	83
rect	91	83	92	84
rect	91	84	92	85
rect	91	85	92	86
rect	91	86	92	87
rect	91	87	92	88
rect	91	88	92	89
rect	91	89	92	90
rect	91	90	92	91
rect	91	91	92	92
rect	91	92	92	93
rect	91	93	92	94
rect	91	94	92	95
rect	91	95	92	96
rect	91	96	92	97
rect	91	97	92	98
rect	91	98	92	99
rect	91	99	92	100
rect	91	100	92	101
rect	91	101	92	102
rect	91	102	92	103
rect	91	103	92	104
rect	91	104	92	105
rect	111	0	112	1
rect	111	1	112	2
rect	111	2	112	3
rect	111	3	112	4
rect	111	4	112	5
rect	111	5	112	6
rect	111	6	112	7
rect	111	7	112	8
rect	111	8	112	9
rect	111	9	112	10
rect	111	10	112	11
rect	111	11	112	12
rect	111	12	112	13
rect	111	13	112	14
rect	111	14	112	15
rect	111	15	112	16
rect	111	16	112	17
rect	111	17	112	18
rect	111	18	112	19
rect	111	19	112	20
rect	111	20	112	21
rect	111	21	112	22
rect	111	22	112	23
rect	111	23	112	24
rect	111	24	112	25
rect	111	25	112	26
rect	111	26	112	27
rect	111	27	112	28
rect	111	28	112	29
rect	111	29	112	30
rect	111	30	112	31
rect	111	31	112	32
rect	111	32	112	33
rect	111	33	112	34
rect	111	34	112	35
rect	111	35	112	36
rect	111	36	112	37
rect	111	37	112	38
rect	111	38	112	39
rect	111	39	112	40
rect	111	40	112	41
rect	111	41	112	42
rect	111	42	112	43
rect	111	43	112	44
rect	111	44	112	45
rect	111	45	112	46
rect	111	46	112	47
rect	111	47	112	48
rect	111	48	112	49
rect	111	49	112	50
rect	111	50	112	51
rect	111	51	112	52
rect	111	52	112	53
rect	111	53	112	54
rect	111	54	112	55
rect	111	55	112	56
rect	111	56	112	57
rect	111	57	112	58
rect	111	58	112	59
rect	111	59	112	60
rect	111	60	112	61
rect	111	61	112	62
rect	111	62	112	63
rect	111	63	112	64
rect	111	64	112	65
rect	111	65	112	66
rect	111	66	112	67
rect	111	67	112	68
rect	111	68	112	69
rect	111	69	112	70
rect	111	70	112	71
rect	111	71	112	72
rect	111	72	112	73
rect	111	73	112	74
rect	111	74	112	75
rect	111	75	112	76
rect	111	76	112	77
rect	111	77	112	78
rect	112	0	113	1
rect	112	1	113	2
rect	112	2	113	3
rect	112	3	113	4
rect	112	4	113	5
rect	112	5	113	6
rect	112	6	113	7
rect	112	7	113	8
rect	112	8	113	9
rect	112	9	113	10
rect	112	10	113	11
rect	112	11	113	12
rect	112	12	113	13
rect	112	13	113	14
rect	112	14	113	15
rect	112	15	113	16
rect	112	16	113	17
rect	112	17	113	18
rect	112	18	113	19
rect	112	19	113	20
rect	112	20	113	21
rect	112	21	113	22
rect	112	22	113	23
rect	112	23	113	24
rect	112	24	113	25
rect	112	25	113	26
rect	112	26	113	27
rect	112	27	113	28
rect	112	28	113	29
rect	112	29	113	30
rect	112	30	113	31
rect	112	31	113	32
rect	112	32	113	33
rect	112	33	113	34
rect	112	34	113	35
rect	112	35	113	36
rect	112	36	113	37
rect	112	37	113	38
rect	112	38	113	39
rect	112	39	113	40
rect	112	40	113	41
rect	112	41	113	42
rect	112	42	113	43
rect	112	43	113	44
rect	112	44	113	45
rect	112	45	113	46
rect	112	46	113	47
rect	112	47	113	48
rect	112	48	113	49
rect	112	49	113	50
rect	112	50	113	51
rect	112	51	113	52
rect	112	52	113	53
rect	112	53	113	54
rect	112	54	113	55
rect	112	55	113	56
rect	112	56	113	57
rect	112	57	113	58
rect	112	58	113	59
rect	112	59	113	60
rect	112	60	113	61
rect	112	61	113	62
rect	112	62	113	63
rect	112	63	113	64
rect	112	64	113	65
rect	112	65	113	66
rect	112	66	113	67
rect	112	67	113	68
rect	112	68	113	69
rect	112	69	113	70
rect	112	70	113	71
rect	112	71	113	72
rect	112	72	113	73
rect	112	73	113	74
rect	112	74	113	75
rect	112	75	113	76
rect	112	76	113	77
rect	112	77	113	78
rect	113	0	114	1
rect	113	1	114	2
rect	113	2	114	3
rect	113	3	114	4
rect	113	4	114	5
rect	113	5	114	6
rect	113	6	114	7
rect	113	7	114	8
rect	113	8	114	9
rect	113	9	114	10
rect	113	10	114	11
rect	113	11	114	12
rect	113	12	114	13
rect	113	13	114	14
rect	113	14	114	15
rect	113	15	114	16
rect	113	16	114	17
rect	113	17	114	18
rect	113	18	114	19
rect	113	19	114	20
rect	113	20	114	21
rect	113	21	114	22
rect	113	22	114	23
rect	113	23	114	24
rect	113	24	114	25
rect	113	25	114	26
rect	113	26	114	27
rect	113	27	114	28
rect	113	28	114	29
rect	113	29	114	30
rect	113	30	114	31
rect	113	31	114	32
rect	113	32	114	33
rect	113	33	114	34
rect	113	34	114	35
rect	113	35	114	36
rect	113	36	114	37
rect	113	37	114	38
rect	113	38	114	39
rect	113	39	114	40
rect	113	40	114	41
rect	113	41	114	42
rect	113	42	114	43
rect	113	43	114	44
rect	113	44	114	45
rect	113	45	114	46
rect	113	46	114	47
rect	113	47	114	48
rect	113	48	114	49
rect	113	49	114	50
rect	113	50	114	51
rect	113	51	114	52
rect	113	52	114	53
rect	113	53	114	54
rect	113	54	114	55
rect	113	55	114	56
rect	113	56	114	57
rect	113	57	114	58
rect	113	58	114	59
rect	113	59	114	60
rect	113	60	114	61
rect	113	61	114	62
rect	113	62	114	63
rect	113	63	114	64
rect	113	64	114	65
rect	113	65	114	66
rect	113	66	114	67
rect	113	67	114	68
rect	113	68	114	69
rect	113	69	114	70
rect	113	70	114	71
rect	113	71	114	72
rect	113	72	114	73
rect	113	73	114	74
rect	113	74	114	75
rect	113	75	114	76
rect	113	76	114	77
rect	113	77	114	78
rect	114	0	115	1
rect	114	1	115	2
rect	114	2	115	3
rect	114	3	115	4
rect	114	4	115	5
rect	114	5	115	6
rect	114	6	115	7
rect	114	7	115	8
rect	114	8	115	9
rect	114	9	115	10
rect	114	10	115	11
rect	114	11	115	12
rect	114	12	115	13
rect	114	13	115	14
rect	114	14	115	15
rect	114	15	115	16
rect	114	16	115	17
rect	114	17	115	18
rect	114	18	115	19
rect	114	19	115	20
rect	114	20	115	21
rect	114	21	115	22
rect	114	22	115	23
rect	114	23	115	24
rect	114	24	115	25
rect	114	25	115	26
rect	114	26	115	27
rect	114	27	115	28
rect	114	28	115	29
rect	114	29	115	30
rect	114	30	115	31
rect	114	31	115	32
rect	114	32	115	33
rect	114	33	115	34
rect	114	34	115	35
rect	114	35	115	36
rect	114	36	115	37
rect	114	37	115	38
rect	114	38	115	39
rect	114	39	115	40
rect	114	40	115	41
rect	114	41	115	42
rect	114	42	115	43
rect	114	43	115	44
rect	114	44	115	45
rect	114	45	115	46
rect	114	46	115	47
rect	114	47	115	48
rect	114	48	115	49
rect	114	49	115	50
rect	114	50	115	51
rect	114	51	115	52
rect	114	52	115	53
rect	114	53	115	54
rect	114	54	115	55
rect	114	55	115	56
rect	114	56	115	57
rect	114	57	115	58
rect	114	58	115	59
rect	114	59	115	60
rect	114	60	115	61
rect	114	61	115	62
rect	114	62	115	63
rect	114	63	115	64
rect	114	64	115	65
rect	114	65	115	66
rect	114	66	115	67
rect	114	67	115	68
rect	114	68	115	69
rect	114	69	115	70
rect	114	70	115	71
rect	114	71	115	72
rect	114	72	115	73
rect	114	73	115	74
rect	114	74	115	75
rect	114	75	115	76
rect	114	76	115	77
rect	114	77	115	78
rect	115	0	116	1
rect	115	1	116	2
rect	115	2	116	3
rect	115	3	116	4
rect	115	4	116	5
rect	115	5	116	6
rect	115	6	116	7
rect	115	7	116	8
rect	115	8	116	9
rect	115	9	116	10
rect	115	10	116	11
rect	115	11	116	12
rect	115	12	116	13
rect	115	13	116	14
rect	115	14	116	15
rect	115	15	116	16
rect	115	16	116	17
rect	115	17	116	18
rect	115	18	116	19
rect	115	19	116	20
rect	115	20	116	21
rect	115	21	116	22
rect	115	22	116	23
rect	115	23	116	24
rect	115	24	116	25
rect	115	25	116	26
rect	115	26	116	27
rect	115	27	116	28
rect	115	28	116	29
rect	115	29	116	30
rect	115	30	116	31
rect	115	31	116	32
rect	115	32	116	33
rect	115	33	116	34
rect	115	34	116	35
rect	115	35	116	36
rect	115	36	116	37
rect	115	37	116	38
rect	115	38	116	39
rect	115	39	116	40
rect	115	40	116	41
rect	115	41	116	42
rect	115	42	116	43
rect	115	43	116	44
rect	115	44	116	45
rect	115	45	116	46
rect	115	46	116	47
rect	115	47	116	48
rect	115	48	116	49
rect	115	49	116	50
rect	115	50	116	51
rect	115	51	116	52
rect	115	52	116	53
rect	115	53	116	54
rect	115	54	116	55
rect	115	55	116	56
rect	115	56	116	57
rect	115	57	116	58
rect	115	58	116	59
rect	115	59	116	60
rect	115	60	116	61
rect	115	61	116	62
rect	115	62	116	63
rect	115	63	116	64
rect	115	64	116	65
rect	115	65	116	66
rect	115	66	116	67
rect	115	67	116	68
rect	115	68	116	69
rect	115	69	116	70
rect	115	70	116	71
rect	115	71	116	72
rect	115	72	116	73
rect	115	73	116	74
rect	115	74	116	75
rect	115	75	116	76
rect	115	76	116	77
rect	115	77	116	78
rect	116	0	117	1
rect	116	1	117	2
rect	116	2	117	3
rect	116	3	117	4
rect	116	4	117	5
rect	116	5	117	6
rect	116	6	117	7
rect	116	7	117	8
rect	116	8	117	9
rect	116	9	117	10
rect	116	10	117	11
rect	116	11	117	12
rect	116	12	117	13
rect	116	13	117	14
rect	116	14	117	15
rect	116	15	117	16
rect	116	16	117	17
rect	116	17	117	18
rect	116	18	117	19
rect	116	19	117	20
rect	116	20	117	21
rect	116	21	117	22
rect	116	22	117	23
rect	116	23	117	24
rect	116	24	117	25
rect	116	25	117	26
rect	116	26	117	27
rect	116	27	117	28
rect	116	28	117	29
rect	116	29	117	30
rect	116	30	117	31
rect	116	31	117	32
rect	116	32	117	33
rect	116	33	117	34
rect	116	34	117	35
rect	116	35	117	36
rect	116	36	117	37
rect	116	37	117	38
rect	116	38	117	39
rect	116	39	117	40
rect	116	40	117	41
rect	116	41	117	42
rect	116	42	117	43
rect	116	43	117	44
rect	116	44	117	45
rect	116	45	117	46
rect	116	46	117	47
rect	116	47	117	48
rect	116	48	117	49
rect	116	49	117	50
rect	116	50	117	51
rect	116	51	117	52
rect	116	52	117	53
rect	116	53	117	54
rect	116	54	117	55
rect	116	55	117	56
rect	116	56	117	57
rect	116	57	117	58
rect	116	58	117	59
rect	116	59	117	60
rect	116	60	117	61
rect	116	61	117	62
rect	116	62	117	63
rect	116	63	117	64
rect	116	64	117	65
rect	116	65	117	66
rect	116	66	117	67
rect	116	67	117	68
rect	116	68	117	69
rect	116	69	117	70
rect	116	70	117	71
rect	116	71	117	72
rect	116	72	117	73
rect	116	73	117	74
rect	116	74	117	75
rect	116	75	117	76
rect	116	76	117	77
rect	116	77	117	78
rect	132	0	133	1
rect	132	1	133	2
rect	132	2	133	3
rect	132	3	133	4
rect	132	4	133	5
rect	132	5	133	6
rect	132	6	133	7
rect	132	7	133	8
rect	132	8	133	9
rect	132	9	133	10
rect	132	10	133	11
rect	132	11	133	12
rect	132	12	133	13
rect	132	13	133	14
rect	132	14	133	15
rect	132	15	133	16
rect	132	16	133	17
rect	132	17	133	18
rect	132	18	133	19
rect	132	19	133	20
rect	132	20	133	21
rect	132	21	133	22
rect	132	22	133	23
rect	132	23	133	24
rect	132	24	133	25
rect	132	25	133	26
rect	132	26	133	27
rect	133	0	134	1
rect	133	1	134	2
rect	133	2	134	3
rect	133	3	134	4
rect	133	4	134	5
rect	133	5	134	6
rect	133	6	134	7
rect	133	7	134	8
rect	133	8	134	9
rect	133	9	134	10
rect	133	10	134	11
rect	133	11	134	12
rect	133	12	134	13
rect	133	13	134	14
rect	133	14	134	15
rect	133	15	134	16
rect	133	16	134	17
rect	133	17	134	18
rect	133	18	134	19
rect	133	19	134	20
rect	133	20	134	21
rect	133	21	134	22
rect	133	22	134	23
rect	133	23	134	24
rect	133	24	134	25
rect	133	25	134	26
rect	133	26	134	27
rect	134	0	135	1
rect	134	1	135	2
rect	134	2	135	3
rect	134	3	135	4
rect	134	4	135	5
rect	134	5	135	6
rect	134	6	135	7
rect	134	7	135	8
rect	134	8	135	9
rect	134	9	135	10
rect	134	10	135	11
rect	134	11	135	12
rect	134	12	135	13
rect	134	13	135	14
rect	134	14	135	15
rect	134	15	135	16
rect	134	16	135	17
rect	134	17	135	18
rect	134	18	135	19
rect	134	19	135	20
rect	134	20	135	21
rect	134	21	135	22
rect	134	22	135	23
rect	134	23	135	24
rect	134	24	135	25
rect	134	25	135	26
rect	134	26	135	27
rect	135	0	136	1
rect	135	1	136	2
rect	135	2	136	3
rect	135	3	136	4
rect	135	4	136	5
rect	135	5	136	6
rect	135	6	136	7
rect	135	7	136	8
rect	135	8	136	9
rect	135	9	136	10
rect	135	10	136	11
rect	135	11	136	12
rect	135	12	136	13
rect	135	13	136	14
rect	135	14	136	15
rect	135	15	136	16
rect	135	16	136	17
rect	135	17	136	18
rect	135	18	136	19
rect	135	19	136	20
rect	135	20	136	21
rect	135	21	136	22
rect	135	22	136	23
rect	135	23	136	24
rect	135	24	136	25
rect	135	25	136	26
rect	135	26	136	27
rect	136	0	137	1
rect	136	1	137	2
rect	136	2	137	3
rect	136	3	137	4
rect	136	4	137	5
rect	136	5	137	6
rect	136	6	137	7
rect	136	7	137	8
rect	136	8	137	9
rect	136	9	137	10
rect	136	10	137	11
rect	136	11	137	12
rect	136	12	137	13
rect	136	13	137	14
rect	136	14	137	15
rect	136	15	137	16
rect	136	16	137	17
rect	136	17	137	18
rect	136	18	137	19
rect	136	19	137	20
rect	136	20	137	21
rect	136	21	137	22
rect	136	22	137	23
rect	136	23	137	24
rect	136	24	137	25
rect	136	25	137	26
rect	136	26	137	27
rect	137	0	138	1
rect	137	1	138	2
rect	137	2	138	3
rect	137	3	138	4
rect	137	4	138	5
rect	137	5	138	6
rect	137	6	138	7
rect	137	7	138	8
rect	137	8	138	9
rect	137	9	138	10
rect	137	10	138	11
rect	137	11	138	12
rect	137	12	138	13
rect	137	13	138	14
rect	137	14	138	15
rect	137	15	138	16
rect	137	16	138	17
rect	137	17	138	18
rect	137	18	138	19
rect	137	19	138	20
rect	137	20	138	21
rect	137	21	138	22
rect	137	22	138	23
rect	137	23	138	24
rect	137	24	138	25
rect	137	25	138	26
rect	137	26	138	27
<< metal1 >>
rect	0	5	1	6
rect	0	6	1	7
rect	0	7	1	8
rect	0	8	1	9
rect	0	9	1	10
rect	0	10	1	11
rect	0	11	1	12
rect	0	12	1	13
rect	0	13	1	14
rect	0	14	1	15
rect	0	15	1	16
rect	0	16	1	17
rect	0	17	1	18
rect	0	18	1	19
rect	0	19	1	20
rect	0	20	1	21
rect	0	21	1	22
rect	0	22	1	23
rect	0	23	1	24
rect	0	24	1	25
rect	0	25	1	26
rect	0	26	1	27
rect	0	27	1	28
rect	0	28	1	29
rect	0	29	1	30
rect	0	30	1	31
rect	0	31	1	32
rect	0	32	1	33
rect	0	33	1	34
rect	0	34	1	35
rect	0	35	1	36
rect	0	36	1	37
rect	0	37	1	38
rect	0	38	1	39
rect	0	39	1	40
rect	0	40	1	41
rect	0	41	1	42
rect	0	42	1	43
rect	0	43	1	44
rect	0	44	1	45
rect	0	45	1	46
rect	0	46	1	47
rect	0	47	1	48
rect	0	48	1	49
rect	2	2	3	3
rect	2	3	3	4
rect	2	5	3	6
rect	2	6	3	7
rect	2	11	3	12
rect	2	12	3	13
rect	2	17	3	18
rect	2	18	3	19
rect	2	47	3	48
rect	2	48	3	49
rect	2	50	3	51
rect	2	51	3	52
rect	11	26	12	27
rect	11	27	12	28
rect	11	28	12	29
rect	11	29	12	30
rect	11	30	12	31
rect	11	47	12	48
rect	11	48	12	49
rect	11	50	12	51
rect	11	51	12	52
rect	11	53	12	54
rect	11	54	12	55
rect	11	55	12	56
rect	11	56	12	57
rect	11	57	12	58
rect	11	58	12	59
rect	11	59	12	60
rect	11	60	12	61
rect	11	61	12	62
rect	11	62	12	63
rect	11	63	12	64
rect	11	64	12	65
rect	11	65	12	66
rect	11	66	12	67
rect	13	20	14	21
rect	13	21	14	22
rect	13	22	14	23
rect	13	23	14	24
rect	13	24	14	25
rect	13	26	14	27
rect	13	27	14	28
rect	13	38	14	39
rect	13	39	14	40
rect	13	40	14	41
rect	13	41	14	42
rect	13	42	14	43
rect	13	43	14	44
rect	13	44	14	45
rect	13	45	14	46
rect	15	14	16	15
rect	15	15	16	16
rect	15	16	16	17
rect	15	17	16	18
rect	15	18	16	19
rect	15	19	16	20
rect	15	20	16	21
rect	15	21	16	22
rect	15	22	16	23
rect	15	23	16	24
rect	15	24	16	25
rect	15	26	16	27
rect	15	27	16	28
rect	15	29	16	30
rect	15	30	16	31
rect	15	31	16	32
rect	15	32	16	33
rect	15	33	16	34
rect	15	34	16	35
rect	15	35	16	36
rect	15	36	16	37
rect	15	38	16	39
rect	15	39	16	40
rect	15	40	16	41
rect	15	41	16	42
rect	15	42	16	43
rect	15	43	16	44
rect	15	44	16	45
rect	15	45	16	46
rect	15	47	16	48
rect	15	48	16	49
rect	15	50	16	51
rect	15	51	16	52
rect	15	53	16	54
rect	15	54	16	55
rect	15	55	16	56
rect	15	56	16	57
rect	15	57	16	58
rect	15	58	16	59
rect	15	59	16	60
rect	15	60	16	61
rect	17	11	18	12
rect	17	12	18	13
rect	17	14	18	15
rect	17	15	18	16
rect	17	20	18	21
rect	17	21	18	22
rect	17	22	18	23
rect	17	23	18	24
rect	17	24	18	25
rect	17	26	18	27
rect	17	27	18	28
rect	17	29	18	30
rect	17	30	18	31
rect	17	31	18	32
rect	17	32	18	33
rect	17	33	18	34
rect	17	34	18	35
rect	17	35	18	36
rect	17	36	18	37
rect	17	38	18	39
rect	17	39	18	40
rect	17	59	18	60
rect	17	60	18	61
rect	17	62	18	63
rect	17	63	18	64
rect	17	64	18	65
rect	17	65	18	66
rect	17	66	18	67
rect	17	68	18	69
rect	17	69	18	70
rect	17	70	18	71
rect	17	71	18	72
rect	17	72	18	73
rect	19	2	20	3
rect	19	3	20	4
rect	19	4	20	5
rect	19	5	20	6
rect	19	6	20	7
rect	19	11	20	12
rect	19	12	20	13
rect	19	14	20	15
rect	19	15	20	16
rect	19	17	20	18
rect	19	18	20	19
rect	19	20	20	21
rect	19	21	20	22
rect	19	22	20	23
rect	19	23	20	24
rect	19	24	20	25
rect	19	26	20	27
rect	19	27	20	28
rect	19	29	20	30
rect	19	30	20	31
rect	19	31	20	32
rect	19	32	20	33
rect	19	33	20	34
rect	19	34	20	35
rect	19	35	20	36
rect	19	36	20	37
rect	19	38	20	39
rect	19	39	20	40
rect	19	41	20	42
rect	19	42	20	43
rect	19	43	20	44
rect	19	44	20	45
rect	19	45	20	46
rect	19	47	20	48
rect	19	48	20	49
rect	19	50	20	51
rect	19	51	20	52
rect	19	56	20	57
rect	19	57	20	58
rect	19	59	20	60
rect	19	60	20	61
rect	19	62	20	63
rect	19	63	20	64
rect	28	65	29	66
rect	28	66	29	67
rect	28	68	29	69
rect	28	69	29	70
rect	28	71	29	72
rect	28	72	29	73
rect	30	20	31	21
rect	30	21	31	22
rect	30	22	31	23
rect	30	23	31	24
rect	30	24	31	25
rect	30	26	31	27
rect	30	27	31	28
rect	30	29	31	30
rect	30	30	31	31
rect	30	31	31	32
rect	30	32	31	33
rect	30	33	31	34
rect	30	34	31	35
rect	30	35	31	36
rect	30	36	31	37
rect	30	50	31	51
rect	30	51	31	52
rect	30	52	31	53
rect	30	53	31	54
rect	30	54	31	55
rect	30	62	31	63
rect	30	63	31	64
rect	30	64	31	65
rect	30	65	31	66
rect	30	66	31	67
rect	30	68	31	69
rect	30	69	31	70
rect	30	71	31	72
rect	30	72	31	73
rect	30	74	31	75
rect	30	75	31	76
rect	30	76	31	77
rect	30	77	31	78
rect	30	78	31	79
rect	32	14	33	15
rect	32	15	33	16
rect	32	17	33	18
rect	32	18	33	19
rect	32	19	33	20
rect	32	20	33	21
rect	32	21	33	22
rect	32	44	33	45
rect	32	45	33	46
rect	32	47	33	48
rect	32	48	33	49
rect	32	49	33	50
rect	32	50	33	51
rect	32	51	33	52
rect	32	52	33	53
rect	32	53	33	54
rect	32	54	33	55
rect	32	56	33	57
rect	32	57	33	58
rect	32	59	33	60
rect	32	60	33	61
rect	32	61	33	62
rect	32	62	33	63
rect	32	63	33	64
rect	32	68	33	69
rect	32	69	33	70
rect	32	71	33	72
rect	32	72	33	73
rect	32	74	33	75
rect	32	75	33	76
rect	34	2	35	3
rect	34	3	35	4
rect	34	4	35	5
rect	34	5	35	6
rect	34	6	35	7
rect	34	14	35	15
rect	34	15	35	16
rect	34	17	35	18
rect	34	18	35	19
rect	34	19	35	20
rect	34	20	35	21
rect	34	21	35	22
rect	34	23	35	24
rect	34	24	35	25
rect	34	26	35	27
rect	34	27	35	28
rect	34	29	35	30
rect	34	30	35	31
rect	34	31	35	32
rect	34	32	35	33
rect	34	33	35	34
rect	34	34	35	35
rect	34	35	35	36
rect	34	36	35	37
rect	34	37	35	38
rect	34	38	35	39
rect	34	39	35	40
rect	34	41	35	42
rect	34	42	35	43
rect	34	43	35	44
rect	34	44	35	45
rect	34	45	35	46
rect	34	47	35	48
rect	34	48	35	49
rect	34	49	35	50
rect	34	50	35	51
rect	34	51	35	52
rect	34	52	35	53
rect	34	53	35	54
rect	34	54	35	55
rect	34	56	35	57
rect	34	57	35	58
rect	34	59	35	60
rect	34	60	35	61
rect	34	61	35	62
rect	34	62	35	63
rect	34	63	35	64
rect	34	65	35	66
rect	34	66	35	67
rect	34	67	35	68
rect	34	68	35	69
rect	34	69	35	70
rect	34	71	35	72
rect	34	72	35	73
rect	34	74	35	75
rect	34	75	35	76
rect	34	77	35	78
rect	34	78	35	79
rect	34	80	35	81
rect	34	81	35	82
rect	34	82	35	83
rect	34	83	35	84
rect	34	84	35	85
rect	36	2	37	3
rect	36	3	37	4
rect	36	4	37	5
rect	36	5	37	6
rect	36	6	37	7
rect	36	11	37	12
rect	36	12	37	13
rect	36	14	37	15
rect	36	15	37	16
rect	36	20	37	21
rect	36	21	37	22
rect	36	23	37	24
rect	36	24	37	25
rect	36	26	37	27
rect	36	27	37	28
rect	36	29	37	30
rect	36	30	37	31
rect	36	41	37	42
rect	36	42	37	43
rect	36	47	37	48
rect	36	48	37	49
rect	36	49	37	50
rect	36	50	37	51
rect	36	51	37	52
rect	36	62	37	63
rect	36	63	37	64
rect	36	65	37	66
rect	36	66	37	67
rect	45	59	46	60
rect	45	60	46	61
rect	47	29	48	30
rect	47	30	48	31
rect	47	32	48	33
rect	47	33	48	34
rect	47	34	48	35
rect	47	35	48	36
rect	47	36	48	37
rect	47	38	48	39
rect	47	39	48	40
rect	47	56	48	57
rect	47	57	48	58
rect	47	58	48	59
rect	47	59	48	60
rect	47	60	48	61
rect	47	61	48	62
rect	47	62	48	63
rect	47	63	48	64
rect	49	29	50	30
rect	49	30	50	31
rect	49	38	50	39
rect	49	39	50	40
rect	49	41	50	42
rect	49	42	50	43
rect	49	44	50	45
rect	49	45	50	46
rect	49	47	50	48
rect	49	48	50	49
rect	49	49	50	50
rect	49	50	50	51
rect	49	51	50	52
rect	49	53	50	54
rect	49	54	50	55
rect	49	55	50	56
rect	49	56	50	57
rect	49	57	50	58
rect	49	68	50	69
rect	49	69	50	70
rect	49	71	50	72
rect	49	72	50	73
rect	49	74	50	75
rect	49	75	50	76
rect	49	77	50	78
rect	49	78	50	79
rect	51	23	52	24
rect	51	24	52	25
rect	51	26	52	27
rect	51	27	52	28
rect	51	29	52	30
rect	51	30	52	31
rect	51	31	52	32
rect	51	32	52	33
rect	51	33	52	34
rect	51	34	52	35
rect	51	35	52	36
rect	51	36	52	37
rect	51	53	52	54
rect	51	54	52	55
rect	51	77	52	78
rect	51	78	52	79
rect	53	5	54	6
rect	53	6	54	7
rect	53	11	54	12
rect	53	12	54	13
rect	53	17	54	18
rect	53	18	54	19
rect	53	20	54	21
rect	53	21	54	22
rect	53	22	54	23
rect	53	23	54	24
rect	53	24	54	25
rect	53	26	54	27
rect	53	27	54	28
rect	53	29	54	30
rect	53	30	54	31
rect	53	31	54	32
rect	53	32	54	33
rect	53	33	54	34
rect	53	34	54	35
rect	53	35	54	36
rect	53	36	54	37
rect	53	38	54	39
rect	53	39	54	40
rect	53	41	54	42
rect	53	42	54	43
rect	53	44	54	45
rect	53	45	54	46
rect	53	47	54	48
rect	53	48	54	49
rect	53	49	54	50
rect	53	50	54	51
rect	53	51	54	52
rect	53	71	54	72
rect	53	72	54	73
rect	53	74	54	75
rect	53	75	54	76
rect	55	2	56	3
rect	55	3	56	4
rect	55	4	56	5
rect	55	5	56	6
rect	55	6	56	7
rect	55	7	56	8
rect	55	8	56	9
rect	55	9	56	10
rect	55	17	56	18
rect	55	18	56	19
rect	55	23	56	24
rect	55	24	56	25
rect	55	26	56	27
rect	55	27	56	28
rect	55	29	56	30
rect	55	30	56	31
rect	55	44	56	45
rect	55	45	56	46
rect	55	71	56	72
rect	55	72	56	73
rect	57	2	58	3
rect	57	3	58	4
rect	57	4	58	5
rect	57	5	58	6
rect	57	6	58	7
rect	57	20	58	21
rect	57	21	58	22
rect	57	23	58	24
rect	57	24	58	25
rect	57	35	58	36
rect	57	36	58	37
rect	57	38	58	39
rect	57	39	58	40
rect	57	41	58	42
rect	57	42	58	43
rect	57	47	58	48
rect	57	48	58	49
rect	57	62	58	63
rect	57	63	58	64
rect	57	74	58	75
rect	57	75	58	76
rect	57	77	58	78
rect	57	78	58	79
rect	57	80	58	81
rect	57	81	58	82
rect	57	86	58	87
rect	57	87	58	88
rect	66	77	67	78
rect	66	78	67	79
rect	66	80	67	81
rect	66	81	67	82
rect	66	83	67	84
rect	66	84	67	85
rect	68	65	69	66
rect	68	66	69	67
rect	68	67	69	68
rect	68	68	69	69
rect	68	69	69	70
rect	68	71	69	72
rect	68	72	69	73
rect	68	74	69	75
rect	68	75	69	76
rect	68	76	69	77
rect	68	77	69	78
rect	68	78	69	79
rect	68	80	69	81
rect	68	81	69	82
rect	68	83	69	84
rect	68	84	69	85
rect	70	62	71	63
rect	70	63	71	64
rect	70	64	71	65
rect	70	65	71	66
rect	70	66	71	67
rect	70	67	71	68
rect	70	68	71	69
rect	70	69	71	70
rect	70	71	71	72
rect	70	72	71	73
rect	72	2	73	3
rect	72	3	73	4
rect	72	14	73	15
rect	72	15	73	16
rect	72	17	73	18
rect	72	18	73	19
rect	72	20	73	21
rect	72	21	73	22
rect	72	22	73	23
rect	72	23	73	24
rect	72	24	73	25
rect	72	56	73	57
rect	72	57	73	58
rect	72	58	73	59
rect	72	59	73	60
rect	72	60	73	61
rect	72	62	73	63
rect	72	63	73	64
rect	74	5	75	6
rect	74	6	75	7
rect	74	7	75	8
rect	74	8	75	9
rect	74	9	75	10
rect	74	11	75	12
rect	74	12	75	13
rect	74	13	75	14
rect	74	14	75	15
rect	74	15	75	16
rect	74	17	75	18
rect	74	18	75	19
rect	74	47	75	48
rect	74	48	75	49
rect	74	50	75	51
rect	74	51	75	52
rect	74	53	75	54
rect	74	54	75	55
rect	74	55	75	56
rect	74	56	75	57
rect	74	57	75	58
rect	74	58	75	59
rect	74	59	75	60
rect	74	60	75	61
rect	74	62	75	63
rect	74	63	75	64
rect	74	65	75	66
rect	74	66	75	67
rect	74	67	75	68
rect	74	68	75	69
rect	74	69	75	70
rect	74	71	75	72
rect	74	72	75	73
rect	76	14	77	15
rect	76	15	77	16
rect	76	17	77	18
rect	76	18	77	19
rect	76	47	77	48
rect	76	48	77	49
rect	76	53	77	54
rect	76	54	77	55
rect	76	77	77	78
rect	76	78	77	79
rect	76	80	77	81
rect	76	81	77	82
rect	78	11	79	12
rect	78	12	79	13
rect	78	14	79	15
rect	78	15	79	16
rect	78	17	79	18
rect	78	18	79	19
rect	78	20	79	21
rect	78	21	79	22
rect	78	44	79	45
rect	78	45	79	46
rect	78	47	79	48
rect	78	48	79	49
rect	78	49	79	50
rect	78	50	79	51
rect	78	51	79	52
rect	78	71	79	72
rect	78	72	79	73
rect	78	74	79	75
rect	78	75	79	76
rect	78	77	79	78
rect	78	78	79	79
rect	78	83	79	84
rect	78	84	79	85
rect	78	86	79	87
rect	78	87	79	88
rect	80	11	81	12
rect	80	12	81	13
rect	80	14	81	15
rect	80	15	81	16
rect	80	17	81	18
rect	80	18	81	19
rect	80	20	81	21
rect	80	21	81	22
rect	80	23	81	24
rect	80	24	81	25
rect	80	25	81	26
rect	80	26	81	27
rect	80	27	81	28
rect	80	29	81	30
rect	80	30	81	31
rect	80	32	81	33
rect	80	33	81	34
rect	80	35	81	36
rect	80	36	81	37
rect	80	38	81	39
rect	80	39	81	40
rect	80	41	81	42
rect	80	42	81	43
rect	80	44	81	45
rect	80	45	81	46
rect	80	47	81	48
rect	80	48	81	49
rect	80	49	81	50
rect	80	50	81	51
rect	80	51	81	52
rect	80	53	81	54
rect	80	54	81	55
rect	80	56	81	57
rect	80	57	81	58
rect	80	58	81	59
rect	80	59	81	60
rect	80	60	81	61
rect	80	62	81	63
rect	80	63	81	64
rect	80	65	81	66
rect	80	66	81	67
rect	80	67	81	68
rect	80	68	81	69
rect	80	69	81	70
rect	80	70	81	71
rect	80	71	81	72
rect	80	72	81	73
rect	80	74	81	75
rect	80	75	81	76
rect	80	77	81	78
rect	80	78	81	79
rect	80	79	81	80
rect	80	80	81	81
rect	80	81	81	82
rect	80	83	81	84
rect	80	84	81	85
rect	80	86	81	87
rect	80	87	81	88
rect	80	89	81	90
rect	80	90	81	91
rect	80	92	81	93
rect	80	93	81	94
rect	82	8	83	9
rect	82	9	83	10
rect	82	11	83	12
rect	82	12	83	13
rect	82	14	83	15
rect	82	15	83	16
rect	82	26	83	27
rect	82	27	83	28
rect	82	38	83	39
rect	82	39	83	40
rect	82	41	83	42
rect	82	42	83	43
rect	82	44	83	45
rect	82	45	83	46
rect	82	47	83	48
rect	82	48	83	49
rect	82	49	83	50
rect	82	50	83	51
rect	82	51	83	52
rect	82	53	83	54
rect	82	54	83	55
rect	82	56	83	57
rect	82	57	83	58
rect	82	58	83	59
rect	82	59	83	60
rect	82	60	83	61
rect	82	62	83	63
rect	82	63	83	64
rect	82	65	83	66
rect	82	66	83	67
rect	82	67	83	68
rect	82	68	83	69
rect	82	69	83	70
rect	82	70	83	71
rect	82	71	83	72
rect	82	72	83	73
rect	82	74	83	75
rect	82	75	83	76
rect	82	77	83	78
rect	82	78	83	79
rect	82	79	83	80
rect	82	80	83	81
rect	82	81	83	82
rect	82	83	83	84
rect	82	84	83	85
rect	82	86	83	87
rect	82	87	83	88
rect	82	89	83	90
rect	82	90	83	91
rect	84	2	85	3
rect	84	3	85	4
rect	84	5	85	6
rect	84	6	85	7
rect	84	8	85	9
rect	84	9	85	10
rect	84	11	85	12
rect	84	12	85	13
rect	84	14	85	15
rect	84	15	85	16
rect	84	29	85	30
rect	84	30	85	31
rect	84	32	85	33
rect	84	33	85	34
rect	84	35	85	36
rect	84	36	85	37
rect	84	41	85	42
rect	84	42	85	43
rect	84	44	85	45
rect	84	45	85	46
rect	84	47	85	48
rect	84	48	85	49
rect	84	59	85	60
rect	84	60	85	61
rect	84	62	85	63
rect	84	63	85	64
rect	84	65	85	66
rect	84	66	85	67
rect	84	80	85	81
rect	84	81	85	82
rect	84	83	85	84
rect	84	84	85	85
rect	84	86	85	87
rect	84	87	85	88
rect	84	89	85	90
rect	84	90	85	91
rect	84	98	85	99
rect	84	99	85	100
rect	84	100	85	101
rect	84	101	85	102
rect	84	102	85	103
rect	93	14	94	15
rect	93	15	94	16
rect	93	17	94	18
rect	93	18	94	19
rect	93	20	94	21
rect	93	21	94	22
rect	93	23	94	24
rect	93	24	94	25
rect	93	26	94	27
rect	93	27	94	28
rect	93	29	94	30
rect	93	30	94	31
rect	93	32	94	33
rect	93	33	94	34
rect	95	32	96	33
rect	95	33	96	34
rect	97	32	98	33
rect	97	33	98	34
rect	97	35	98	36
rect	97	36	98	37
rect	97	38	98	39
rect	97	39	98	40
rect	97	41	98	42
rect	97	42	98	43
rect	99	20	100	21
rect	99	21	100	22
rect	99	23	100	24
rect	99	24	100	25
rect	99	26	100	27
rect	99	27	100	28
rect	99	29	100	30
rect	99	30	100	31
rect	99	32	100	33
rect	99	33	100	34
rect	99	35	100	36
rect	99	36	100	37
rect	99	62	100	63
rect	99	63	100	64
rect	99	65	100	66
rect	99	66	100	67
rect	99	68	100	69
rect	99	69	100	70
rect	101	17	102	18
rect	101	18	102	19
rect	101	19	102	20
rect	101	20	102	21
rect	101	21	102	22
rect	101	23	102	24
rect	101	24	102	25
rect	101	26	102	27
rect	101	27	102	28
rect	101	29	102	30
rect	101	30	102	31
rect	101	32	102	33
rect	101	33	102	34
rect	101	35	102	36
rect	101	36	102	37
rect	101	37	102	38
rect	101	38	102	39
rect	101	39	102	40
rect	101	47	102	48
rect	101	48	102	49
rect	101	50	102	51
rect	101	51	102	52
rect	101	71	102	72
rect	101	72	102	73
rect	101	74	102	75
rect	101	75	102	76
rect	103	11	104	12
rect	103	12	104	13
rect	103	13	104	14
rect	103	14	104	15
rect	103	15	104	16
rect	103	16	104	17
rect	103	17	104	18
rect	103	18	104	19
rect	103	19	104	20
rect	103	20	104	21
rect	103	21	104	22
rect	103	23	104	24
rect	103	24	104	25
rect	103	26	104	27
rect	103	27	104	28
rect	103	29	104	30
rect	103	30	104	31
rect	103	32	104	33
rect	103	33	104	34
rect	103	35	104	36
rect	103	36	104	37
rect	103	37	104	38
rect	103	38	104	39
rect	103	39	104	40
rect	103	40	104	41
rect	103	41	104	42
rect	103	42	104	43
rect	103	43	104	44
rect	103	44	104	45
rect	103	45	104	46
rect	103	46	104	47
rect	103	47	104	48
rect	103	48	104	49
rect	103	50	104	51
rect	103	51	104	52
rect	103	53	104	54
rect	103	54	104	55
rect	103	55	104	56
rect	103	56	104	57
rect	103	57	104	58
rect	103	65	104	66
rect	103	66	104	67
rect	103	77	104	78
rect	103	78	104	79
rect	103	80	104	81
rect	103	81	104	82
rect	105	11	106	12
rect	105	12	106	13
rect	105	13	106	14
rect	105	14	106	15
rect	105	15	106	16
rect	105	16	106	17
rect	105	17	106	18
rect	105	18	106	19
rect	105	19	106	20
rect	105	20	106	21
rect	105	21	106	22
rect	105	44	106	45
rect	105	45	106	46
rect	105	46	106	47
rect	105	47	106	48
rect	105	48	106	49
rect	105	62	106	63
rect	105	63	106	64
rect	105	64	106	65
rect	105	65	106	66
rect	105	66	106	67
rect	105	74	106	75
rect	105	75	106	76
rect	105	77	106	78
rect	105	78	106	79
rect	105	80	106	81
rect	105	81	106	82
rect	105	82	106	83
rect	105	83	106	84
rect	105	84	106	85
rect	105	86	106	87
rect	105	87	106	88
rect	105	95	106	96
rect	105	96	106	97
rect	105	98	106	99
rect	105	99	106	100
rect	105	101	106	102
rect	105	102	106	103
rect	107	8	108	9
rect	107	9	108	10
rect	107	11	108	12
rect	107	12	108	13
rect	107	13	108	14
rect	107	14	108	15
rect	107	15	108	16
rect	107	16	108	17
rect	107	17	108	18
rect	107	18	108	19
rect	107	23	108	24
rect	107	24	108	25
rect	107	26	108	27
rect	107	27	108	28
rect	107	29	108	30
rect	107	30	108	31
rect	107	32	108	33
rect	107	33	108	34
rect	107	35	108	36
rect	107	36	108	37
rect	107	37	108	38
rect	107	38	108	39
rect	107	39	108	40
rect	107	40	108	41
rect	107	41	108	42
rect	107	42	108	43
rect	107	44	108	45
rect	107	45	108	46
rect	107	59	108	60
rect	107	60	108	61
rect	107	62	108	63
rect	107	63	108	64
rect	107	64	108	65
rect	107	65	108	66
rect	107	66	108	67
rect	107	68	108	69
rect	107	69	108	70
rect	107	71	108	72
rect	107	72	108	73
rect	107	73	108	74
rect	107	74	108	75
rect	107	75	108	76
rect	107	77	108	78
rect	107	78	108	79
rect	107	86	108	87
rect	107	87	108	88
rect	107	88	108	89
rect	107	89	108	90
rect	107	90	108	91
rect	107	91	108	92
rect	107	92	108	93
rect	107	93	108	94
rect	107	94	108	95
rect	107	95	108	96
rect	107	96	108	97
rect	107	98	108	99
rect	107	99	108	100
rect	109	5	110	6
rect	109	6	110	7
rect	109	7	110	8
rect	109	8	110	9
rect	109	9	110	10
rect	109	11	110	12
rect	109	12	110	13
rect	109	17	110	18
rect	109	18	110	19
rect	109	20	110	21
rect	109	21	110	22
rect	109	23	110	24
rect	109	24	110	25
rect	109	41	110	42
rect	109	42	110	43
rect	109	44	110	45
rect	109	45	110	46
rect	109	47	110	48
rect	109	48	110	49
rect	109	49	110	50
rect	109	50	110	51
rect	109	51	110	52
rect	109	53	110	54
rect	109	54	110	55
rect	109	55	110	56
rect	109	56	110	57
rect	109	57	110	58
rect	109	59	110	60
rect	109	60	110	61
rect	109	62	110	63
rect	109	63	110	64
rect	109	74	110	75
rect	109	75	110	76
rect	109	77	110	78
rect	109	78	110	79
rect	109	79	110	80
rect	109	80	110	81
rect	109	81	110	82
rect	109	82	110	83
rect	109	83	110	84
rect	109	84	110	85
rect	109	85	110	86
rect	109	86	110	87
rect	109	87	110	88
rect	109	88	110	89
rect	109	89	110	90
rect	109	90	110	91
rect	109	91	110	92
rect	109	92	110	93
rect	109	93	110	94
rect	109	94	110	95
rect	109	95	110	96
rect	109	96	110	97
rect	118	29	119	30
rect	118	30	119	31
rect	118	32	119	33
rect	118	33	119	34
rect	118	35	119	36
rect	118	36	119	37
rect	118	37	119	38
rect	118	38	119	39
rect	118	39	119	40
rect	120	8	121	9
rect	120	9	121	10
rect	120	11	121	12
rect	120	12	121	13
rect	120	14	121	15
rect	120	15	121	16
rect	120	17	121	18
rect	120	18	121	19
rect	120	26	121	27
rect	120	27	121	28
rect	120	28	121	29
rect	120	29	121	30
rect	120	30	121	31
rect	120	32	121	33
rect	120	33	121	34
rect	120	35	121	36
rect	120	36	121	37
rect	120	37	121	38
rect	120	38	121	39
rect	120	39	121	40
rect	120	40	121	41
rect	120	41	121	42
rect	120	42	121	43
rect	120	44	121	45
rect	120	45	121	46
rect	120	47	121	48
rect	120	48	121	49
rect	120	50	121	51
rect	120	51	121	52
rect	120	53	121	54
rect	120	54	121	55
rect	120	55	121	56
rect	120	56	121	57
rect	120	57	121	58
rect	120	58	121	59
rect	120	59	121	60
rect	120	60	121	61
rect	120	62	121	63
rect	120	63	121	64
rect	120	64	121	65
rect	120	65	121	66
rect	120	66	121	67
rect	120	67	121	68
rect	120	68	121	69
rect	120	69	121	70
rect	120	71	121	72
rect	120	72	121	73
rect	120	74	121	75
rect	120	75	121	76
rect	122	20	123	21
rect	122	21	123	22
rect	122	22	123	23
rect	122	23	123	24
rect	122	24	123	25
rect	122	26	123	27
rect	122	27	123	28
rect	122	28	123	29
rect	122	29	123	30
rect	122	30	123	31
rect	122	32	123	33
rect	122	33	123	34
rect	122	35	123	36
rect	122	36	123	37
rect	122	37	123	38
rect	122	38	123	39
rect	122	39	123	40
rect	122	40	123	41
rect	122	41	123	42
rect	122	42	123	43
rect	122	44	123	45
rect	122	45	123	46
rect	122	47	123	48
rect	122	48	123	49
rect	122	50	123	51
rect	122	51	123	52
rect	122	53	123	54
rect	122	54	123	55
rect	122	55	123	56
rect	122	56	123	57
rect	122	57	123	58
rect	122	58	123	59
rect	122	59	123	60
rect	122	60	123	61
rect	122	62	123	63
rect	122	63	123	64
rect	122	64	123	65
rect	122	65	123	66
rect	122	66	123	67
rect	122	67	123	68
rect	122	68	123	69
rect	122	69	123	70
rect	122	71	123	72
rect	122	72	123	73
rect	124	11	125	12
rect	124	12	125	13
rect	124	14	125	15
rect	124	15	125	16
rect	124	17	125	18
rect	124	18	125	19
rect	124	20	125	21
rect	124	21	125	22
rect	124	22	125	23
rect	124	23	125	24
rect	124	24	125	25
rect	124	26	125	27
rect	124	27	125	28
rect	124	28	125	29
rect	124	29	125	30
rect	124	30	125	31
rect	124	32	125	33
rect	124	33	125	34
rect	126	11	127	12
rect	126	12	127	13
rect	126	14	127	15
rect	126	15	127	16
rect	126	17	127	18
rect	126	18	127	19
rect	126	20	127	21
rect	126	21	127	22
rect	126	22	127	23
rect	126	23	127	24
rect	126	24	127	25
rect	126	26	127	27
rect	126	27	127	28
rect	126	28	127	29
rect	126	29	127	30
rect	126	30	127	31
rect	126	32	127	33
rect	126	33	127	34
rect	126	34	127	35
rect	126	35	127	36
rect	126	36	127	37
rect	126	37	127	38
rect	126	38	127	39
rect	126	39	127	40
rect	126	40	127	41
rect	126	41	127	42
rect	126	42	127	43
rect	126	44	127	45
rect	126	45	127	46
rect	126	47	127	48
rect	126	48	127	49
rect	126	50	127	51
rect	126	51	127	52
rect	126	53	127	54
rect	126	54	127	55
rect	126	55	127	56
rect	126	56	127	57
rect	126	57	127	58
rect	126	58	127	59
rect	126	59	127	60
rect	126	60	127	61
rect	126	62	127	63
rect	126	63	127	64
rect	126	64	127	65
rect	126	65	127	66
rect	126	66	127	67
rect	126	67	127	68
rect	126	68	127	69
rect	126	69	127	70
rect	128	5	129	6
rect	128	6	129	7
rect	128	7	129	8
rect	128	8	129	9
rect	128	9	129	10
rect	128	11	129	12
rect	128	12	129	13
rect	128	14	129	15
rect	128	15	129	16
rect	128	17	129	18
rect	128	18	129	19
rect	128	20	129	21
rect	128	21	129	22
rect	128	22	129	23
rect	128	23	129	24
rect	128	24	129	25
rect	128	26	129	27
rect	128	27	129	28
rect	128	28	129	29
rect	128	29	129	30
rect	128	30	129	31
rect	128	44	129	45
rect	128	45	129	46
rect	128	50	129	51
rect	128	51	129	52
rect	130	5	131	6
rect	130	6	131	7
rect	130	7	131	8
rect	130	8	131	9
rect	130	9	131	10
rect	130	11	131	12
rect	130	12	131	13
rect	130	14	131	15
rect	130	15	131	16
rect	130	17	131	18
rect	130	18	131	19
rect	130	20	131	21
rect	130	21	131	22
rect	130	22	131	23
rect	130	23	131	24
rect	130	24	131	25
rect	130	26	131	27
rect	130	27	131	28
rect	130	28	131	29
rect	130	29	131	30
rect	130	30	131	31
rect	130	31	131	32
rect	130	32	131	33
rect	130	33	131	34
rect	130	34	131	35
rect	130	35	131	36
rect	130	36	131	37
rect	130	37	131	38
rect	130	38	131	39
rect	130	39	131	40
rect	130	40	131	41
rect	130	41	131	42
rect	130	42	131	43
rect	130	43	131	44
rect	130	44	131	45
rect	130	45	131	46
rect	130	46	131	47
rect	130	47	131	48
rect	130	48	131	49
rect	130	49	131	50
rect	130	50	131	51
rect	130	51	131	52
rect	130	52	131	53
rect	130	53	131	54
rect	130	54	131	55
rect	130	55	131	56
rect	130	56	131	57
rect	130	57	131	58
rect	130	58	131	59
rect	130	59	131	60
rect	130	60	131	61
rect	139	14	140	15
rect	139	15	140	16
rect	139	17	140	18
rect	139	18	140	19
rect	141	11	142	12
rect	141	12	142	13
rect	141	13	142	14
rect	141	14	142	15
rect	141	15	142	16
rect	141	17	142	18
rect	141	18	142	19
rect	141	19	142	20
rect	141	20	142	21
rect	141	21	142	22
rect	141	22	142	23
rect	141	23	142	24
rect	141	24	142	25
rect	143	8	144	9
rect	143	9	144	10
rect	143	10	144	11
rect	143	11	144	12
rect	143	12	144	13
rect	143	13	144	14
rect	143	14	144	15
rect	143	15	144	16
<< metal2 >>
rect	1	4	2	5
rect	1	49	2	50
rect	2	4	3	5
rect	2	49	3	50
rect	3	1	4	2
rect	3	4	4	5
rect	3	7	4	8
rect	3	10	4	11
rect	3	13	4	14
rect	3	16	4	17
rect	3	19	4	20
rect	3	46	4	47
rect	3	49	4	50
rect	3	52	4	53
rect	10	7	11	8
rect	10	10	11	11
rect	10	19	11	20
rect	10	31	11	32
rect	10	46	11	47
rect	10	49	11	50
rect	10	52	11	53
rect	11	7	12	8
rect	11	10	12	11
rect	11	19	12	20
rect	11	49	12	50
rect	11	52	12	53
rect	12	7	13	8
rect	12	10	13	11
rect	12	19	13	20
rect	12	25	13	26
rect	12	49	13	50
rect	12	52	13	53
rect	12	67	13	68
rect	13	7	14	8
rect	13	10	14	11
rect	13	25	14	26
rect	13	49	14	50
rect	13	52	14	53
rect	13	67	14	68
rect	14	7	15	8
rect	14	10	15	11
rect	14	25	15	26
rect	14	28	15	29
rect	14	37	15	38
rect	14	46	15	47
rect	14	49	15	50
rect	14	52	15	53
rect	14	67	15	68
rect	15	7	16	8
rect	15	10	16	11
rect	15	25	16	26
rect	15	28	16	29
rect	15	37	16	38
rect	15	46	16	47
rect	15	49	16	50
rect	15	52	16	53
rect	15	67	16	68
rect	16	7	17	8
rect	16	10	17	11
rect	16	13	17	14
rect	16	25	17	26
rect	16	28	17	29
rect	16	37	17	38
rect	16	46	17	47
rect	16	49	17	50
rect	16	52	17	53
rect	16	61	17	62
rect	16	67	17	68
rect	17	7	18	8
rect	17	13	18	14
rect	17	25	18	26
rect	17	28	18	29
rect	17	37	18	38
rect	17	46	18	47
rect	17	49	18	50
rect	17	52	18	53
rect	17	61	18	62
rect	17	67	18	68
rect	18	7	19	8
rect	18	13	19	14
rect	18	16	19	17
rect	18	19	19	20
rect	18	25	19	26
rect	18	28	19	29
rect	18	37	19	38
rect	18	40	19	41
rect	18	46	19	47
rect	18	49	19	50
rect	18	52	19	53
rect	18	58	19	59
rect	18	61	19	62
rect	18	67	19	68
rect	18	73	19	74
rect	19	13	20	14
rect	19	16	20	17
rect	19	19	20	20
rect	19	25	20	26
rect	19	28	20	29
rect	19	37	20	38
rect	19	40	20	41
rect	19	46	20	47
rect	19	49	20	50
rect	19	58	20	59
rect	19	61	20	62
rect	19	67	20	68
rect	19	73	20	74
rect	20	1	21	2
rect	20	10	21	11
rect	20	13	21	14
rect	20	16	21	17
rect	20	19	21	20
rect	20	25	21	26
rect	20	28	21	29
rect	20	37	21	38
rect	20	40	21	41
rect	20	46	21	47
rect	20	49	21	50
rect	20	55	21	56
rect	20	58	21	59
rect	20	61	21	62
rect	20	64	21	65
rect	20	67	21	68
rect	20	73	21	74
rect	27	1	28	2
rect	27	7	28	8
rect	27	13	28	14
rect	27	16	28	17
rect	27	19	28	20
rect	27	25	28	26
rect	27	28	28	29
rect	27	37	28	38
rect	27	40	28	41
rect	27	43	28	44
rect	27	46	28	47
rect	27	49	28	50
rect	27	58	28	59
rect	27	61	28	62
rect	27	64	28	65
rect	27	67	28	68
rect	27	70	28	71
rect	28	1	29	2
rect	28	7	29	8
rect	28	13	29	14
rect	28	16	29	17
rect	28	19	29	20
rect	28	25	29	26
rect	28	28	29	29
rect	28	37	29	38
rect	28	40	29	41
rect	28	43	29	44
rect	28	46	29	47
rect	28	49	29	50
rect	28	58	29	59
rect	28	61	29	62
rect	28	67	29	68
rect	28	70	29	71
rect	29	1	30	2
rect	29	7	30	8
rect	29	13	30	14
rect	29	16	30	17
rect	29	19	30	20
rect	29	25	30	26
rect	29	28	30	29
rect	29	37	30	38
rect	29	40	30	41
rect	29	43	30	44
rect	29	46	30	47
rect	29	49	30	50
rect	29	58	30	59
rect	29	61	30	62
rect	29	67	30	68
rect	29	70	30	71
rect	29	73	30	74
rect	30	1	31	2
rect	30	7	31	8
rect	30	13	31	14
rect	30	16	31	17
rect	30	25	31	26
rect	30	28	31	29
rect	30	40	31	41
rect	30	43	31	44
rect	30	46	31	47
rect	30	58	31	59
rect	30	67	31	68
rect	30	70	31	71
rect	30	73	31	74
rect	31	1	32	2
rect	31	7	32	8
rect	31	13	32	14
rect	31	16	32	17
rect	31	25	32	26
rect	31	28	32	29
rect	31	40	32	41
rect	31	43	32	44
rect	31	46	32	47
rect	31	55	32	56
rect	31	58	32	59
rect	31	67	32	68
rect	31	70	32	71
rect	31	73	32	74
rect	31	79	32	80
rect	32	1	33	2
rect	32	7	33	8
rect	32	16	33	17
rect	32	25	33	26
rect	32	28	33	29
rect	32	40	33	41
rect	32	46	33	47
rect	32	55	33	56
rect	32	58	33	59
rect	32	70	33	71
rect	32	73	33	74
rect	32	79	33	80
rect	33	1	34	2
rect	33	7	34	8
rect	33	16	34	17
rect	33	22	34	23
rect	33	25	34	26
rect	33	28	34	29
rect	33	40	34	41
rect	33	46	34	47
rect	33	55	34	56
rect	33	58	34	59
rect	33	64	34	65
rect	33	70	34	71
rect	33	73	34	74
rect	33	76	34	77
rect	33	79	34	80
rect	34	16	35	17
rect	34	22	35	23
rect	34	25	35	26
rect	34	28	35	29
rect	34	40	35	41
rect	34	46	35	47
rect	34	55	35	56
rect	34	58	35	59
rect	34	64	35	65
rect	34	70	35	71
rect	34	73	35	74
rect	34	76	35	77
rect	34	79	35	80
rect	35	13	36	14
rect	35	16	36	17
rect	35	22	36	23
rect	35	25	36	26
rect	35	28	36	29
rect	35	40	36	41
rect	35	46	36	47
rect	35	55	36	56
rect	35	58	36	59
rect	35	64	36	65
rect	35	70	36	71
rect	35	73	36	74
rect	35	76	36	77
rect	35	79	36	80
rect	35	85	36	86
rect	36	13	37	14
rect	36	22	37	23
rect	36	25	37	26
rect	36	28	37	29
rect	36	55	37	56
rect	36	58	37	59
rect	36	64	37	65
rect	36	70	37	71
rect	36	73	37	74
rect	36	76	37	77
rect	36	79	37	80
rect	36	85	37	86
rect	37	1	38	2
rect	37	7	38	8
rect	37	10	38	11
rect	37	13	38	14
rect	37	19	38	20
rect	37	22	38	23
rect	37	25	38	26
rect	37	28	38	29
rect	37	31	38	32
rect	37	43	38	44
rect	37	52	38	53
rect	37	55	38	56
rect	37	58	38	59
rect	37	61	38	62
rect	37	64	38	65
rect	37	67	38	68
rect	37	70	38	71
rect	37	73	38	74
rect	37	76	38	77
rect	37	79	38	80
rect	37	85	38	86
rect	44	1	45	2
rect	44	4	45	5
rect	44	7	45	8
rect	44	10	45	11
rect	44	16	45	17
rect	44	19	45	20
rect	44	22	45	23
rect	44	25	45	26
rect	44	28	45	29
rect	44	31	45	32
rect	44	37	45	38
rect	44	43	45	44
rect	44	46	45	47
rect	44	52	45	53
rect	44	55	45	56
rect	44	58	45	59
rect	44	61	45	62
rect	44	64	45	65
rect	44	67	45	68
rect	44	70	45	71
rect	44	73	45	74
rect	44	76	45	77
rect	44	79	45	80
rect	44	85	45	86
rect	45	1	46	2
rect	45	4	46	5
rect	45	7	46	8
rect	45	10	46	11
rect	45	16	46	17
rect	45	19	46	20
rect	45	22	46	23
rect	45	25	46	26
rect	45	28	46	29
rect	45	31	46	32
rect	45	37	46	38
rect	45	43	46	44
rect	45	46	46	47
rect	45	52	46	53
rect	45	55	46	56
rect	45	64	46	65
rect	45	67	46	68
rect	45	70	46	71
rect	45	73	46	74
rect	45	76	46	77
rect	45	79	46	80
rect	45	85	46	86
rect	46	1	47	2
rect	46	4	47	5
rect	46	7	47	8
rect	46	10	47	11
rect	46	16	47	17
rect	46	19	47	20
rect	46	22	47	23
rect	46	25	47	26
rect	46	28	47	29
rect	46	31	47	32
rect	46	37	47	38
rect	46	43	47	44
rect	46	46	47	47
rect	46	52	47	53
rect	46	55	47	56
rect	46	64	47	65
rect	46	67	47	68
rect	46	70	47	71
rect	46	73	47	74
rect	46	76	47	77
rect	46	79	47	80
rect	46	85	47	86
rect	47	1	48	2
rect	47	4	48	5
rect	47	7	48	8
rect	47	10	48	11
rect	47	16	48	17
rect	47	19	48	20
rect	47	22	48	23
rect	47	25	48	26
rect	47	31	48	32
rect	47	37	48	38
rect	47	43	48	44
rect	47	46	48	47
rect	47	52	48	53
rect	47	67	48	68
rect	47	70	48	71
rect	47	73	48	74
rect	47	76	48	77
rect	47	79	48	80
rect	47	85	48	86
rect	48	1	49	2
rect	48	4	49	5
rect	48	7	49	8
rect	48	10	49	11
rect	48	16	49	17
rect	48	19	49	20
rect	48	22	49	23
rect	48	25	49	26
rect	48	31	49	32
rect	48	37	49	38
rect	48	40	49	41
rect	48	43	49	44
rect	48	46	49	47
rect	48	52	49	53
rect	48	67	49	68
rect	48	70	49	71
rect	48	73	49	74
rect	48	76	49	77
rect	48	79	49	80
rect	48	85	49	86
rect	49	1	50	2
rect	49	4	50	5
rect	49	7	50	8
rect	49	10	50	11
rect	49	16	50	17
rect	49	19	50	20
rect	49	22	50	23
rect	49	25	50	26
rect	49	40	50	41
rect	49	43	50	44
rect	49	46	50	47
rect	49	52	50	53
rect	49	70	50	71
rect	49	73	50	74
rect	49	76	50	77
rect	49	85	50	86
rect	50	1	51	2
rect	50	4	51	5
rect	50	7	51	8
rect	50	10	51	11
rect	50	16	51	17
rect	50	19	51	20
rect	50	22	51	23
rect	50	25	51	26
rect	50	28	51	29
rect	50	40	51	41
rect	50	43	51	44
rect	50	46	51	47
rect	50	52	51	53
rect	50	58	51	59
rect	50	70	51	71
rect	50	73	51	74
rect	50	76	51	77
rect	50	85	51	86
rect	51	1	52	2
rect	51	4	52	5
rect	51	7	52	8
rect	51	10	52	11
rect	51	16	52	17
rect	51	19	52	20
rect	51	25	52	26
rect	51	28	52	29
rect	51	40	52	41
rect	51	43	52	44
rect	51	46	52	47
rect	51	58	52	59
rect	51	70	52	71
rect	51	73	52	74
rect	51	85	52	86
rect	52	1	53	2
rect	52	4	53	5
rect	52	7	53	8
rect	52	10	53	11
rect	52	16	53	17
rect	52	19	53	20
rect	52	25	53	26
rect	52	28	53	29
rect	52	37	53	38
rect	52	40	53	41
rect	52	43	53	44
rect	52	46	53	47
rect	52	55	53	56
rect	52	58	53	59
rect	52	70	53	71
rect	52	73	53	74
rect	52	79	53	80
rect	52	85	53	86
rect	53	1	54	2
rect	53	19	54	20
rect	53	25	54	26
rect	53	28	54	29
rect	53	37	54	38
rect	53	40	54	41
rect	53	43	54	44
rect	53	46	54	47
rect	53	55	54	56
rect	53	58	54	59
rect	53	73	54	74
rect	53	79	54	80
rect	53	85	54	86
rect	54	1	55	2
rect	54	13	55	14
rect	54	19	55	20
rect	54	25	55	26
rect	54	28	55	29
rect	54	37	55	38
rect	54	40	55	41
rect	54	43	55	44
rect	54	46	55	47
rect	54	52	55	53
rect	54	55	55	56
rect	54	58	55	59
rect	54	73	55	74
rect	54	76	55	77
rect	54	79	55	80
rect	54	85	55	86
rect	55	13	56	14
rect	55	25	56	26
rect	55	28	56	29
rect	55	37	56	38
rect	55	40	56	41
rect	55	52	56	53
rect	55	55	56	56
rect	55	58	56	59
rect	55	76	56	77
rect	55	79	56	80
rect	55	85	56	86
rect	56	10	57	11
rect	56	13	57	14
rect	56	16	57	17
rect	56	22	57	23
rect	56	25	57	26
rect	56	28	57	29
rect	56	31	57	32
rect	56	37	57	38
rect	56	40	57	41
rect	56	52	57	53
rect	56	55	57	56
rect	56	58	57	59
rect	56	70	57	71
rect	56	76	57	77
rect	56	79	57	80
rect	56	85	57	86
rect	57	10	58	11
rect	57	13	58	14
rect	57	16	58	17
rect	57	22	58	23
rect	57	28	58	29
rect	57	31	58	32
rect	57	37	58	38
rect	57	40	58	41
rect	57	52	58	53
rect	57	55	58	56
rect	57	58	58	59
rect	57	70	58	71
rect	57	76	58	77
rect	57	79	58	80
rect	58	1	59	2
rect	58	7	59	8
rect	58	10	59	11
rect	58	13	59	14
rect	58	16	59	17
rect	58	19	59	20
rect	58	22	59	23
rect	58	28	59	29
rect	58	31	59	32
rect	58	34	59	35
rect	58	37	59	38
rect	58	40	59	41
rect	58	43	59	44
rect	58	46	59	47
rect	58	49	59	50
rect	58	52	59	53
rect	58	55	59	56
rect	58	58	59	59
rect	58	61	59	62
rect	58	64	59	65
rect	58	70	59	71
rect	58	73	59	74
rect	58	76	59	77
rect	58	79	59	80
rect	58	82	59	83
rect	58	88	59	89
rect	65	1	66	2
rect	65	4	66	5
rect	65	10	66	11
rect	65	13	66	14
rect	65	16	66	17
rect	65	19	66	20
rect	65	25	66	26
rect	65	28	66	29
rect	65	31	66	32
rect	65	34	66	35
rect	65	37	66	38
rect	65	40	66	41
rect	65	46	66	47
rect	65	49	66	50
rect	65	52	66	53
rect	65	55	66	56
rect	65	64	66	65
rect	65	70	66	71
rect	65	73	66	74
rect	65	76	66	77
rect	65	79	66	80
rect	65	82	66	83
rect	65	85	66	86
rect	65	91	66	92
rect	66	1	67	2
rect	66	4	67	5
rect	66	10	67	11
rect	66	13	67	14
rect	66	16	67	17
rect	66	19	67	20
rect	66	25	67	26
rect	66	28	67	29
rect	66	31	67	32
rect	66	34	67	35
rect	66	37	67	38
rect	66	40	67	41
rect	66	46	67	47
rect	66	49	67	50
rect	66	52	67	53
rect	66	55	67	56
rect	66	64	67	65
rect	66	70	67	71
rect	66	73	67	74
rect	66	79	67	80
rect	66	82	67	83
rect	66	91	67	92
rect	67	1	68	2
rect	67	4	68	5
rect	67	10	68	11
rect	67	13	68	14
rect	67	16	68	17
rect	67	19	68	20
rect	67	25	68	26
rect	67	28	68	29
rect	67	31	68	32
rect	67	34	68	35
rect	67	37	68	38
rect	67	40	68	41
rect	67	46	68	47
rect	67	49	68	50
rect	67	52	68	53
rect	67	55	68	56
rect	67	64	68	65
rect	67	70	68	71
rect	67	73	68	74
rect	67	79	68	80
rect	67	82	68	83
rect	67	91	68	92
rect	68	1	69	2
rect	68	4	69	5
rect	68	10	69	11
rect	68	13	69	14
rect	68	16	69	17
rect	68	19	69	20
rect	68	25	69	26
rect	68	28	69	29
rect	68	31	69	32
rect	68	34	69	35
rect	68	37	69	38
rect	68	40	69	41
rect	68	46	69	47
rect	68	49	69	50
rect	68	52	69	53
rect	68	55	69	56
rect	68	70	69	71
rect	68	73	69	74
rect	68	79	69	80
rect	68	82	69	83
rect	68	91	69	92
rect	69	1	70	2
rect	69	4	70	5
rect	69	10	70	11
rect	69	13	70	14
rect	69	16	70	17
rect	69	19	70	20
rect	69	25	70	26
rect	69	28	70	29
rect	69	31	70	32
rect	69	34	70	35
rect	69	37	70	38
rect	69	40	70	41
rect	69	46	70	47
rect	69	49	70	50
rect	69	52	70	53
rect	69	55	70	56
rect	69	70	70	71
rect	69	73	70	74
rect	69	79	70	80
rect	69	82	70	83
rect	69	85	70	86
rect	69	91	70	92
rect	70	1	71	2
rect	70	4	71	5
rect	70	10	71	11
rect	70	13	71	14
rect	70	16	71	17
rect	70	19	71	20
rect	70	25	71	26
rect	70	28	71	29
rect	70	31	71	32
rect	70	34	71	35
rect	70	37	71	38
rect	70	40	71	41
rect	70	46	71	47
rect	70	49	71	50
rect	70	52	71	53
rect	70	55	71	56
rect	70	70	71	71
rect	70	79	71	80
rect	70	82	71	83
rect	70	85	71	86
rect	70	91	71	92
rect	71	1	72	2
rect	71	4	72	5
rect	71	10	72	11
rect	71	13	72	14
rect	71	16	72	17
rect	71	19	72	20
rect	71	25	72	26
rect	71	28	72	29
rect	71	31	72	32
rect	71	34	72	35
rect	71	37	72	38
rect	71	40	72	41
rect	71	46	72	47
rect	71	49	72	50
rect	71	52	72	53
rect	71	55	72	56
rect	71	61	72	62
rect	71	70	72	71
rect	71	79	72	80
rect	71	82	72	83
rect	71	85	72	86
rect	71	91	72	92
rect	72	10	73	11
rect	72	16	73	17
rect	72	19	73	20
rect	72	28	73	29
rect	72	31	73	32
rect	72	34	73	35
rect	72	37	73	38
rect	72	40	73	41
rect	72	46	73	47
rect	72	49	73	50
rect	72	52	73	53
rect	72	61	73	62
rect	72	70	73	71
rect	72	79	73	80
rect	72	82	73	83
rect	72	85	73	86
rect	72	91	73	92
rect	73	10	74	11
rect	73	16	74	17
rect	73	19	74	20
rect	73	28	74	29
rect	73	31	74	32
rect	73	34	74	35
rect	73	37	74	38
rect	73	40	74	41
rect	73	46	74	47
rect	73	49	74	50
rect	73	52	74	53
rect	73	61	74	62
rect	73	64	74	65
rect	73	70	74	71
rect	73	79	74	80
rect	73	82	74	83
rect	73	85	74	86
rect	73	91	74	92
rect	74	10	75	11
rect	74	16	75	17
rect	74	28	75	29
rect	74	31	75	32
rect	74	34	75	35
rect	74	37	75	38
rect	74	40	75	41
rect	74	49	75	50
rect	74	52	75	53
rect	74	61	75	62
rect	74	64	75	65
rect	74	70	75	71
rect	74	79	75	80
rect	74	82	75	83
rect	74	85	75	86
rect	74	91	75	92
rect	75	4	76	5
rect	75	10	76	11
rect	75	16	76	17
rect	75	28	76	29
rect	75	31	76	32
rect	75	34	76	35
rect	75	37	76	38
rect	75	40	76	41
rect	75	49	76	50
rect	75	52	76	53
rect	75	61	76	62
rect	75	64	76	65
rect	75	70	76	71
rect	75	73	76	74
rect	75	79	76	80
rect	75	82	76	83
rect	75	85	76	86
rect	75	91	76	92
rect	76	4	77	5
rect	76	10	77	11
rect	76	16	77	17
rect	76	28	77	29
rect	76	31	77	32
rect	76	34	77	35
rect	76	37	77	38
rect	76	40	77	41
rect	76	61	77	62
rect	76	64	77	65
rect	76	70	77	71
rect	76	73	77	74
rect	76	79	77	80
rect	76	85	77	86
rect	76	91	77	92
rect	77	4	78	5
rect	77	10	78	11
rect	77	13	78	14
rect	77	16	78	17
rect	77	19	78	20
rect	77	28	78	29
rect	77	31	78	32
rect	77	34	78	35
rect	77	37	78	38
rect	77	40	78	41
rect	77	46	78	47
rect	77	55	78	56
rect	77	61	78	62
rect	77	64	78	65
rect	77	70	78	71
rect	77	73	78	74
rect	77	76	78	77
rect	77	79	78	80
rect	77	85	78	86
rect	77	91	78	92
rect	78	4	79	5
rect	78	13	79	14
rect	78	16	79	17
rect	78	19	79	20
rect	78	28	79	29
rect	78	31	79	32
rect	78	34	79	35
rect	78	37	79	38
rect	78	40	79	41
rect	78	46	79	47
rect	78	55	79	56
rect	78	61	79	62
rect	78	64	79	65
rect	78	73	79	74
rect	78	76	79	77
rect	78	85	79	86
rect	78	91	79	92
rect	79	4	80	5
rect	79	13	80	14
rect	79	16	80	17
rect	79	19	80	20
rect	79	22	80	23
rect	79	28	80	29
rect	79	31	80	32
rect	79	34	80	35
rect	79	37	80	38
rect	79	40	80	41
rect	79	43	80	44
rect	79	46	80	47
rect	79	52	80	53
rect	79	55	80	56
rect	79	61	80	62
rect	79	64	80	65
rect	79	73	80	74
rect	79	76	80	77
rect	79	82	80	83
rect	79	85	80	86
rect	79	88	80	89
rect	79	91	80	92
rect	80	4	81	5
rect	80	13	81	14
rect	80	16	81	17
rect	80	19	81	20
rect	80	22	81	23
rect	80	28	81	29
rect	80	31	81	32
rect	80	34	81	35
rect	80	37	81	38
rect	80	40	81	41
rect	80	43	81	44
rect	80	46	81	47
rect	80	52	81	53
rect	80	55	81	56
rect	80	61	81	62
rect	80	64	81	65
rect	80	73	81	74
rect	80	76	81	77
rect	80	82	81	83
rect	80	85	81	86
rect	80	88	81	89
rect	80	91	81	92
rect	81	4	82	5
rect	81	10	82	11
rect	81	13	82	14
rect	81	16	82	17
rect	81	19	82	20
rect	81	22	82	23
rect	81	28	82	29
rect	81	31	82	32
rect	81	34	82	35
rect	81	37	82	38
rect	81	40	82	41
rect	81	43	82	44
rect	81	46	82	47
rect	81	52	82	53
rect	81	55	82	56
rect	81	61	82	62
rect	81	64	82	65
rect	81	73	82	74
rect	81	76	82	77
rect	81	82	82	83
rect	81	85	82	86
rect	81	88	82	89
rect	81	91	82	92
rect	81	94	82	95
rect	82	4	83	5
rect	82	10	83	11
rect	82	13	83	14
rect	82	19	83	20
rect	82	22	83	23
rect	82	31	83	32
rect	82	34	83	35
rect	82	40	83	41
rect	82	43	83	44
rect	82	46	83	47
rect	82	52	83	53
rect	82	55	83	56
rect	82	61	83	62
rect	82	64	83	65
rect	82	73	83	74
rect	82	76	83	77
rect	82	82	83	83
rect	82	85	83	86
rect	82	88	83	89
rect	82	94	83	95
rect	83	4	84	5
rect	83	7	84	8
rect	83	10	84	11
rect	83	13	84	14
rect	83	19	84	20
rect	83	22	84	23
rect	83	25	84	26
rect	83	31	84	32
rect	83	34	84	35
rect	83	40	84	41
rect	83	43	84	44
rect	83	46	84	47
rect	83	52	84	53
rect	83	55	84	56
rect	83	61	84	62
rect	83	64	84	65
rect	83	73	84	74
rect	83	76	84	77
rect	83	82	84	83
rect	83	85	84	86
rect	83	88	84	89
rect	83	94	84	95
rect	84	4	85	5
rect	84	7	85	8
rect	84	10	85	11
rect	84	13	85	14
rect	84	19	85	20
rect	84	22	85	23
rect	84	25	85	26
rect	84	31	85	32
rect	84	34	85	35
rect	84	43	85	44
rect	84	46	85	47
rect	84	52	85	53
rect	84	55	85	56
rect	84	61	85	62
rect	84	64	85	65
rect	84	73	85	74
rect	84	76	85	77
rect	84	82	85	83
rect	84	85	85	86
rect	84	88	85	89
rect	84	94	85	95
rect	85	1	86	2
rect	85	4	86	5
rect	85	7	86	8
rect	85	10	86	11
rect	85	13	86	14
rect	85	16	86	17
rect	85	19	86	20
rect	85	22	86	23
rect	85	25	86	26
rect	85	28	86	29
rect	85	31	86	32
rect	85	34	86	35
rect	85	37	86	38
rect	85	43	86	44
rect	85	46	86	47
rect	85	49	86	50
rect	85	52	86	53
rect	85	55	86	56
rect	85	58	86	59
rect	85	61	86	62
rect	85	64	86	65
rect	85	67	86	68
rect	85	73	86	74
rect	85	76	86	77
rect	85	79	86	80
rect	85	82	86	83
rect	85	85	86	86
rect	85	88	86	89
rect	85	91	86	92
rect	85	94	86	95
rect	85	97	86	98
rect	85	103	86	104
rect	92	7	93	8
rect	92	10	93	11
rect	92	13	93	14
rect	92	16	93	17
rect	92	19	93	20
rect	92	22	93	23
rect	92	25	93	26
rect	92	28	93	29
rect	92	31	93	32
rect	92	34	93	35
rect	92	37	93	38
rect	92	40	93	41
rect	92	43	93	44
rect	92	46	93	47
rect	92	49	93	50
rect	92	58	93	59
rect	92	61	93	62
rect	92	64	93	65
rect	92	67	93	68
rect	92	70	93	71
rect	92	73	93	74
rect	92	76	93	77
rect	92	79	93	80
rect	92	82	93	83
rect	92	85	93	86
rect	92	88	93	89
rect	92	94	93	95
rect	92	97	93	98
rect	92	100	93	101
rect	92	103	93	104
rect	93	7	94	8
rect	93	10	94	11
rect	93	16	94	17
rect	93	19	94	20
rect	93	22	94	23
rect	93	25	94	26
rect	93	28	94	29
rect	93	31	94	32
rect	93	37	94	38
rect	93	40	94	41
rect	93	43	94	44
rect	93	46	94	47
rect	93	49	94	50
rect	93	58	94	59
rect	93	61	94	62
rect	93	64	94	65
rect	93	67	94	68
rect	93	70	94	71
rect	93	73	94	74
rect	93	76	94	77
rect	93	79	94	80
rect	93	82	94	83
rect	93	85	94	86
rect	93	88	94	89
rect	93	94	94	95
rect	93	97	94	98
rect	93	100	94	101
rect	93	103	94	104
rect	94	7	95	8
rect	94	10	95	11
rect	94	16	95	17
rect	94	19	95	20
rect	94	22	95	23
rect	94	25	95	26
rect	94	28	95	29
rect	94	31	95	32
rect	94	37	95	38
rect	94	40	95	41
rect	94	43	95	44
rect	94	46	95	47
rect	94	49	95	50
rect	94	58	95	59
rect	94	61	95	62
rect	94	64	95	65
rect	94	67	95	68
rect	94	70	95	71
rect	94	73	95	74
rect	94	76	95	77
rect	94	79	95	80
rect	94	82	95	83
rect	94	85	95	86
rect	94	88	95	89
rect	94	94	95	95
rect	94	97	95	98
rect	94	100	95	101
rect	94	103	95	104
rect	95	7	96	8
rect	95	10	96	11
rect	95	16	96	17
rect	95	19	96	20
rect	95	22	96	23
rect	95	25	96	26
rect	95	28	96	29
rect	95	37	96	38
rect	95	40	96	41
rect	95	43	96	44
rect	95	46	96	47
rect	95	49	96	50
rect	95	58	96	59
rect	95	61	96	62
rect	95	64	96	65
rect	95	67	96	68
rect	95	70	96	71
rect	95	73	96	74
rect	95	76	96	77
rect	95	79	96	80
rect	95	82	96	83
rect	95	85	96	86
rect	95	88	96	89
rect	95	94	96	95
rect	95	97	96	98
rect	95	100	96	101
rect	95	103	96	104
rect	96	7	97	8
rect	96	10	97	11
rect	96	16	97	17
rect	96	19	97	20
rect	96	22	97	23
rect	96	25	97	26
rect	96	28	97	29
rect	96	34	97	35
rect	96	37	97	38
rect	96	40	97	41
rect	96	43	97	44
rect	96	46	97	47
rect	96	49	97	50
rect	96	58	97	59
rect	96	61	97	62
rect	96	64	97	65
rect	96	67	97	68
rect	96	70	97	71
rect	96	73	97	74
rect	96	76	97	77
rect	96	79	97	80
rect	96	82	97	83
rect	96	85	97	86
rect	96	88	97	89
rect	96	94	97	95
rect	96	97	97	98
rect	96	100	97	101
rect	96	103	97	104
rect	97	7	98	8
rect	97	10	98	11
rect	97	16	98	17
rect	97	19	98	20
rect	97	22	98	23
rect	97	25	98	26
rect	97	28	98	29
rect	97	34	98	35
rect	97	37	98	38
rect	97	40	98	41
rect	97	46	98	47
rect	97	49	98	50
rect	97	58	98	59
rect	97	61	98	62
rect	97	64	98	65
rect	97	67	98	68
rect	97	70	98	71
rect	97	73	98	74
rect	97	76	98	77
rect	97	79	98	80
rect	97	82	98	83
rect	97	85	98	86
rect	97	88	98	89
rect	97	94	98	95
rect	97	97	98	98
rect	97	100	98	101
rect	97	103	98	104
rect	98	7	99	8
rect	98	10	99	11
rect	98	16	99	17
rect	98	19	99	20
rect	98	22	99	23
rect	98	25	99	26
rect	98	28	99	29
rect	98	31	99	32
rect	98	34	99	35
rect	98	37	99	38
rect	98	40	99	41
rect	98	46	99	47
rect	98	49	99	50
rect	98	58	99	59
rect	98	61	99	62
rect	98	64	99	65
rect	98	67	99	68
rect	98	70	99	71
rect	98	73	99	74
rect	98	76	99	77
rect	98	79	99	80
rect	98	82	99	83
rect	98	85	99	86
rect	98	88	99	89
rect	98	94	99	95
rect	98	97	99	98
rect	98	100	99	101
rect	98	103	99	104
rect	99	7	100	8
rect	99	10	100	11
rect	99	16	100	17
rect	99	22	100	23
rect	99	25	100	26
rect	99	28	100	29
rect	99	31	100	32
rect	99	34	100	35
rect	99	40	100	41
rect	99	46	100	47
rect	99	49	100	50
rect	99	58	100	59
rect	99	64	100	65
rect	99	67	100	68
rect	99	73	100	74
rect	99	76	100	77
rect	99	79	100	80
rect	99	82	100	83
rect	99	85	100	86
rect	99	88	100	89
rect	99	94	100	95
rect	99	97	100	98
rect	99	100	100	101
rect	99	103	100	104
rect	100	7	101	8
rect	100	10	101	11
rect	100	16	101	17
rect	100	22	101	23
rect	100	25	101	26
rect	100	28	101	29
rect	100	31	101	32
rect	100	34	101	35
rect	100	40	101	41
rect	100	46	101	47
rect	100	49	101	50
rect	100	58	101	59
rect	100	64	101	65
rect	100	67	101	68
rect	100	73	101	74
rect	100	76	101	77
rect	100	79	101	80
rect	100	82	101	83
rect	100	85	101	86
rect	100	88	101	89
rect	100	94	101	95
rect	100	97	101	98
rect	100	100	101	101
rect	100	103	101	104
rect	101	7	102	8
rect	101	10	102	11
rect	101	22	102	23
rect	101	25	102	26
rect	101	28	102	29
rect	101	31	102	32
rect	101	34	102	35
rect	101	49	102	50
rect	101	58	102	59
rect	101	64	102	65
rect	101	67	102	68
rect	101	73	102	74
rect	101	79	102	80
rect	101	82	102	83
rect	101	85	102	86
rect	101	88	102	89
rect	101	94	102	95
rect	101	97	102	98
rect	101	100	102	101
rect	101	103	102	104
rect	102	7	103	8
rect	102	10	103	11
rect	102	22	103	23
rect	102	25	103	26
rect	102	28	103	29
rect	102	31	103	32
rect	102	34	103	35
rect	102	49	103	50
rect	102	52	103	53
rect	102	58	103	59
rect	102	64	103	65
rect	102	67	103	68
rect	102	70	103	71
rect	102	73	103	74
rect	102	79	103	80
rect	102	82	103	83
rect	102	85	103	86
rect	102	88	103	89
rect	102	94	103	95
rect	102	97	103	98
rect	102	100	103	101
rect	102	103	103	104
rect	103	7	104	8
rect	103	22	104	23
rect	103	25	104	26
rect	103	28	104	29
rect	103	31	104	32
rect	103	34	104	35
rect	103	49	104	50
rect	103	52	104	53
rect	103	70	104	71
rect	103	73	104	74
rect	103	79	104	80
rect	103	85	104	86
rect	103	88	104	89
rect	103	94	104	95
rect	103	97	104	98
rect	103	100	104	101
rect	103	103	104	104
rect	104	7	105	8
rect	104	22	105	23
rect	104	25	105	26
rect	104	28	105	29
rect	104	31	105	32
rect	104	34	105	35
rect	104	49	105	50
rect	104	52	105	53
rect	104	70	105	71
rect	104	73	105	74
rect	104	76	105	77
rect	104	79	105	80
rect	104	85	105	86
rect	104	88	105	89
rect	104	94	105	95
rect	104	97	105	98
rect	104	100	105	101
rect	104	103	105	104
rect	105	7	106	8
rect	105	25	106	26
rect	105	28	106	29
rect	105	31	106	32
rect	105	34	106	35
rect	105	52	106	53
rect	105	70	106	71
rect	105	76	106	77
rect	105	79	106	80
rect	105	85	106	86
rect	105	97	106	98
rect	105	100	106	101
rect	106	7	107	8
rect	106	10	107	11
rect	106	25	107	26
rect	106	28	107	29
rect	106	31	107	32
rect	106	34	107	35
rect	106	43	107	44
rect	106	52	107	53
rect	106	61	107	62
rect	106	67	107	68
rect	106	70	107	71
rect	106	76	107	77
rect	106	79	107	80
rect	106	85	107	86
rect	106	97	107	98
rect	106	100	107	101
rect	107	10	108	11
rect	107	25	108	26
rect	107	28	108	29
rect	107	31	108	32
rect	107	34	108	35
rect	107	43	108	44
rect	107	52	108	53
rect	107	61	108	62
rect	107	67	108	68
rect	107	70	108	71
rect	107	76	108	77
rect	107	97	108	98
rect	108	10	109	11
rect	108	19	109	20
rect	108	22	109	23
rect	108	25	109	26
rect	108	28	109	29
rect	108	31	109	32
rect	108	34	109	35
rect	108	43	109	44
rect	108	46	109	47
rect	108	52	109	53
rect	108	58	109	59
rect	108	61	109	62
rect	108	67	109	68
rect	108	70	109	71
rect	108	76	109	77
rect	108	97	109	98
rect	109	10	110	11
rect	109	19	110	20
rect	109	22	110	23
rect	109	28	110	29
rect	109	31	110	32
rect	109	34	110	35
rect	109	43	110	44
rect	109	46	110	47
rect	109	52	110	53
rect	109	58	110	59
rect	109	61	110	62
rect	109	67	110	68
rect	109	70	110	71
rect	109	76	110	77
rect	110	4	111	5
rect	110	10	111	11
rect	110	13	111	14
rect	110	16	111	17
rect	110	19	111	20
rect	110	22	111	23
rect	110	28	111	29
rect	110	31	111	32
rect	110	34	111	35
rect	110	40	111	41
rect	110	43	111	44
rect	110	46	111	47
rect	110	52	111	53
rect	110	58	111	59
rect	110	61	111	62
rect	110	64	111	65
rect	110	67	111	68
rect	110	70	111	71
rect	110	73	111	74
rect	110	76	111	77
rect	117	4	118	5
rect	117	7	118	8
rect	117	10	118	11
rect	117	13	118	14
rect	117	16	118	17
rect	117	19	118	20
rect	117	28	118	29
rect	117	31	118	32
rect	117	34	118	35
rect	117	40	118	41
rect	117	43	118	44
rect	117	46	118	47
rect	117	49	118	50
rect	117	52	118	53
rect	117	61	118	62
rect	117	70	118	71
rect	117	73	118	74
rect	117	76	118	77
rect	118	4	119	5
rect	118	7	119	8
rect	118	10	119	11
rect	118	13	119	14
rect	118	16	119	17
rect	118	19	119	20
rect	118	31	119	32
rect	118	34	119	35
rect	118	43	119	44
rect	118	46	119	47
rect	118	49	119	50
rect	118	52	119	53
rect	118	61	119	62
rect	118	70	119	71
rect	118	73	119	74
rect	118	76	119	77
rect	119	4	120	5
rect	119	7	120	8
rect	119	10	120	11
rect	119	13	120	14
rect	119	16	120	17
rect	119	19	120	20
rect	119	31	120	32
rect	119	34	120	35
rect	119	43	120	44
rect	119	46	120	47
rect	119	49	120	50
rect	119	52	120	53
rect	119	61	120	62
rect	119	70	120	71
rect	119	73	120	74
rect	119	76	120	77
rect	120	4	121	5
rect	120	10	121	11
rect	120	13	121	14
rect	120	16	121	17
rect	120	31	121	32
rect	120	34	121	35
rect	120	43	121	44
rect	120	46	121	47
rect	120	49	121	50
rect	120	52	121	53
rect	120	61	121	62
rect	120	70	121	71
rect	120	73	121	74
rect	121	4	122	5
rect	121	10	122	11
rect	121	13	122	14
rect	121	16	122	17
rect	121	25	122	26
rect	121	31	122	32
rect	121	34	122	35
rect	121	43	122	44
rect	121	46	122	47
rect	121	49	122	50
rect	121	52	122	53
rect	121	61	122	62
rect	121	70	122	71
rect	121	73	122	74
rect	122	4	123	5
rect	122	10	123	11
rect	122	13	123	14
rect	122	16	123	17
rect	122	25	123	26
rect	122	31	123	32
rect	122	34	123	35
rect	122	43	123	44
rect	122	46	123	47
rect	122	49	123	50
rect	122	52	123	53
rect	122	61	123	62
rect	122	70	123	71
rect	123	4	124	5
rect	123	10	124	11
rect	123	13	124	14
rect	123	16	124	17
rect	123	19	124	20
rect	123	25	124	26
rect	123	31	124	32
rect	123	34	124	35
rect	123	43	124	44
rect	123	46	124	47
rect	123	49	124	50
rect	123	52	124	53
rect	123	61	124	62
rect	123	70	124	71
rect	124	4	125	5
rect	124	13	125	14
rect	124	16	125	17
rect	124	19	125	20
rect	124	25	125	26
rect	124	31	125	32
rect	124	43	125	44
rect	124	46	125	47
rect	124	49	125	50
rect	124	52	125	53
rect	124	61	125	62
rect	124	70	125	71
rect	125	4	126	5
rect	125	13	126	14
rect	125	16	126	17
rect	125	19	126	20
rect	125	25	126	26
rect	125	31	126	32
rect	125	43	126	44
rect	125	46	126	47
rect	125	49	126	50
rect	125	52	126	53
rect	125	61	126	62
rect	125	70	126	71
rect	126	4	127	5
rect	126	13	127	14
rect	126	16	127	17
rect	126	19	127	20
rect	126	25	127	26
rect	126	31	127	32
rect	126	43	127	44
rect	126	46	127	47
rect	126	49	127	50
rect	126	52	127	53
rect	126	61	127	62
rect	127	4	128	5
rect	127	10	128	11
rect	127	13	128	14
rect	127	16	128	17
rect	127	19	128	20
rect	127	25	128	26
rect	127	31	128	32
rect	127	43	128	44
rect	127	46	128	47
rect	127	49	128	50
rect	127	52	128	53
rect	127	61	128	62
rect	128	10	129	11
rect	128	13	129	14
rect	128	16	129	17
rect	128	19	129	20
rect	128	25	129	26
rect	128	61	129	62
rect	129	10	130	11
rect	129	13	130	14
rect	129	16	130	17
rect	129	19	130	20
rect	129	25	130	26
rect	129	61	130	62
rect	130	10	131	11
rect	130	13	131	14
rect	130	16	131	17
rect	130	19	131	20
rect	130	25	131	26
rect	131	4	132	5
rect	131	10	132	11
rect	131	13	132	14
rect	131	16	132	17
rect	131	19	132	20
rect	131	25	132	26
rect	138	7	139	8
rect	138	10	139	11
rect	138	13	139	14
rect	138	16	139	17
rect	138	19	139	20
rect	138	25	139	26
rect	139	7	140	8
rect	139	10	140	11
rect	139	16	140	17
rect	139	25	140	26
rect	140	7	141	8
rect	140	10	141	11
rect	140	16	141	17
rect	140	25	141	26
rect	141	7	142	8
rect	141	16	142	17
rect	142	7	143	8
rect	142	16	143	17
