magic
tech scmos
timestamp
<< pdiffusion >>
rect	6	0	7	1
rect	6	2	7	3
rect	6	3	7	4
rect	6	5	7	6
rect	6	6	7	7
rect	6	8	7	9
rect	6	9	7	10
rect	6	11	7	12
rect	6	12	7	13
rect	6	14	7	15
rect	6	15	7	16
rect	6	17	7	18
rect	6	18	7	19
rect	6	20	7	21
rect	6	21	7	22
rect	6	23	7	24
rect	6	24	7	25
rect	6	26	7	27
rect	6	27	7	28
rect	6	29	7	30
rect	6	30	7	31
rect	6	32	7	33
rect	6	33	7	34
rect	6	35	7	36
rect	6	36	7	37
rect	6	38	7	39
rect	6	39	7	40
rect	6	41	7	42
rect	6	42	7	43
rect	6	44	7	45
rect	6	45	7	46
rect	6	47	7	48
rect	6	48	7	49
rect	6	50	7	51
rect	6	51	7	52
rect	6	53	7	54
rect	6	54	7	55
rect	6	56	7	57
rect	6	57	7	58
rect	6	59	7	60
rect	6	60	7	61
rect	6	62	7	63
rect	6	63	7	64
rect	6	65	7	66
rect	6	66	7	67
rect	6	68	7	69
rect	6	69	7	70
rect	6	71	7	72
rect	6	72	7	73
rect	6	74	7	75
rect	6	75	7	76
rect	6	77	7	78
rect	6	78	7	79
rect	6	80	7	81
rect	6	81	7	82
rect	6	83	7	84
rect	6	84	7	85
rect	6	86	7	87
rect	6	87	7	88
rect	6	89	7	90
rect	6	90	7	91
rect	6	92	7	93
rect	6	93	7	94
rect	6	95	7	96
rect	6	96	7	97
rect	6	98	7	99
rect	6	99	7	100
rect	6	101	7	102
rect	6	102	7	103
rect	6	104	7	105
rect	6	105	7	106
rect	6	107	7	108
rect	6	108	7	109
rect	6	110	7	111
rect	6	111	7	112
rect	6	113	7	114
rect	6	114	7	115
rect	6	116	7	117
rect	6	117	7	118
rect	6	119	7	120
rect	6	120	7	121
rect	6	122	7	123
rect	6	123	7	124
rect	6	125	7	126
rect	6	126	7	127
rect	6	128	7	129
rect	6	129	7	130
rect	6	131	7	132
rect	6	132	7	133
rect	6	134	7	135
rect	6	135	7	136
rect	6	137	7	138
rect	6	138	7	139
rect	6	140	7	141
rect	6	141	7	142
rect	6	143	7	144
rect	6	144	7	145
rect	6	146	7	147
rect	6	147	7	148
rect	6	149	7	150
rect	6	150	7	151
rect	6	152	7	153
rect	6	153	7	154
rect	6	155	7	156
rect	6	156	7	157
rect	6	158	7	159
rect	6	159	7	160
rect	6	161	7	162
rect	6	162	7	163
rect	6	164	7	165
rect	6	165	7	166
rect	6	167	7	168
rect	6	168	7	169
rect	6	170	7	171
rect	6	171	7	172
rect	6	173	7	174
rect	7	0	8	1
rect	7	2	8	3
rect	7	3	8	4
rect	7	5	8	6
rect	7	6	8	7
rect	7	8	8	9
rect	7	9	8	10
rect	7	11	8	12
rect	7	12	8	13
rect	7	14	8	15
rect	7	15	8	16
rect	7	17	8	18
rect	7	18	8	19
rect	7	20	8	21
rect	7	21	8	22
rect	7	23	8	24
rect	7	24	8	25
rect	7	26	8	27
rect	7	27	8	28
rect	7	29	8	30
rect	7	30	8	31
rect	7	32	8	33
rect	7	33	8	34
rect	7	35	8	36
rect	7	36	8	37
rect	7	38	8	39
rect	7	39	8	40
rect	7	41	8	42
rect	7	42	8	43
rect	7	44	8	45
rect	7	45	8	46
rect	7	47	8	48
rect	7	48	8	49
rect	7	50	8	51
rect	7	51	8	52
rect	7	53	8	54
rect	7	54	8	55
rect	7	56	8	57
rect	7	57	8	58
rect	7	59	8	60
rect	7	60	8	61
rect	7	62	8	63
rect	7	63	8	64
rect	7	65	8	66
rect	7	66	8	67
rect	7	68	8	69
rect	7	69	8	70
rect	7	71	8	72
rect	7	72	8	73
rect	7	74	8	75
rect	7	75	8	76
rect	7	77	8	78
rect	7	78	8	79
rect	7	80	8	81
rect	7	81	8	82
rect	7	83	8	84
rect	7	84	8	85
rect	7	86	8	87
rect	7	87	8	88
rect	7	89	8	90
rect	7	90	8	91
rect	7	92	8	93
rect	7	93	8	94
rect	7	95	8	96
rect	7	96	8	97
rect	7	98	8	99
rect	7	99	8	100
rect	7	101	8	102
rect	7	102	8	103
rect	7	104	8	105
rect	7	105	8	106
rect	7	107	8	108
rect	7	108	8	109
rect	7	110	8	111
rect	7	111	8	112
rect	7	113	8	114
rect	7	114	8	115
rect	7	116	8	117
rect	7	117	8	118
rect	7	119	8	120
rect	7	120	8	121
rect	7	122	8	123
rect	7	123	8	124
rect	7	125	8	126
rect	7	126	8	127
rect	7	128	8	129
rect	7	129	8	130
rect	7	131	8	132
rect	7	132	8	133
rect	7	134	8	135
rect	7	135	8	136
rect	7	137	8	138
rect	7	138	8	139
rect	7	140	8	141
rect	7	141	8	142
rect	7	143	8	144
rect	7	144	8	145
rect	7	146	8	147
rect	7	147	8	148
rect	7	149	8	150
rect	7	150	8	151
rect	7	152	8	153
rect	7	153	8	154
rect	7	155	8	156
rect	7	156	8	157
rect	7	158	8	159
rect	7	159	8	160
rect	7	161	8	162
rect	7	162	8	163
rect	7	164	8	165
rect	7	165	8	166
rect	7	167	8	168
rect	7	168	8	169
rect	7	170	8	171
rect	7	171	8	172
rect	7	173	8	174
rect	8	0	9	1
rect	8	2	9	3
rect	8	3	9	4
rect	8	5	9	6
rect	8	6	9	7
rect	8	8	9	9
rect	8	9	9	10
rect	8	11	9	12
rect	8	12	9	13
rect	8	14	9	15
rect	8	15	9	16
rect	8	17	9	18
rect	8	18	9	19
rect	8	20	9	21
rect	8	21	9	22
rect	8	23	9	24
rect	8	24	9	25
rect	8	26	9	27
rect	8	27	9	28
rect	8	29	9	30
rect	8	30	9	31
rect	8	32	9	33
rect	8	33	9	34
rect	8	35	9	36
rect	8	36	9	37
rect	8	38	9	39
rect	8	39	9	40
rect	8	41	9	42
rect	8	42	9	43
rect	8	44	9	45
rect	8	45	9	46
rect	8	47	9	48
rect	8	48	9	49
rect	8	50	9	51
rect	8	51	9	52
rect	8	53	9	54
rect	8	54	9	55
rect	8	56	9	57
rect	8	57	9	58
rect	8	59	9	60
rect	8	60	9	61
rect	8	62	9	63
rect	8	63	9	64
rect	8	65	9	66
rect	8	66	9	67
rect	8	68	9	69
rect	8	69	9	70
rect	8	71	9	72
rect	8	72	9	73
rect	8	74	9	75
rect	8	75	9	76
rect	8	77	9	78
rect	8	78	9	79
rect	8	80	9	81
rect	8	81	9	82
rect	8	83	9	84
rect	8	84	9	85
rect	8	86	9	87
rect	8	87	9	88
rect	8	89	9	90
rect	8	90	9	91
rect	8	92	9	93
rect	8	93	9	94
rect	8	95	9	96
rect	8	96	9	97
rect	8	98	9	99
rect	8	99	9	100
rect	8	101	9	102
rect	8	102	9	103
rect	8	104	9	105
rect	8	105	9	106
rect	8	107	9	108
rect	8	108	9	109
rect	8	110	9	111
rect	8	111	9	112
rect	8	113	9	114
rect	8	114	9	115
rect	8	116	9	117
rect	8	117	9	118
rect	8	119	9	120
rect	8	120	9	121
rect	8	122	9	123
rect	8	123	9	124
rect	8	125	9	126
rect	8	126	9	127
rect	8	128	9	129
rect	8	129	9	130
rect	8	131	9	132
rect	8	132	9	133
rect	8	134	9	135
rect	8	135	9	136
rect	8	137	9	138
rect	8	138	9	139
rect	8	140	9	141
rect	8	141	9	142
rect	8	143	9	144
rect	8	144	9	145
rect	8	146	9	147
rect	8	147	9	148
rect	8	149	9	150
rect	8	150	9	151
rect	8	152	9	153
rect	8	153	9	154
rect	8	155	9	156
rect	8	156	9	157
rect	8	158	9	159
rect	8	159	9	160
rect	8	161	9	162
rect	8	162	9	163
rect	8	164	9	165
rect	8	165	9	166
rect	8	167	9	168
rect	8	168	9	169
rect	8	170	9	171
rect	8	171	9	172
rect	8	173	9	174
rect	9	0	10	1
rect	9	2	10	3
rect	9	3	10	4
rect	9	5	10	6
rect	9	6	10	7
rect	9	8	10	9
rect	9	9	10	10
rect	9	11	10	12
rect	9	12	10	13
rect	9	14	10	15
rect	9	15	10	16
rect	9	17	10	18
rect	9	18	10	19
rect	9	20	10	21
rect	9	21	10	22
rect	9	23	10	24
rect	9	24	10	25
rect	9	26	10	27
rect	9	27	10	28
rect	9	29	10	30
rect	9	30	10	31
rect	9	32	10	33
rect	9	33	10	34
rect	9	35	10	36
rect	9	36	10	37
rect	9	38	10	39
rect	9	39	10	40
rect	9	41	10	42
rect	9	42	10	43
rect	9	44	10	45
rect	9	45	10	46
rect	9	47	10	48
rect	9	48	10	49
rect	9	50	10	51
rect	9	51	10	52
rect	9	53	10	54
rect	9	54	10	55
rect	9	56	10	57
rect	9	57	10	58
rect	9	59	10	60
rect	9	60	10	61
rect	9	62	10	63
rect	9	63	10	64
rect	9	65	10	66
rect	9	66	10	67
rect	9	68	10	69
rect	9	69	10	70
rect	9	71	10	72
rect	9	72	10	73
rect	9	74	10	75
rect	9	75	10	76
rect	9	77	10	78
rect	9	78	10	79
rect	9	80	10	81
rect	9	81	10	82
rect	9	83	10	84
rect	9	84	10	85
rect	9	86	10	87
rect	9	87	10	88
rect	9	89	10	90
rect	9	90	10	91
rect	9	92	10	93
rect	9	93	10	94
rect	9	95	10	96
rect	9	96	10	97
rect	9	98	10	99
rect	9	99	10	100
rect	9	101	10	102
rect	9	102	10	103
rect	9	104	10	105
rect	9	105	10	106
rect	9	107	10	108
rect	9	108	10	109
rect	9	110	10	111
rect	9	111	10	112
rect	9	113	10	114
rect	9	114	10	115
rect	9	116	10	117
rect	9	117	10	118
rect	9	119	10	120
rect	9	120	10	121
rect	9	122	10	123
rect	9	123	10	124
rect	9	125	10	126
rect	9	126	10	127
rect	9	128	10	129
rect	9	129	10	130
rect	9	131	10	132
rect	9	132	10	133
rect	9	134	10	135
rect	9	135	10	136
rect	9	137	10	138
rect	9	138	10	139
rect	9	140	10	141
rect	9	141	10	142
rect	9	143	10	144
rect	9	144	10	145
rect	9	146	10	147
rect	9	147	10	148
rect	9	149	10	150
rect	9	150	10	151
rect	9	152	10	153
rect	9	153	10	154
rect	9	155	10	156
rect	9	156	10	157
rect	9	158	10	159
rect	9	159	10	160
rect	9	161	10	162
rect	9	162	10	163
rect	9	164	10	165
rect	9	165	10	166
rect	9	167	10	168
rect	9	168	10	169
rect	9	170	10	171
rect	9	171	10	172
rect	9	173	10	174
rect	10	0	11	1
rect	10	2	11	3
rect	10	3	11	4
rect	10	5	11	6
rect	10	6	11	7
rect	10	8	11	9
rect	10	9	11	10
rect	10	11	11	12
rect	10	12	11	13
rect	10	14	11	15
rect	10	15	11	16
rect	10	17	11	18
rect	10	18	11	19
rect	10	20	11	21
rect	10	21	11	22
rect	10	23	11	24
rect	10	24	11	25
rect	10	26	11	27
rect	10	27	11	28
rect	10	29	11	30
rect	10	30	11	31
rect	10	32	11	33
rect	10	33	11	34
rect	10	35	11	36
rect	10	36	11	37
rect	10	38	11	39
rect	10	39	11	40
rect	10	41	11	42
rect	10	42	11	43
rect	10	44	11	45
rect	10	45	11	46
rect	10	47	11	48
rect	10	48	11	49
rect	10	50	11	51
rect	10	51	11	52
rect	10	53	11	54
rect	10	54	11	55
rect	10	56	11	57
rect	10	57	11	58
rect	10	59	11	60
rect	10	60	11	61
rect	10	62	11	63
rect	10	63	11	64
rect	10	65	11	66
rect	10	66	11	67
rect	10	68	11	69
rect	10	69	11	70
rect	10	71	11	72
rect	10	72	11	73
rect	10	74	11	75
rect	10	75	11	76
rect	10	77	11	78
rect	10	78	11	79
rect	10	80	11	81
rect	10	81	11	82
rect	10	83	11	84
rect	10	84	11	85
rect	10	86	11	87
rect	10	87	11	88
rect	10	89	11	90
rect	10	90	11	91
rect	10	92	11	93
rect	10	93	11	94
rect	10	95	11	96
rect	10	96	11	97
rect	10	98	11	99
rect	10	99	11	100
rect	10	101	11	102
rect	10	102	11	103
rect	10	104	11	105
rect	10	105	11	106
rect	10	107	11	108
rect	10	108	11	109
rect	10	110	11	111
rect	10	111	11	112
rect	10	113	11	114
rect	10	114	11	115
rect	10	116	11	117
rect	10	117	11	118
rect	10	119	11	120
rect	10	120	11	121
rect	10	122	11	123
rect	10	123	11	124
rect	10	125	11	126
rect	10	126	11	127
rect	10	128	11	129
rect	10	129	11	130
rect	10	131	11	132
rect	10	132	11	133
rect	10	134	11	135
rect	10	135	11	136
rect	10	137	11	138
rect	10	138	11	139
rect	10	140	11	141
rect	10	141	11	142
rect	10	143	11	144
rect	10	144	11	145
rect	10	146	11	147
rect	10	147	11	148
rect	10	149	11	150
rect	10	150	11	151
rect	10	152	11	153
rect	10	153	11	154
rect	10	155	11	156
rect	10	156	11	157
rect	10	158	11	159
rect	10	159	11	160
rect	10	161	11	162
rect	10	162	11	163
rect	10	164	11	165
rect	10	165	11	166
rect	10	167	11	168
rect	10	168	11	169
rect	10	170	11	171
rect	10	171	11	172
rect	10	173	11	174
rect	11	0	12	1
rect	11	2	12	3
rect	11	3	12	4
rect	11	5	12	6
rect	11	6	12	7
rect	11	8	12	9
rect	11	9	12	10
rect	11	11	12	12
rect	11	12	12	13
rect	11	14	12	15
rect	11	15	12	16
rect	11	17	12	18
rect	11	18	12	19
rect	11	20	12	21
rect	11	21	12	22
rect	11	23	12	24
rect	11	24	12	25
rect	11	26	12	27
rect	11	27	12	28
rect	11	29	12	30
rect	11	30	12	31
rect	11	32	12	33
rect	11	33	12	34
rect	11	35	12	36
rect	11	36	12	37
rect	11	38	12	39
rect	11	39	12	40
rect	11	41	12	42
rect	11	42	12	43
rect	11	44	12	45
rect	11	45	12	46
rect	11	47	12	48
rect	11	48	12	49
rect	11	50	12	51
rect	11	51	12	52
rect	11	53	12	54
rect	11	54	12	55
rect	11	56	12	57
rect	11	57	12	58
rect	11	59	12	60
rect	11	60	12	61
rect	11	62	12	63
rect	11	63	12	64
rect	11	65	12	66
rect	11	66	12	67
rect	11	68	12	69
rect	11	69	12	70
rect	11	71	12	72
rect	11	72	12	73
rect	11	74	12	75
rect	11	75	12	76
rect	11	77	12	78
rect	11	78	12	79
rect	11	80	12	81
rect	11	81	12	82
rect	11	83	12	84
rect	11	84	12	85
rect	11	86	12	87
rect	11	87	12	88
rect	11	89	12	90
rect	11	90	12	91
rect	11	92	12	93
rect	11	93	12	94
rect	11	95	12	96
rect	11	96	12	97
rect	11	98	12	99
rect	11	99	12	100
rect	11	101	12	102
rect	11	102	12	103
rect	11	104	12	105
rect	11	105	12	106
rect	11	107	12	108
rect	11	108	12	109
rect	11	110	12	111
rect	11	111	12	112
rect	11	113	12	114
rect	11	114	12	115
rect	11	116	12	117
rect	11	117	12	118
rect	11	119	12	120
rect	11	120	12	121
rect	11	122	12	123
rect	11	123	12	124
rect	11	125	12	126
rect	11	126	12	127
rect	11	128	12	129
rect	11	129	12	130
rect	11	131	12	132
rect	11	132	12	133
rect	11	134	12	135
rect	11	135	12	136
rect	11	137	12	138
rect	11	138	12	139
rect	11	140	12	141
rect	11	141	12	142
rect	11	143	12	144
rect	11	144	12	145
rect	11	146	12	147
rect	11	147	12	148
rect	11	149	12	150
rect	11	150	12	151
rect	11	152	12	153
rect	11	153	12	154
rect	11	155	12	156
rect	11	156	12	157
rect	11	158	12	159
rect	11	159	12	160
rect	11	161	12	162
rect	11	162	12	163
rect	11	164	12	165
rect	11	165	12	166
rect	11	167	12	168
rect	11	168	12	169
rect	11	170	12	171
rect	11	171	12	172
rect	11	173	12	174
rect	13	0	14	1
rect	13	2	14	3
rect	13	3	14	4
rect	13	5	14	6
rect	13	6	14	7
rect	13	8	14	9
rect	13	9	14	10
rect	13	11	14	12
rect	13	12	14	13
rect	13	14	14	15
rect	13	15	14	16
rect	13	17	14	18
rect	13	18	14	19
rect	13	20	14	21
rect	13	21	14	22
rect	13	23	14	24
rect	13	24	14	25
rect	13	26	14	27
rect	13	27	14	28
rect	13	29	14	30
rect	13	30	14	31
rect	13	32	14	33
rect	13	33	14	34
rect	13	35	14	36
rect	13	36	14	37
rect	13	38	14	39
rect	13	39	14	40
rect	13	41	14	42
rect	13	42	14	43
rect	13	44	14	45
rect	13	45	14	46
rect	13	47	14	48
rect	13	48	14	49
rect	13	50	14	51
rect	13	51	14	52
rect	13	53	14	54
rect	13	54	14	55
rect	13	56	14	57
rect	13	57	14	58
rect	13	59	14	60
rect	13	60	14	61
rect	13	62	14	63
rect	13	63	14	64
rect	13	65	14	66
rect	13	66	14	67
rect	13	68	14	69
rect	13	69	14	70
rect	13	71	14	72
rect	13	72	14	73
rect	13	74	14	75
rect	13	75	14	76
rect	13	77	14	78
rect	13	78	14	79
rect	13	80	14	81
rect	13	81	14	82
rect	13	83	14	84
rect	13	84	14	85
rect	13	86	14	87
rect	13	87	14	88
rect	13	89	14	90
rect	13	90	14	91
rect	13	92	14	93
rect	13	93	14	94
rect	13	95	14	96
rect	13	96	14	97
rect	13	98	14	99
rect	13	99	14	100
rect	13	101	14	102
rect	13	102	14	103
rect	13	104	14	105
rect	13	105	14	106
rect	13	107	14	108
rect	13	108	14	109
rect	13	110	14	111
rect	13	111	14	112
rect	13	113	14	114
rect	13	114	14	115
rect	13	116	14	117
rect	13	117	14	118
rect	13	119	14	120
rect	13	120	14	121
rect	13	122	14	123
rect	13	123	14	124
rect	13	125	14	126
rect	13	126	14	127
rect	13	128	14	129
rect	13	129	14	130
rect	13	131	14	132
rect	13	132	14	133
rect	13	134	14	135
rect	13	135	14	136
rect	13	137	14	138
rect	13	138	14	139
rect	13	140	14	141
rect	13	141	14	142
rect	13	143	14	144
rect	13	144	14	145
rect	13	146	14	147
rect	13	147	14	148
rect	13	149	14	150
rect	13	150	14	151
rect	13	152	14	153
rect	13	153	14	154
rect	13	155	14	156
rect	13	156	14	157
rect	13	158	14	159
rect	13	159	14	160
rect	13	161	14	162
rect	13	162	14	163
rect	13	164	14	165
rect	13	165	14	166
rect	13	167	14	168
rect	13	168	14	169
rect	13	170	14	171
rect	13	171	14	172
rect	13	173	14	174
rect	13	174	14	175
rect	13	176	14	177
rect	13	177	14	178
rect	13	179	14	180
rect	13	180	14	181
rect	13	182	14	183
rect	13	183	14	184
rect	13	185	14	186
rect	13	186	14	187
rect	13	188	14	189
rect	13	189	14	190
rect	13	191	14	192
rect	13	192	14	193
rect	13	194	14	195
rect	13	195	14	196
rect	13	197	14	198
rect	13	198	14	199
rect	13	200	14	201
rect	13	201	14	202
rect	13	203	14	204
rect	13	204	14	205
rect	13	206	14	207
rect	13	207	14	208
rect	13	209	14	210
rect	13	210	14	211
rect	13	212	14	213
rect	13	213	14	214
rect	13	215	14	216
rect	14	0	15	1
rect	14	2	15	3
rect	14	3	15	4
rect	14	5	15	6
rect	14	6	15	7
rect	14	8	15	9
rect	14	9	15	10
rect	14	11	15	12
rect	14	12	15	13
rect	14	14	15	15
rect	14	15	15	16
rect	14	17	15	18
rect	14	18	15	19
rect	14	20	15	21
rect	14	21	15	22
rect	14	23	15	24
rect	14	24	15	25
rect	14	26	15	27
rect	14	27	15	28
rect	14	29	15	30
rect	14	30	15	31
rect	14	32	15	33
rect	14	33	15	34
rect	14	35	15	36
rect	14	36	15	37
rect	14	38	15	39
rect	14	39	15	40
rect	14	41	15	42
rect	14	42	15	43
rect	14	44	15	45
rect	14	45	15	46
rect	14	47	15	48
rect	14	48	15	49
rect	14	50	15	51
rect	14	51	15	52
rect	14	53	15	54
rect	14	54	15	55
rect	14	56	15	57
rect	14	57	15	58
rect	14	59	15	60
rect	14	60	15	61
rect	14	62	15	63
rect	14	63	15	64
rect	14	65	15	66
rect	14	66	15	67
rect	14	68	15	69
rect	14	69	15	70
rect	14	71	15	72
rect	14	72	15	73
rect	14	74	15	75
rect	14	75	15	76
rect	14	77	15	78
rect	14	78	15	79
rect	14	80	15	81
rect	14	81	15	82
rect	14	83	15	84
rect	14	84	15	85
rect	14	86	15	87
rect	14	87	15	88
rect	14	89	15	90
rect	14	90	15	91
rect	14	92	15	93
rect	14	93	15	94
rect	14	95	15	96
rect	14	96	15	97
rect	14	98	15	99
rect	14	99	15	100
rect	14	101	15	102
rect	14	102	15	103
rect	14	104	15	105
rect	14	105	15	106
rect	14	107	15	108
rect	14	108	15	109
rect	14	110	15	111
rect	14	111	15	112
rect	14	113	15	114
rect	14	114	15	115
rect	14	116	15	117
rect	14	117	15	118
rect	14	119	15	120
rect	14	120	15	121
rect	14	122	15	123
rect	14	123	15	124
rect	14	125	15	126
rect	14	126	15	127
rect	14	128	15	129
rect	14	129	15	130
rect	14	131	15	132
rect	14	132	15	133
rect	14	134	15	135
rect	14	135	15	136
rect	14	137	15	138
rect	14	138	15	139
rect	14	140	15	141
rect	14	141	15	142
rect	14	143	15	144
rect	14	144	15	145
rect	14	146	15	147
rect	14	147	15	148
rect	14	149	15	150
rect	14	150	15	151
rect	14	152	15	153
rect	14	153	15	154
rect	14	155	15	156
rect	14	156	15	157
rect	14	158	15	159
rect	14	159	15	160
rect	14	161	15	162
rect	14	162	15	163
rect	14	164	15	165
rect	14	165	15	166
rect	14	167	15	168
rect	14	168	15	169
rect	14	170	15	171
rect	14	171	15	172
rect	14	173	15	174
rect	14	174	15	175
rect	14	176	15	177
rect	14	177	15	178
rect	14	179	15	180
rect	14	180	15	181
rect	14	182	15	183
rect	14	183	15	184
rect	14	185	15	186
rect	14	186	15	187
rect	14	188	15	189
rect	14	189	15	190
rect	14	191	15	192
rect	14	192	15	193
rect	14	194	15	195
rect	14	195	15	196
rect	14	197	15	198
rect	14	198	15	199
rect	14	200	15	201
rect	14	201	15	202
rect	14	203	15	204
rect	14	204	15	205
rect	14	206	15	207
rect	14	207	15	208
rect	14	209	15	210
rect	14	210	15	211
rect	14	212	15	213
rect	14	213	15	214
rect	14	215	15	216
rect	15	0	16	1
rect	15	2	16	3
rect	15	3	16	4
rect	15	5	16	6
rect	15	6	16	7
rect	15	8	16	9
rect	15	9	16	10
rect	15	11	16	12
rect	15	12	16	13
rect	15	14	16	15
rect	15	15	16	16
rect	15	17	16	18
rect	15	18	16	19
rect	15	20	16	21
rect	15	21	16	22
rect	15	23	16	24
rect	15	24	16	25
rect	15	26	16	27
rect	15	27	16	28
rect	15	29	16	30
rect	15	30	16	31
rect	15	32	16	33
rect	15	33	16	34
rect	15	35	16	36
rect	15	36	16	37
rect	15	38	16	39
rect	15	39	16	40
rect	15	41	16	42
rect	15	42	16	43
rect	15	44	16	45
rect	15	45	16	46
rect	15	47	16	48
rect	15	48	16	49
rect	15	50	16	51
rect	15	51	16	52
rect	15	53	16	54
rect	15	54	16	55
rect	15	56	16	57
rect	15	57	16	58
rect	15	59	16	60
rect	15	60	16	61
rect	15	62	16	63
rect	15	63	16	64
rect	15	65	16	66
rect	15	66	16	67
rect	15	68	16	69
rect	15	69	16	70
rect	15	71	16	72
rect	15	72	16	73
rect	15	74	16	75
rect	15	75	16	76
rect	15	77	16	78
rect	15	78	16	79
rect	15	80	16	81
rect	15	81	16	82
rect	15	83	16	84
rect	15	84	16	85
rect	15	86	16	87
rect	15	87	16	88
rect	15	89	16	90
rect	15	90	16	91
rect	15	92	16	93
rect	15	93	16	94
rect	15	95	16	96
rect	15	96	16	97
rect	15	98	16	99
rect	15	99	16	100
rect	15	101	16	102
rect	15	102	16	103
rect	15	104	16	105
rect	15	105	16	106
rect	15	107	16	108
rect	15	108	16	109
rect	15	110	16	111
rect	15	111	16	112
rect	15	113	16	114
rect	15	114	16	115
rect	15	116	16	117
rect	15	117	16	118
rect	15	119	16	120
rect	15	120	16	121
rect	15	122	16	123
rect	15	123	16	124
rect	15	125	16	126
rect	15	126	16	127
rect	15	128	16	129
rect	15	129	16	130
rect	15	131	16	132
rect	15	132	16	133
rect	15	134	16	135
rect	15	135	16	136
rect	15	137	16	138
rect	15	138	16	139
rect	15	140	16	141
rect	15	141	16	142
rect	15	143	16	144
rect	15	144	16	145
rect	15	146	16	147
rect	15	147	16	148
rect	15	149	16	150
rect	15	150	16	151
rect	15	152	16	153
rect	15	153	16	154
rect	15	155	16	156
rect	15	156	16	157
rect	15	158	16	159
rect	15	159	16	160
rect	15	161	16	162
rect	15	162	16	163
rect	15	164	16	165
rect	15	165	16	166
rect	15	167	16	168
rect	15	168	16	169
rect	15	170	16	171
rect	15	171	16	172
rect	15	173	16	174
rect	15	174	16	175
rect	15	176	16	177
rect	15	177	16	178
rect	15	179	16	180
rect	15	180	16	181
rect	15	182	16	183
rect	15	183	16	184
rect	15	185	16	186
rect	15	186	16	187
rect	15	188	16	189
rect	15	189	16	190
rect	15	191	16	192
rect	15	192	16	193
rect	15	194	16	195
rect	15	195	16	196
rect	15	197	16	198
rect	15	198	16	199
rect	15	200	16	201
rect	15	201	16	202
rect	15	203	16	204
rect	15	204	16	205
rect	15	206	16	207
rect	15	207	16	208
rect	15	209	16	210
rect	15	210	16	211
rect	15	212	16	213
rect	15	213	16	214
rect	15	215	16	216
rect	16	0	17	1
rect	16	2	17	3
rect	16	3	17	4
rect	16	5	17	6
rect	16	6	17	7
rect	16	8	17	9
rect	16	9	17	10
rect	16	11	17	12
rect	16	12	17	13
rect	16	14	17	15
rect	16	15	17	16
rect	16	17	17	18
rect	16	18	17	19
rect	16	20	17	21
rect	16	21	17	22
rect	16	23	17	24
rect	16	24	17	25
rect	16	26	17	27
rect	16	27	17	28
rect	16	29	17	30
rect	16	30	17	31
rect	16	32	17	33
rect	16	33	17	34
rect	16	35	17	36
rect	16	36	17	37
rect	16	38	17	39
rect	16	39	17	40
rect	16	41	17	42
rect	16	42	17	43
rect	16	44	17	45
rect	16	45	17	46
rect	16	47	17	48
rect	16	48	17	49
rect	16	50	17	51
rect	16	51	17	52
rect	16	53	17	54
rect	16	54	17	55
rect	16	56	17	57
rect	16	57	17	58
rect	16	59	17	60
rect	16	60	17	61
rect	16	62	17	63
rect	16	63	17	64
rect	16	65	17	66
rect	16	66	17	67
rect	16	68	17	69
rect	16	69	17	70
rect	16	71	17	72
rect	16	72	17	73
rect	16	74	17	75
rect	16	75	17	76
rect	16	77	17	78
rect	16	78	17	79
rect	16	80	17	81
rect	16	81	17	82
rect	16	83	17	84
rect	16	84	17	85
rect	16	86	17	87
rect	16	87	17	88
rect	16	89	17	90
rect	16	90	17	91
rect	16	92	17	93
rect	16	93	17	94
rect	16	95	17	96
rect	16	96	17	97
rect	16	98	17	99
rect	16	99	17	100
rect	16	101	17	102
rect	16	102	17	103
rect	16	104	17	105
rect	16	105	17	106
rect	16	107	17	108
rect	16	108	17	109
rect	16	110	17	111
rect	16	111	17	112
rect	16	113	17	114
rect	16	114	17	115
rect	16	116	17	117
rect	16	117	17	118
rect	16	119	17	120
rect	16	120	17	121
rect	16	122	17	123
rect	16	123	17	124
rect	16	125	17	126
rect	16	126	17	127
rect	16	128	17	129
rect	16	129	17	130
rect	16	131	17	132
rect	16	132	17	133
rect	16	134	17	135
rect	16	135	17	136
rect	16	137	17	138
rect	16	138	17	139
rect	16	140	17	141
rect	16	141	17	142
rect	16	143	17	144
rect	16	144	17	145
rect	16	146	17	147
rect	16	147	17	148
rect	16	149	17	150
rect	16	150	17	151
rect	16	152	17	153
rect	16	153	17	154
rect	16	155	17	156
rect	16	156	17	157
rect	16	158	17	159
rect	16	159	17	160
rect	16	161	17	162
rect	16	162	17	163
rect	16	164	17	165
rect	16	165	17	166
rect	16	167	17	168
rect	16	168	17	169
rect	16	170	17	171
rect	16	171	17	172
rect	16	173	17	174
rect	16	174	17	175
rect	16	176	17	177
rect	16	177	17	178
rect	16	179	17	180
rect	16	180	17	181
rect	16	182	17	183
rect	16	183	17	184
rect	16	185	17	186
rect	16	186	17	187
rect	16	188	17	189
rect	16	189	17	190
rect	16	191	17	192
rect	16	192	17	193
rect	16	194	17	195
rect	16	195	17	196
rect	16	197	17	198
rect	16	198	17	199
rect	16	200	17	201
rect	16	201	17	202
rect	16	203	17	204
rect	16	204	17	205
rect	16	206	17	207
rect	16	207	17	208
rect	16	209	17	210
rect	16	210	17	211
rect	16	212	17	213
rect	16	213	17	214
rect	16	215	17	216
rect	17	0	18	1
rect	17	2	18	3
rect	17	3	18	4
rect	17	5	18	6
rect	17	6	18	7
rect	17	8	18	9
rect	17	9	18	10
rect	17	11	18	12
rect	17	12	18	13
rect	17	14	18	15
rect	17	15	18	16
rect	17	17	18	18
rect	17	18	18	19
rect	17	20	18	21
rect	17	21	18	22
rect	17	23	18	24
rect	17	24	18	25
rect	17	26	18	27
rect	17	27	18	28
rect	17	29	18	30
rect	17	30	18	31
rect	17	32	18	33
rect	17	33	18	34
rect	17	35	18	36
rect	17	36	18	37
rect	17	38	18	39
rect	17	39	18	40
rect	17	41	18	42
rect	17	42	18	43
rect	17	44	18	45
rect	17	45	18	46
rect	17	47	18	48
rect	17	48	18	49
rect	17	50	18	51
rect	17	51	18	52
rect	17	53	18	54
rect	17	54	18	55
rect	17	56	18	57
rect	17	57	18	58
rect	17	59	18	60
rect	17	60	18	61
rect	17	62	18	63
rect	17	63	18	64
rect	17	65	18	66
rect	17	66	18	67
rect	17	68	18	69
rect	17	69	18	70
rect	17	71	18	72
rect	17	72	18	73
rect	17	74	18	75
rect	17	75	18	76
rect	17	77	18	78
rect	17	78	18	79
rect	17	80	18	81
rect	17	81	18	82
rect	17	83	18	84
rect	17	84	18	85
rect	17	86	18	87
rect	17	87	18	88
rect	17	89	18	90
rect	17	90	18	91
rect	17	92	18	93
rect	17	93	18	94
rect	17	95	18	96
rect	17	96	18	97
rect	17	98	18	99
rect	17	99	18	100
rect	17	101	18	102
rect	17	102	18	103
rect	17	104	18	105
rect	17	105	18	106
rect	17	107	18	108
rect	17	108	18	109
rect	17	110	18	111
rect	17	111	18	112
rect	17	113	18	114
rect	17	114	18	115
rect	17	116	18	117
rect	17	117	18	118
rect	17	119	18	120
rect	17	120	18	121
rect	17	122	18	123
rect	17	123	18	124
rect	17	125	18	126
rect	17	126	18	127
rect	17	128	18	129
rect	17	129	18	130
rect	17	131	18	132
rect	17	132	18	133
rect	17	134	18	135
rect	17	135	18	136
rect	17	137	18	138
rect	17	138	18	139
rect	17	140	18	141
rect	17	141	18	142
rect	17	143	18	144
rect	17	144	18	145
rect	17	146	18	147
rect	17	147	18	148
rect	17	149	18	150
rect	17	150	18	151
rect	17	152	18	153
rect	17	153	18	154
rect	17	155	18	156
rect	17	156	18	157
rect	17	158	18	159
rect	17	159	18	160
rect	17	161	18	162
rect	17	162	18	163
rect	17	164	18	165
rect	17	165	18	166
rect	17	167	18	168
rect	17	168	18	169
rect	17	170	18	171
rect	17	171	18	172
rect	17	173	18	174
rect	17	174	18	175
rect	17	176	18	177
rect	17	177	18	178
rect	17	179	18	180
rect	17	180	18	181
rect	17	182	18	183
rect	17	183	18	184
rect	17	185	18	186
rect	17	186	18	187
rect	17	188	18	189
rect	17	189	18	190
rect	17	191	18	192
rect	17	192	18	193
rect	17	194	18	195
rect	17	195	18	196
rect	17	197	18	198
rect	17	198	18	199
rect	17	200	18	201
rect	17	201	18	202
rect	17	203	18	204
rect	17	204	18	205
rect	17	206	18	207
rect	17	207	18	208
rect	17	209	18	210
rect	17	210	18	211
rect	17	212	18	213
rect	17	213	18	214
rect	17	215	18	216
rect	22	0	23	1
rect	22	2	23	3
rect	22	3	23	4
rect	22	5	23	6
rect	22	6	23	7
rect	22	8	23	9
rect	22	9	23	10
rect	22	11	23	12
rect	22	12	23	13
rect	22	14	23	15
rect	22	15	23	16
rect	22	17	23	18
rect	22	18	23	19
rect	22	20	23	21
rect	22	21	23	22
rect	22	23	23	24
rect	22	24	23	25
rect	22	26	23	27
rect	22	27	23	28
rect	22	29	23	30
rect	22	30	23	31
rect	22	32	23	33
rect	22	33	23	34
rect	22	35	23	36
rect	22	36	23	37
rect	22	38	23	39
rect	22	39	23	40
rect	22	41	23	42
rect	22	42	23	43
rect	22	44	23	45
rect	22	45	23	46
rect	22	47	23	48
rect	22	48	23	49
rect	22	50	23	51
rect	22	51	23	52
rect	22	53	23	54
rect	22	54	23	55
rect	22	56	23	57
rect	22	57	23	58
rect	22	59	23	60
rect	22	60	23	61
rect	22	62	23	63
rect	22	63	23	64
rect	22	65	23	66
rect	22	66	23	67
rect	22	68	23	69
rect	22	69	23	70
rect	22	71	23	72
rect	22	72	23	73
rect	22	74	23	75
rect	22	75	23	76
rect	22	77	23	78
rect	22	78	23	79
rect	22	80	23	81
rect	22	81	23	82
rect	22	83	23	84
rect	22	84	23	85
rect	22	86	23	87
rect	22	87	23	88
rect	22	89	23	90
rect	22	90	23	91
rect	22	92	23	93
rect	22	93	23	94
rect	22	95	23	96
rect	22	96	23	97
rect	22	98	23	99
rect	22	99	23	100
rect	22	101	23	102
rect	22	102	23	103
rect	22	104	23	105
rect	22	105	23	106
rect	22	107	23	108
rect	22	108	23	109
rect	22	110	23	111
rect	22	111	23	112
rect	22	113	23	114
rect	22	114	23	115
rect	22	116	23	117
rect	22	117	23	118
rect	22	119	23	120
rect	22	120	23	121
rect	22	122	23	123
rect	22	123	23	124
rect	22	125	23	126
rect	22	126	23	127
rect	22	128	23	129
rect	22	129	23	130
rect	22	131	23	132
rect	22	132	23	133
rect	22	134	23	135
rect	22	135	23	136
rect	22	137	23	138
rect	22	138	23	139
rect	22	140	23	141
rect	22	141	23	142
rect	22	143	23	144
rect	22	144	23	145
rect	22	146	23	147
rect	22	147	23	148
rect	22	149	23	150
rect	22	150	23	151
rect	22	152	23	153
rect	22	153	23	154
rect	22	155	23	156
rect	22	156	23	157
rect	22	158	23	159
rect	22	159	23	160
rect	22	161	23	162
rect	22	162	23	163
rect	22	164	23	165
rect	22	165	23	166
rect	22	167	23	168
rect	22	168	23	169
rect	22	170	23	171
rect	22	171	23	172
rect	22	173	23	174
rect	22	174	23	175
rect	22	176	23	177
rect	22	177	23	178
rect	22	179	23	180
rect	22	180	23	181
rect	22	182	23	183
rect	22	183	23	184
rect	22	185	23	186
rect	22	186	23	187
rect	22	188	23	189
rect	22	189	23	190
rect	22	191	23	192
rect	22	192	23	193
rect	22	194	23	195
rect	22	195	23	196
rect	22	197	23	198
rect	22	198	23	199
rect	22	200	23	201
rect	22	201	23	202
rect	22	203	23	204
rect	22	204	23	205
rect	22	206	23	207
rect	22	207	23	208
rect	22	209	23	210
rect	22	210	23	211
rect	22	212	23	213
rect	22	213	23	214
rect	22	215	23	216
rect	24	0	25	1
rect	24	2	25	3
rect	24	3	25	4
rect	24	5	25	6
rect	24	6	25	7
rect	24	8	25	9
rect	24	9	25	10
rect	24	11	25	12
rect	24	12	25	13
rect	24	14	25	15
rect	24	15	25	16
rect	24	17	25	18
rect	24	18	25	19
rect	24	20	25	21
rect	24	21	25	22
rect	24	23	25	24
rect	24	24	25	25
rect	24	26	25	27
rect	24	27	25	28
rect	24	29	25	30
rect	24	30	25	31
rect	24	32	25	33
rect	24	33	25	34
rect	24	35	25	36
rect	24	36	25	37
rect	24	38	25	39
rect	24	39	25	40
rect	24	41	25	42
rect	24	42	25	43
rect	24	44	25	45
rect	24	45	25	46
rect	24	47	25	48
rect	24	48	25	49
rect	24	50	25	51
rect	24	51	25	52
rect	24	53	25	54
rect	24	54	25	55
rect	24	56	25	57
rect	24	57	25	58
rect	24	59	25	60
rect	24	60	25	61
rect	24	62	25	63
rect	24	63	25	64
rect	24	65	25	66
rect	24	66	25	67
rect	24	68	25	69
rect	24	69	25	70
rect	24	71	25	72
rect	24	72	25	73
rect	24	74	25	75
rect	24	75	25	76
rect	24	77	25	78
rect	24	78	25	79
rect	24	80	25	81
rect	24	81	25	82
rect	24	83	25	84
rect	24	84	25	85
rect	24	86	25	87
rect	24	87	25	88
rect	24	89	25	90
rect	24	90	25	91
rect	24	92	25	93
rect	24	93	25	94
rect	24	95	25	96
rect	24	96	25	97
rect	24	98	25	99
rect	24	99	25	100
rect	24	101	25	102
rect	24	102	25	103
rect	24	104	25	105
rect	24	105	25	106
rect	24	107	25	108
rect	24	108	25	109
rect	24	110	25	111
rect	24	111	25	112
rect	24	113	25	114
rect	24	114	25	115
rect	24	116	25	117
rect	24	117	25	118
rect	24	119	25	120
rect	24	120	25	121
rect	24	122	25	123
rect	24	123	25	124
rect	24	125	25	126
rect	24	126	25	127
rect	24	128	25	129
rect	24	129	25	130
rect	24	131	25	132
rect	24	132	25	133
rect	24	134	25	135
rect	24	135	25	136
rect	24	137	25	138
rect	24	138	25	139
rect	24	140	25	141
rect	24	141	25	142
rect	24	143	25	144
rect	24	144	25	145
rect	24	146	25	147
rect	24	147	25	148
rect	24	149	25	150
rect	24	150	25	151
rect	24	152	25	153
rect	24	153	25	154
rect	24	155	25	156
rect	24	156	25	157
rect	24	158	25	159
rect	24	159	25	160
rect	24	161	25	162
rect	24	162	25	163
rect	24	164	25	165
rect	24	165	25	166
rect	24	167	25	168
rect	24	168	25	169
rect	24	170	25	171
rect	24	171	25	172
rect	24	173	25	174
rect	24	174	25	175
rect	24	176	25	177
rect	24	177	25	178
rect	24	179	25	180
rect	24	180	25	181
rect	24	182	25	183
rect	24	183	25	184
rect	24	185	25	186
rect	24	186	25	187
rect	24	188	25	189
rect	24	189	25	190
rect	24	191	25	192
rect	24	192	25	193
rect	24	194	25	195
rect	24	195	25	196
rect	24	197	25	198
rect	24	198	25	199
rect	24	200	25	201
rect	24	201	25	202
rect	24	203	25	204
rect	24	204	25	205
rect	24	206	25	207
rect	24	207	25	208
rect	24	209	25	210
rect	24	210	25	211
rect	24	212	25	213
rect	24	213	25	214
rect	24	215	25	216
rect	24	216	25	217
rect	24	218	25	219
rect	24	219	25	220
rect	24	221	25	222
rect	24	222	25	223
rect	24	224	25	225
rect	24	225	25	226
rect	24	227	25	228
rect	24	228	25	229
rect	24	230	25	231
rect	24	231	25	232
rect	24	233	25	234
rect	24	234	25	235
rect	24	236	25	237
rect	24	237	25	238
rect	24	239	25	240
rect	24	240	25	241
rect	24	242	25	243
rect	25	0	26	1
rect	25	2	26	3
rect	25	3	26	4
rect	25	5	26	6
rect	25	6	26	7
rect	25	8	26	9
rect	25	9	26	10
rect	25	11	26	12
rect	25	12	26	13
rect	25	14	26	15
rect	25	15	26	16
rect	25	17	26	18
rect	25	18	26	19
rect	25	20	26	21
rect	25	21	26	22
rect	25	23	26	24
rect	25	24	26	25
rect	25	26	26	27
rect	25	27	26	28
rect	25	29	26	30
rect	25	30	26	31
rect	25	32	26	33
rect	25	33	26	34
rect	25	35	26	36
rect	25	36	26	37
rect	25	38	26	39
rect	25	39	26	40
rect	25	41	26	42
rect	25	42	26	43
rect	25	44	26	45
rect	25	45	26	46
rect	25	47	26	48
rect	25	48	26	49
rect	25	50	26	51
rect	25	51	26	52
rect	25	53	26	54
rect	25	54	26	55
rect	25	56	26	57
rect	25	57	26	58
rect	25	59	26	60
rect	25	60	26	61
rect	25	62	26	63
rect	25	63	26	64
rect	25	65	26	66
rect	25	66	26	67
rect	25	68	26	69
rect	25	69	26	70
rect	25	71	26	72
rect	25	72	26	73
rect	25	74	26	75
rect	25	75	26	76
rect	25	77	26	78
rect	25	78	26	79
rect	25	80	26	81
rect	25	81	26	82
rect	25	83	26	84
rect	25	84	26	85
rect	25	86	26	87
rect	25	87	26	88
rect	25	89	26	90
rect	25	90	26	91
rect	25	92	26	93
rect	25	93	26	94
rect	25	95	26	96
rect	25	96	26	97
rect	25	98	26	99
rect	25	99	26	100
rect	25	101	26	102
rect	25	102	26	103
rect	25	104	26	105
rect	25	105	26	106
rect	25	107	26	108
rect	25	108	26	109
rect	25	110	26	111
rect	25	111	26	112
rect	25	113	26	114
rect	25	114	26	115
rect	25	116	26	117
rect	25	117	26	118
rect	25	119	26	120
rect	25	120	26	121
rect	25	122	26	123
rect	25	123	26	124
rect	25	125	26	126
rect	25	126	26	127
rect	25	128	26	129
rect	25	129	26	130
rect	25	131	26	132
rect	25	132	26	133
rect	25	134	26	135
rect	25	135	26	136
rect	25	137	26	138
rect	25	138	26	139
rect	25	140	26	141
rect	25	141	26	142
rect	25	143	26	144
rect	25	144	26	145
rect	25	146	26	147
rect	25	147	26	148
rect	25	149	26	150
rect	25	150	26	151
rect	25	152	26	153
rect	25	153	26	154
rect	25	155	26	156
rect	25	156	26	157
rect	25	158	26	159
rect	25	159	26	160
rect	25	161	26	162
rect	25	162	26	163
rect	25	164	26	165
rect	25	165	26	166
rect	25	167	26	168
rect	25	168	26	169
rect	25	170	26	171
rect	25	171	26	172
rect	25	173	26	174
rect	25	174	26	175
rect	25	176	26	177
rect	25	177	26	178
rect	25	179	26	180
rect	25	180	26	181
rect	25	182	26	183
rect	25	183	26	184
rect	25	185	26	186
rect	25	186	26	187
rect	25	188	26	189
rect	25	189	26	190
rect	25	191	26	192
rect	25	192	26	193
rect	25	194	26	195
rect	25	195	26	196
rect	25	197	26	198
rect	25	198	26	199
rect	25	200	26	201
rect	25	201	26	202
rect	25	203	26	204
rect	25	204	26	205
rect	25	206	26	207
rect	25	207	26	208
rect	25	209	26	210
rect	25	210	26	211
rect	25	212	26	213
rect	25	213	26	214
rect	25	215	26	216
rect	25	216	26	217
rect	25	218	26	219
rect	25	219	26	220
rect	25	221	26	222
rect	25	222	26	223
rect	25	224	26	225
rect	25	225	26	226
rect	25	227	26	228
rect	25	228	26	229
rect	25	230	26	231
rect	25	231	26	232
rect	25	233	26	234
rect	25	234	26	235
rect	25	236	26	237
rect	25	237	26	238
rect	25	239	26	240
rect	25	240	26	241
rect	25	242	26	243
rect	26	0	27	1
rect	26	2	27	3
rect	26	3	27	4
rect	26	5	27	6
rect	26	6	27	7
rect	26	8	27	9
rect	26	9	27	10
rect	26	11	27	12
rect	26	12	27	13
rect	26	14	27	15
rect	26	15	27	16
rect	26	17	27	18
rect	26	18	27	19
rect	26	20	27	21
rect	26	21	27	22
rect	26	23	27	24
rect	26	24	27	25
rect	26	26	27	27
rect	26	27	27	28
rect	26	29	27	30
rect	26	30	27	31
rect	26	32	27	33
rect	26	33	27	34
rect	26	35	27	36
rect	26	36	27	37
rect	26	38	27	39
rect	26	39	27	40
rect	26	41	27	42
rect	26	42	27	43
rect	26	44	27	45
rect	26	45	27	46
rect	26	47	27	48
rect	26	48	27	49
rect	26	50	27	51
rect	26	51	27	52
rect	26	53	27	54
rect	26	54	27	55
rect	26	56	27	57
rect	26	57	27	58
rect	26	59	27	60
rect	26	60	27	61
rect	26	62	27	63
rect	26	63	27	64
rect	26	65	27	66
rect	26	66	27	67
rect	26	68	27	69
rect	26	69	27	70
rect	26	71	27	72
rect	26	72	27	73
rect	26	74	27	75
rect	26	75	27	76
rect	26	77	27	78
rect	26	78	27	79
rect	26	80	27	81
rect	26	81	27	82
rect	26	83	27	84
rect	26	84	27	85
rect	26	86	27	87
rect	26	87	27	88
rect	26	89	27	90
rect	26	90	27	91
rect	26	92	27	93
rect	26	93	27	94
rect	26	95	27	96
rect	26	96	27	97
rect	26	98	27	99
rect	26	99	27	100
rect	26	101	27	102
rect	26	102	27	103
rect	26	104	27	105
rect	26	105	27	106
rect	26	107	27	108
rect	26	108	27	109
rect	26	110	27	111
rect	26	111	27	112
rect	26	113	27	114
rect	26	114	27	115
rect	26	116	27	117
rect	26	117	27	118
rect	26	119	27	120
rect	26	120	27	121
rect	26	122	27	123
rect	26	123	27	124
rect	26	125	27	126
rect	26	126	27	127
rect	26	128	27	129
rect	26	129	27	130
rect	26	131	27	132
rect	26	132	27	133
rect	26	134	27	135
rect	26	135	27	136
rect	26	137	27	138
rect	26	138	27	139
rect	26	140	27	141
rect	26	141	27	142
rect	26	143	27	144
rect	26	144	27	145
rect	26	146	27	147
rect	26	147	27	148
rect	26	149	27	150
rect	26	150	27	151
rect	26	152	27	153
rect	26	153	27	154
rect	26	155	27	156
rect	26	156	27	157
rect	26	158	27	159
rect	26	159	27	160
rect	26	161	27	162
rect	26	162	27	163
rect	26	164	27	165
rect	26	165	27	166
rect	26	167	27	168
rect	26	168	27	169
rect	26	170	27	171
rect	26	171	27	172
rect	26	173	27	174
rect	26	174	27	175
rect	26	176	27	177
rect	26	177	27	178
rect	26	179	27	180
rect	26	180	27	181
rect	26	182	27	183
rect	26	183	27	184
rect	26	185	27	186
rect	26	186	27	187
rect	26	188	27	189
rect	26	189	27	190
rect	26	191	27	192
rect	26	192	27	193
rect	26	194	27	195
rect	26	195	27	196
rect	26	197	27	198
rect	26	198	27	199
rect	26	200	27	201
rect	26	201	27	202
rect	26	203	27	204
rect	26	204	27	205
rect	26	206	27	207
rect	26	207	27	208
rect	26	209	27	210
rect	26	210	27	211
rect	26	212	27	213
rect	26	213	27	214
rect	26	215	27	216
rect	26	216	27	217
rect	26	218	27	219
rect	26	219	27	220
rect	26	221	27	222
rect	26	222	27	223
rect	26	224	27	225
rect	26	225	27	226
rect	26	227	27	228
rect	26	228	27	229
rect	26	230	27	231
rect	26	231	27	232
rect	26	233	27	234
rect	26	234	27	235
rect	26	236	27	237
rect	26	237	27	238
rect	26	239	27	240
rect	26	240	27	241
rect	26	242	27	243
rect	27	0	28	1
rect	27	2	28	3
rect	27	3	28	4
rect	27	5	28	6
rect	27	6	28	7
rect	27	8	28	9
rect	27	9	28	10
rect	27	11	28	12
rect	27	12	28	13
rect	27	14	28	15
rect	27	15	28	16
rect	27	17	28	18
rect	27	18	28	19
rect	27	20	28	21
rect	27	21	28	22
rect	27	23	28	24
rect	27	24	28	25
rect	27	26	28	27
rect	27	27	28	28
rect	27	29	28	30
rect	27	30	28	31
rect	27	32	28	33
rect	27	33	28	34
rect	27	35	28	36
rect	27	36	28	37
rect	27	38	28	39
rect	27	39	28	40
rect	27	41	28	42
rect	27	42	28	43
rect	27	44	28	45
rect	27	45	28	46
rect	27	47	28	48
rect	27	48	28	49
rect	27	50	28	51
rect	27	51	28	52
rect	27	53	28	54
rect	27	54	28	55
rect	27	56	28	57
rect	27	57	28	58
rect	27	59	28	60
rect	27	60	28	61
rect	27	62	28	63
rect	27	63	28	64
rect	27	65	28	66
rect	27	66	28	67
rect	27	68	28	69
rect	27	69	28	70
rect	27	71	28	72
rect	27	72	28	73
rect	27	74	28	75
rect	27	75	28	76
rect	27	77	28	78
rect	27	78	28	79
rect	27	80	28	81
rect	27	81	28	82
rect	27	83	28	84
rect	27	84	28	85
rect	27	86	28	87
rect	27	87	28	88
rect	27	89	28	90
rect	27	90	28	91
rect	27	92	28	93
rect	27	93	28	94
rect	27	95	28	96
rect	27	96	28	97
rect	27	98	28	99
rect	27	99	28	100
rect	27	101	28	102
rect	27	102	28	103
rect	27	104	28	105
rect	27	105	28	106
rect	27	107	28	108
rect	27	108	28	109
rect	27	110	28	111
rect	27	111	28	112
rect	27	113	28	114
rect	27	114	28	115
rect	27	116	28	117
rect	27	117	28	118
rect	27	119	28	120
rect	27	120	28	121
rect	27	122	28	123
rect	27	123	28	124
rect	27	125	28	126
rect	27	126	28	127
rect	27	128	28	129
rect	27	129	28	130
rect	27	131	28	132
rect	27	132	28	133
rect	27	134	28	135
rect	27	135	28	136
rect	27	137	28	138
rect	27	138	28	139
rect	27	140	28	141
rect	27	141	28	142
rect	27	143	28	144
rect	27	144	28	145
rect	27	146	28	147
rect	27	147	28	148
rect	27	149	28	150
rect	27	150	28	151
rect	27	152	28	153
rect	27	153	28	154
rect	27	155	28	156
rect	27	156	28	157
rect	27	158	28	159
rect	27	159	28	160
rect	27	161	28	162
rect	27	162	28	163
rect	27	164	28	165
rect	27	165	28	166
rect	27	167	28	168
rect	27	168	28	169
rect	27	170	28	171
rect	27	171	28	172
rect	27	173	28	174
rect	27	174	28	175
rect	27	176	28	177
rect	27	177	28	178
rect	27	179	28	180
rect	27	180	28	181
rect	27	182	28	183
rect	27	183	28	184
rect	27	185	28	186
rect	27	186	28	187
rect	27	188	28	189
rect	27	189	28	190
rect	27	191	28	192
rect	27	192	28	193
rect	27	194	28	195
rect	27	195	28	196
rect	27	197	28	198
rect	27	198	28	199
rect	27	200	28	201
rect	27	201	28	202
rect	27	203	28	204
rect	27	204	28	205
rect	27	206	28	207
rect	27	207	28	208
rect	27	209	28	210
rect	27	210	28	211
rect	27	212	28	213
rect	27	213	28	214
rect	27	215	28	216
rect	27	216	28	217
rect	27	218	28	219
rect	27	219	28	220
rect	27	221	28	222
rect	27	222	28	223
rect	27	224	28	225
rect	27	225	28	226
rect	27	227	28	228
rect	27	228	28	229
rect	27	230	28	231
rect	27	231	28	232
rect	27	233	28	234
rect	27	234	28	235
rect	27	236	28	237
rect	27	237	28	238
rect	27	239	28	240
rect	27	240	28	241
rect	27	242	28	243
rect	28	0	29	1
rect	28	2	29	3
rect	28	3	29	4
rect	28	5	29	6
rect	28	6	29	7
rect	28	8	29	9
rect	28	9	29	10
rect	28	11	29	12
rect	28	12	29	13
rect	28	14	29	15
rect	28	15	29	16
rect	28	17	29	18
rect	28	18	29	19
rect	28	20	29	21
rect	28	21	29	22
rect	28	23	29	24
rect	28	24	29	25
rect	28	26	29	27
rect	28	27	29	28
rect	28	29	29	30
rect	28	30	29	31
rect	28	32	29	33
rect	28	33	29	34
rect	28	35	29	36
rect	28	36	29	37
rect	28	38	29	39
rect	28	39	29	40
rect	28	41	29	42
rect	28	42	29	43
rect	28	44	29	45
rect	28	45	29	46
rect	28	47	29	48
rect	28	48	29	49
rect	28	50	29	51
rect	28	51	29	52
rect	28	53	29	54
rect	28	54	29	55
rect	28	56	29	57
rect	28	57	29	58
rect	28	59	29	60
rect	28	60	29	61
rect	28	62	29	63
rect	28	63	29	64
rect	28	65	29	66
rect	28	66	29	67
rect	28	68	29	69
rect	28	69	29	70
rect	28	71	29	72
rect	28	72	29	73
rect	28	74	29	75
rect	28	75	29	76
rect	28	77	29	78
rect	28	78	29	79
rect	28	80	29	81
rect	28	81	29	82
rect	28	83	29	84
rect	28	84	29	85
rect	28	86	29	87
rect	28	87	29	88
rect	28	89	29	90
rect	28	90	29	91
rect	28	92	29	93
rect	28	93	29	94
rect	28	95	29	96
rect	28	96	29	97
rect	28	98	29	99
rect	28	99	29	100
rect	28	101	29	102
rect	28	102	29	103
rect	28	104	29	105
rect	28	105	29	106
rect	28	107	29	108
rect	28	108	29	109
rect	28	110	29	111
rect	28	111	29	112
rect	28	113	29	114
rect	28	114	29	115
rect	28	116	29	117
rect	28	117	29	118
rect	28	119	29	120
rect	28	120	29	121
rect	28	122	29	123
rect	28	123	29	124
rect	28	125	29	126
rect	28	126	29	127
rect	28	128	29	129
rect	28	129	29	130
rect	28	131	29	132
rect	28	132	29	133
rect	28	134	29	135
rect	28	135	29	136
rect	28	137	29	138
rect	28	138	29	139
rect	28	140	29	141
rect	28	141	29	142
rect	28	143	29	144
rect	28	144	29	145
rect	28	146	29	147
rect	28	147	29	148
rect	28	149	29	150
rect	28	150	29	151
rect	28	152	29	153
rect	28	153	29	154
rect	28	155	29	156
rect	28	156	29	157
rect	28	158	29	159
rect	28	159	29	160
rect	28	161	29	162
rect	28	162	29	163
rect	28	164	29	165
rect	28	165	29	166
rect	28	167	29	168
rect	28	168	29	169
rect	28	170	29	171
rect	28	171	29	172
rect	28	173	29	174
rect	28	174	29	175
rect	28	176	29	177
rect	28	177	29	178
rect	28	179	29	180
rect	28	180	29	181
rect	28	182	29	183
rect	28	183	29	184
rect	28	185	29	186
rect	28	186	29	187
rect	28	188	29	189
rect	28	189	29	190
rect	28	191	29	192
rect	28	192	29	193
rect	28	194	29	195
rect	28	195	29	196
rect	28	197	29	198
rect	28	198	29	199
rect	28	200	29	201
rect	28	201	29	202
rect	28	203	29	204
rect	28	204	29	205
rect	28	206	29	207
rect	28	207	29	208
rect	28	209	29	210
rect	28	210	29	211
rect	28	212	29	213
rect	28	213	29	214
rect	28	215	29	216
rect	28	216	29	217
rect	28	218	29	219
rect	28	219	29	220
rect	28	221	29	222
rect	28	222	29	223
rect	28	224	29	225
rect	28	225	29	226
rect	28	227	29	228
rect	28	228	29	229
rect	28	230	29	231
rect	28	231	29	232
rect	28	233	29	234
rect	28	234	29	235
rect	28	236	29	237
rect	28	237	29	238
rect	28	239	29	240
rect	28	240	29	241
rect	28	242	29	243
rect	37	0	38	1
rect	37	2	38	3
rect	37	3	38	4
rect	37	5	38	6
rect	37	6	38	7
rect	37	8	38	9
rect	37	9	38	10
rect	37	11	38	12
rect	37	12	38	13
rect	37	14	38	15
rect	37	15	38	16
rect	37	17	38	18
rect	37	18	38	19
rect	37	20	38	21
rect	37	21	38	22
rect	37	23	38	24
rect	37	24	38	25
rect	37	26	38	27
rect	37	27	38	28
rect	37	29	38	30
rect	37	30	38	31
rect	37	32	38	33
rect	37	33	38	34
rect	37	35	38	36
rect	37	36	38	37
rect	37	38	38	39
rect	37	39	38	40
rect	37	41	38	42
rect	37	42	38	43
rect	37	44	38	45
rect	37	45	38	46
rect	37	47	38	48
rect	37	48	38	49
rect	37	50	38	51
rect	37	51	38	52
rect	37	53	38	54
rect	37	54	38	55
rect	37	56	38	57
rect	37	57	38	58
rect	37	59	38	60
rect	37	60	38	61
rect	37	62	38	63
rect	37	63	38	64
rect	37	65	38	66
rect	37	66	38	67
rect	37	68	38	69
rect	37	69	38	70
rect	37	71	38	72
rect	37	72	38	73
rect	37	74	38	75
rect	37	75	38	76
rect	37	77	38	78
rect	37	78	38	79
rect	37	80	38	81
rect	37	81	38	82
rect	37	83	38	84
rect	37	84	38	85
rect	37	86	38	87
rect	37	87	38	88
rect	37	89	38	90
rect	37	90	38	91
rect	37	92	38	93
rect	37	93	38	94
rect	37	95	38	96
rect	37	96	38	97
rect	37	98	38	99
rect	37	99	38	100
rect	37	101	38	102
rect	37	102	38	103
rect	37	104	38	105
rect	37	105	38	106
rect	37	107	38	108
rect	37	108	38	109
rect	37	110	38	111
rect	37	111	38	112
rect	37	113	38	114
rect	37	114	38	115
rect	37	116	38	117
rect	37	117	38	118
rect	37	119	38	120
rect	37	120	38	121
rect	37	122	38	123
rect	37	123	38	124
rect	37	125	38	126
rect	37	126	38	127
rect	37	128	38	129
rect	37	129	38	130
rect	37	131	38	132
rect	37	132	38	133
rect	37	134	38	135
rect	37	135	38	136
rect	37	137	38	138
rect	37	138	38	139
rect	37	140	38	141
rect	37	141	38	142
rect	37	143	38	144
rect	37	144	38	145
rect	37	146	38	147
rect	37	147	38	148
rect	37	149	38	150
rect	37	150	38	151
rect	37	152	38	153
rect	37	153	38	154
rect	37	155	38	156
rect	37	156	38	157
rect	37	158	38	159
rect	37	159	38	160
rect	37	161	38	162
rect	37	162	38	163
rect	37	164	38	165
rect	37	165	38	166
rect	37	167	38	168
rect	37	168	38	169
rect	37	170	38	171
rect	37	171	38	172
rect	37	173	38	174
rect	37	174	38	175
rect	37	176	38	177
rect	37	177	38	178
rect	37	179	38	180
rect	37	180	38	181
rect	37	182	38	183
rect	37	183	38	184
rect	37	185	38	186
rect	37	186	38	187
rect	37	188	38	189
rect	37	189	38	190
rect	37	191	38	192
rect	37	192	38	193
rect	37	194	38	195
rect	37	195	38	196
rect	37	197	38	198
rect	37	198	38	199
rect	37	200	38	201
rect	37	201	38	202
rect	37	203	38	204
rect	37	204	38	205
rect	37	206	38	207
rect	37	207	38	208
rect	37	209	38	210
rect	37	210	38	211
rect	37	212	38	213
rect	37	213	38	214
rect	37	215	38	216
rect	37	216	38	217
rect	37	218	38	219
rect	37	219	38	220
rect	37	221	38	222
rect	37	222	38	223
rect	37	224	38	225
rect	37	225	38	226
rect	37	227	38	228
rect	37	228	38	229
rect	37	230	38	231
rect	37	231	38	232
rect	37	233	38	234
rect	37	234	38	235
rect	37	236	38	237
rect	37	237	38	238
rect	37	239	38	240
rect	37	240	38	241
rect	37	242	38	243
rect	39	0	40	1
rect	39	2	40	3
rect	39	3	40	4
rect	39	5	40	6
rect	39	6	40	7
rect	39	8	40	9
rect	39	9	40	10
rect	39	11	40	12
rect	39	12	40	13
rect	39	14	40	15
rect	39	15	40	16
rect	39	17	40	18
rect	39	18	40	19
rect	39	20	40	21
rect	39	21	40	22
rect	39	23	40	24
rect	39	24	40	25
rect	39	26	40	27
rect	39	27	40	28
rect	39	29	40	30
rect	39	30	40	31
rect	39	32	40	33
rect	39	33	40	34
rect	39	35	40	36
rect	39	36	40	37
rect	39	38	40	39
rect	39	39	40	40
rect	39	41	40	42
rect	39	42	40	43
rect	39	44	40	45
rect	39	45	40	46
rect	39	47	40	48
rect	39	48	40	49
rect	39	50	40	51
rect	39	51	40	52
rect	39	53	40	54
rect	39	54	40	55
rect	39	56	40	57
rect	39	57	40	58
rect	39	59	40	60
rect	39	60	40	61
rect	39	62	40	63
rect	39	63	40	64
rect	39	65	40	66
rect	39	66	40	67
rect	39	68	40	69
rect	39	69	40	70
rect	39	71	40	72
rect	39	72	40	73
rect	39	74	40	75
rect	39	75	40	76
rect	39	77	40	78
rect	39	78	40	79
rect	39	80	40	81
rect	39	81	40	82
rect	39	83	40	84
rect	39	84	40	85
rect	39	86	40	87
rect	39	87	40	88
rect	39	89	40	90
rect	39	90	40	91
rect	39	92	40	93
rect	39	93	40	94
rect	39	95	40	96
rect	39	96	40	97
rect	39	98	40	99
rect	39	99	40	100
rect	39	101	40	102
rect	39	102	40	103
rect	39	104	40	105
rect	39	105	40	106
rect	39	107	40	108
rect	39	108	40	109
rect	39	110	40	111
rect	39	111	40	112
rect	39	113	40	114
rect	39	114	40	115
rect	39	116	40	117
rect	39	117	40	118
rect	39	119	40	120
rect	39	120	40	121
rect	39	122	40	123
rect	39	123	40	124
rect	39	125	40	126
rect	39	126	40	127
rect	39	128	40	129
rect	39	129	40	130
rect	39	131	40	132
rect	39	132	40	133
rect	39	134	40	135
rect	39	135	40	136
rect	39	137	40	138
rect	39	138	40	139
rect	39	140	40	141
rect	39	141	40	142
rect	39	143	40	144
rect	39	144	40	145
rect	39	146	40	147
rect	39	147	40	148
rect	39	149	40	150
rect	39	150	40	151
rect	39	152	40	153
rect	39	153	40	154
rect	39	155	40	156
rect	39	156	40	157
rect	39	158	40	159
rect	39	159	40	160
rect	39	161	40	162
rect	39	162	40	163
rect	39	164	40	165
rect	39	165	40	166
rect	39	167	40	168
rect	39	168	40	169
rect	39	170	40	171
rect	39	171	40	172
rect	39	173	40	174
rect	39	174	40	175
rect	39	176	40	177
rect	39	177	40	178
rect	39	179	40	180
rect	39	180	40	181
rect	39	182	40	183
rect	39	183	40	184
rect	39	185	40	186
rect	39	186	40	187
rect	39	188	40	189
rect	39	189	40	190
rect	39	191	40	192
rect	39	192	40	193
rect	39	194	40	195
rect	39	195	40	196
rect	39	197	40	198
rect	39	198	40	199
rect	39	200	40	201
rect	39	201	40	202
rect	39	203	40	204
rect	39	204	40	205
rect	39	206	40	207
rect	39	207	40	208
rect	39	209	40	210
rect	39	210	40	211
rect	39	212	40	213
rect	39	213	40	214
rect	39	215	40	216
rect	39	216	40	217
rect	39	218	40	219
rect	39	219	40	220
rect	39	221	40	222
rect	39	222	40	223
rect	39	224	40	225
rect	39	225	40	226
rect	39	227	40	228
rect	39	228	40	229
rect	39	230	40	231
rect	39	231	40	232
rect	39	233	40	234
rect	39	234	40	235
rect	39	236	40	237
rect	39	237	40	238
rect	39	239	40	240
rect	39	240	40	241
rect	39	242	40	243
rect	39	243	40	244
rect	39	245	40	246
rect	39	246	40	247
rect	39	248	40	249
rect	39	249	40	250
rect	39	251	40	252
rect	39	252	40	253
rect	39	254	40	255
rect	39	255	40	256
rect	39	257	40	258
rect	39	258	40	259
rect	39	260	40	261
rect	39	261	40	262
rect	39	263	40	264
rect	39	264	40	265
rect	39	266	40	267
rect	39	267	40	268
rect	39	269	40	270
rect	39	270	40	271
rect	39	272	40	273
rect	39	273	40	274
rect	39	275	40	276
rect	39	276	40	277
rect	39	278	40	279
rect	39	279	40	280
rect	39	281	40	282
rect	39	282	40	283
rect	39	284	40	285
rect	39	285	40	286
rect	39	287	40	288
rect	39	288	40	289
rect	39	290	40	291
rect	40	0	41	1
rect	40	2	41	3
rect	40	3	41	4
rect	40	5	41	6
rect	40	6	41	7
rect	40	8	41	9
rect	40	9	41	10
rect	40	11	41	12
rect	40	12	41	13
rect	40	14	41	15
rect	40	15	41	16
rect	40	17	41	18
rect	40	18	41	19
rect	40	20	41	21
rect	40	21	41	22
rect	40	23	41	24
rect	40	24	41	25
rect	40	26	41	27
rect	40	27	41	28
rect	40	29	41	30
rect	40	30	41	31
rect	40	32	41	33
rect	40	33	41	34
rect	40	35	41	36
rect	40	36	41	37
rect	40	38	41	39
rect	40	39	41	40
rect	40	41	41	42
rect	40	42	41	43
rect	40	44	41	45
rect	40	45	41	46
rect	40	47	41	48
rect	40	48	41	49
rect	40	50	41	51
rect	40	51	41	52
rect	40	53	41	54
rect	40	54	41	55
rect	40	56	41	57
rect	40	57	41	58
rect	40	59	41	60
rect	40	60	41	61
rect	40	62	41	63
rect	40	63	41	64
rect	40	65	41	66
rect	40	66	41	67
rect	40	68	41	69
rect	40	69	41	70
rect	40	71	41	72
rect	40	72	41	73
rect	40	74	41	75
rect	40	75	41	76
rect	40	77	41	78
rect	40	78	41	79
rect	40	80	41	81
rect	40	81	41	82
rect	40	83	41	84
rect	40	84	41	85
rect	40	86	41	87
rect	40	87	41	88
rect	40	89	41	90
rect	40	90	41	91
rect	40	92	41	93
rect	40	93	41	94
rect	40	95	41	96
rect	40	96	41	97
rect	40	98	41	99
rect	40	99	41	100
rect	40	101	41	102
rect	40	102	41	103
rect	40	104	41	105
rect	40	105	41	106
rect	40	107	41	108
rect	40	108	41	109
rect	40	110	41	111
rect	40	111	41	112
rect	40	113	41	114
rect	40	114	41	115
rect	40	116	41	117
rect	40	117	41	118
rect	40	119	41	120
rect	40	120	41	121
rect	40	122	41	123
rect	40	123	41	124
rect	40	125	41	126
rect	40	126	41	127
rect	40	128	41	129
rect	40	129	41	130
rect	40	131	41	132
rect	40	132	41	133
rect	40	134	41	135
rect	40	135	41	136
rect	40	137	41	138
rect	40	138	41	139
rect	40	140	41	141
rect	40	141	41	142
rect	40	143	41	144
rect	40	144	41	145
rect	40	146	41	147
rect	40	147	41	148
rect	40	149	41	150
rect	40	150	41	151
rect	40	152	41	153
rect	40	153	41	154
rect	40	155	41	156
rect	40	156	41	157
rect	40	158	41	159
rect	40	159	41	160
rect	40	161	41	162
rect	40	162	41	163
rect	40	164	41	165
rect	40	165	41	166
rect	40	167	41	168
rect	40	168	41	169
rect	40	170	41	171
rect	40	171	41	172
rect	40	173	41	174
rect	40	174	41	175
rect	40	176	41	177
rect	40	177	41	178
rect	40	179	41	180
rect	40	180	41	181
rect	40	182	41	183
rect	40	183	41	184
rect	40	185	41	186
rect	40	186	41	187
rect	40	188	41	189
rect	40	189	41	190
rect	40	191	41	192
rect	40	192	41	193
rect	40	194	41	195
rect	40	195	41	196
rect	40	197	41	198
rect	40	198	41	199
rect	40	200	41	201
rect	40	201	41	202
rect	40	203	41	204
rect	40	204	41	205
rect	40	206	41	207
rect	40	207	41	208
rect	40	209	41	210
rect	40	210	41	211
rect	40	212	41	213
rect	40	213	41	214
rect	40	215	41	216
rect	40	216	41	217
rect	40	218	41	219
rect	40	219	41	220
rect	40	221	41	222
rect	40	222	41	223
rect	40	224	41	225
rect	40	225	41	226
rect	40	227	41	228
rect	40	228	41	229
rect	40	230	41	231
rect	40	231	41	232
rect	40	233	41	234
rect	40	234	41	235
rect	40	236	41	237
rect	40	237	41	238
rect	40	239	41	240
rect	40	240	41	241
rect	40	242	41	243
rect	40	243	41	244
rect	40	245	41	246
rect	40	246	41	247
rect	40	248	41	249
rect	40	249	41	250
rect	40	251	41	252
rect	40	252	41	253
rect	40	254	41	255
rect	40	255	41	256
rect	40	257	41	258
rect	40	258	41	259
rect	40	260	41	261
rect	40	261	41	262
rect	40	263	41	264
rect	40	264	41	265
rect	40	266	41	267
rect	40	267	41	268
rect	40	269	41	270
rect	40	270	41	271
rect	40	272	41	273
rect	40	273	41	274
rect	40	275	41	276
rect	40	276	41	277
rect	40	278	41	279
rect	40	279	41	280
rect	40	281	41	282
rect	40	282	41	283
rect	40	284	41	285
rect	40	285	41	286
rect	40	287	41	288
rect	40	288	41	289
rect	40	290	41	291
rect	41	0	42	1
rect	41	2	42	3
rect	41	3	42	4
rect	41	5	42	6
rect	41	6	42	7
rect	41	8	42	9
rect	41	9	42	10
rect	41	11	42	12
rect	41	12	42	13
rect	41	14	42	15
rect	41	15	42	16
rect	41	17	42	18
rect	41	18	42	19
rect	41	20	42	21
rect	41	21	42	22
rect	41	23	42	24
rect	41	24	42	25
rect	41	26	42	27
rect	41	27	42	28
rect	41	29	42	30
rect	41	30	42	31
rect	41	32	42	33
rect	41	33	42	34
rect	41	35	42	36
rect	41	36	42	37
rect	41	38	42	39
rect	41	39	42	40
rect	41	41	42	42
rect	41	42	42	43
rect	41	44	42	45
rect	41	45	42	46
rect	41	47	42	48
rect	41	48	42	49
rect	41	50	42	51
rect	41	51	42	52
rect	41	53	42	54
rect	41	54	42	55
rect	41	56	42	57
rect	41	57	42	58
rect	41	59	42	60
rect	41	60	42	61
rect	41	62	42	63
rect	41	63	42	64
rect	41	65	42	66
rect	41	66	42	67
rect	41	68	42	69
rect	41	69	42	70
rect	41	71	42	72
rect	41	72	42	73
rect	41	74	42	75
rect	41	75	42	76
rect	41	77	42	78
rect	41	78	42	79
rect	41	80	42	81
rect	41	81	42	82
rect	41	83	42	84
rect	41	84	42	85
rect	41	86	42	87
rect	41	87	42	88
rect	41	89	42	90
rect	41	90	42	91
rect	41	92	42	93
rect	41	93	42	94
rect	41	95	42	96
rect	41	96	42	97
rect	41	98	42	99
rect	41	99	42	100
rect	41	101	42	102
rect	41	102	42	103
rect	41	104	42	105
rect	41	105	42	106
rect	41	107	42	108
rect	41	108	42	109
rect	41	110	42	111
rect	41	111	42	112
rect	41	113	42	114
rect	41	114	42	115
rect	41	116	42	117
rect	41	117	42	118
rect	41	119	42	120
rect	41	120	42	121
rect	41	122	42	123
rect	41	123	42	124
rect	41	125	42	126
rect	41	126	42	127
rect	41	128	42	129
rect	41	129	42	130
rect	41	131	42	132
rect	41	132	42	133
rect	41	134	42	135
rect	41	135	42	136
rect	41	137	42	138
rect	41	138	42	139
rect	41	140	42	141
rect	41	141	42	142
rect	41	143	42	144
rect	41	144	42	145
rect	41	146	42	147
rect	41	147	42	148
rect	41	149	42	150
rect	41	150	42	151
rect	41	152	42	153
rect	41	153	42	154
rect	41	155	42	156
rect	41	156	42	157
rect	41	158	42	159
rect	41	159	42	160
rect	41	161	42	162
rect	41	162	42	163
rect	41	164	42	165
rect	41	165	42	166
rect	41	167	42	168
rect	41	168	42	169
rect	41	170	42	171
rect	41	171	42	172
rect	41	173	42	174
rect	41	174	42	175
rect	41	176	42	177
rect	41	177	42	178
rect	41	179	42	180
rect	41	180	42	181
rect	41	182	42	183
rect	41	183	42	184
rect	41	185	42	186
rect	41	186	42	187
rect	41	188	42	189
rect	41	189	42	190
rect	41	191	42	192
rect	41	192	42	193
rect	41	194	42	195
rect	41	195	42	196
rect	41	197	42	198
rect	41	198	42	199
rect	41	200	42	201
rect	41	201	42	202
rect	41	203	42	204
rect	41	204	42	205
rect	41	206	42	207
rect	41	207	42	208
rect	41	209	42	210
rect	41	210	42	211
rect	41	212	42	213
rect	41	213	42	214
rect	41	215	42	216
rect	41	216	42	217
rect	41	218	42	219
rect	41	219	42	220
rect	41	221	42	222
rect	41	222	42	223
rect	41	224	42	225
rect	41	225	42	226
rect	41	227	42	228
rect	41	228	42	229
rect	41	230	42	231
rect	41	231	42	232
rect	41	233	42	234
rect	41	234	42	235
rect	41	236	42	237
rect	41	237	42	238
rect	41	239	42	240
rect	41	240	42	241
rect	41	242	42	243
rect	41	243	42	244
rect	41	245	42	246
rect	41	246	42	247
rect	41	248	42	249
rect	41	249	42	250
rect	41	251	42	252
rect	41	252	42	253
rect	41	254	42	255
rect	41	255	42	256
rect	41	257	42	258
rect	41	258	42	259
rect	41	260	42	261
rect	41	261	42	262
rect	41	263	42	264
rect	41	264	42	265
rect	41	266	42	267
rect	41	267	42	268
rect	41	269	42	270
rect	41	270	42	271
rect	41	272	42	273
rect	41	273	42	274
rect	41	275	42	276
rect	41	276	42	277
rect	41	278	42	279
rect	41	279	42	280
rect	41	281	42	282
rect	41	282	42	283
rect	41	284	42	285
rect	41	285	42	286
rect	41	287	42	288
rect	41	288	42	289
rect	41	290	42	291
rect	42	0	43	1
rect	42	2	43	3
rect	42	3	43	4
rect	42	5	43	6
rect	42	6	43	7
rect	42	8	43	9
rect	42	9	43	10
rect	42	11	43	12
rect	42	12	43	13
rect	42	14	43	15
rect	42	15	43	16
rect	42	17	43	18
rect	42	18	43	19
rect	42	20	43	21
rect	42	21	43	22
rect	42	23	43	24
rect	42	24	43	25
rect	42	26	43	27
rect	42	27	43	28
rect	42	29	43	30
rect	42	30	43	31
rect	42	32	43	33
rect	42	33	43	34
rect	42	35	43	36
rect	42	36	43	37
rect	42	38	43	39
rect	42	39	43	40
rect	42	41	43	42
rect	42	42	43	43
rect	42	44	43	45
rect	42	45	43	46
rect	42	47	43	48
rect	42	48	43	49
rect	42	50	43	51
rect	42	51	43	52
rect	42	53	43	54
rect	42	54	43	55
rect	42	56	43	57
rect	42	57	43	58
rect	42	59	43	60
rect	42	60	43	61
rect	42	62	43	63
rect	42	63	43	64
rect	42	65	43	66
rect	42	66	43	67
rect	42	68	43	69
rect	42	69	43	70
rect	42	71	43	72
rect	42	72	43	73
rect	42	74	43	75
rect	42	75	43	76
rect	42	77	43	78
rect	42	78	43	79
rect	42	80	43	81
rect	42	81	43	82
rect	42	83	43	84
rect	42	84	43	85
rect	42	86	43	87
rect	42	87	43	88
rect	42	89	43	90
rect	42	90	43	91
rect	42	92	43	93
rect	42	93	43	94
rect	42	95	43	96
rect	42	96	43	97
rect	42	98	43	99
rect	42	99	43	100
rect	42	101	43	102
rect	42	102	43	103
rect	42	104	43	105
rect	42	105	43	106
rect	42	107	43	108
rect	42	108	43	109
rect	42	110	43	111
rect	42	111	43	112
rect	42	113	43	114
rect	42	114	43	115
rect	42	116	43	117
rect	42	117	43	118
rect	42	119	43	120
rect	42	120	43	121
rect	42	122	43	123
rect	42	123	43	124
rect	42	125	43	126
rect	42	126	43	127
rect	42	128	43	129
rect	42	129	43	130
rect	42	131	43	132
rect	42	132	43	133
rect	42	134	43	135
rect	42	135	43	136
rect	42	137	43	138
rect	42	138	43	139
rect	42	140	43	141
rect	42	141	43	142
rect	42	143	43	144
rect	42	144	43	145
rect	42	146	43	147
rect	42	147	43	148
rect	42	149	43	150
rect	42	150	43	151
rect	42	152	43	153
rect	42	153	43	154
rect	42	155	43	156
rect	42	156	43	157
rect	42	158	43	159
rect	42	159	43	160
rect	42	161	43	162
rect	42	162	43	163
rect	42	164	43	165
rect	42	165	43	166
rect	42	167	43	168
rect	42	168	43	169
rect	42	170	43	171
rect	42	171	43	172
rect	42	173	43	174
rect	42	174	43	175
rect	42	176	43	177
rect	42	177	43	178
rect	42	179	43	180
rect	42	180	43	181
rect	42	182	43	183
rect	42	183	43	184
rect	42	185	43	186
rect	42	186	43	187
rect	42	188	43	189
rect	42	189	43	190
rect	42	191	43	192
rect	42	192	43	193
rect	42	194	43	195
rect	42	195	43	196
rect	42	197	43	198
rect	42	198	43	199
rect	42	200	43	201
rect	42	201	43	202
rect	42	203	43	204
rect	42	204	43	205
rect	42	206	43	207
rect	42	207	43	208
rect	42	209	43	210
rect	42	210	43	211
rect	42	212	43	213
rect	42	213	43	214
rect	42	215	43	216
rect	42	216	43	217
rect	42	218	43	219
rect	42	219	43	220
rect	42	221	43	222
rect	42	222	43	223
rect	42	224	43	225
rect	42	225	43	226
rect	42	227	43	228
rect	42	228	43	229
rect	42	230	43	231
rect	42	231	43	232
rect	42	233	43	234
rect	42	234	43	235
rect	42	236	43	237
rect	42	237	43	238
rect	42	239	43	240
rect	42	240	43	241
rect	42	242	43	243
rect	42	243	43	244
rect	42	245	43	246
rect	42	246	43	247
rect	42	248	43	249
rect	42	249	43	250
rect	42	251	43	252
rect	42	252	43	253
rect	42	254	43	255
rect	42	255	43	256
rect	42	257	43	258
rect	42	258	43	259
rect	42	260	43	261
rect	42	261	43	262
rect	42	263	43	264
rect	42	264	43	265
rect	42	266	43	267
rect	42	267	43	268
rect	42	269	43	270
rect	42	270	43	271
rect	42	272	43	273
rect	42	273	43	274
rect	42	275	43	276
rect	42	276	43	277
rect	42	278	43	279
rect	42	279	43	280
rect	42	281	43	282
rect	42	282	43	283
rect	42	284	43	285
rect	42	285	43	286
rect	42	287	43	288
rect	42	288	43	289
rect	42	290	43	291
rect	43	0	44	1
rect	43	2	44	3
rect	43	3	44	4
rect	43	5	44	6
rect	43	6	44	7
rect	43	8	44	9
rect	43	9	44	10
rect	43	11	44	12
rect	43	12	44	13
rect	43	14	44	15
rect	43	15	44	16
rect	43	17	44	18
rect	43	18	44	19
rect	43	20	44	21
rect	43	21	44	22
rect	43	23	44	24
rect	43	24	44	25
rect	43	26	44	27
rect	43	27	44	28
rect	43	29	44	30
rect	43	30	44	31
rect	43	32	44	33
rect	43	33	44	34
rect	43	35	44	36
rect	43	36	44	37
rect	43	38	44	39
rect	43	39	44	40
rect	43	41	44	42
rect	43	42	44	43
rect	43	44	44	45
rect	43	45	44	46
rect	43	47	44	48
rect	43	48	44	49
rect	43	50	44	51
rect	43	51	44	52
rect	43	53	44	54
rect	43	54	44	55
rect	43	56	44	57
rect	43	57	44	58
rect	43	59	44	60
rect	43	60	44	61
rect	43	62	44	63
rect	43	63	44	64
rect	43	65	44	66
rect	43	66	44	67
rect	43	68	44	69
rect	43	69	44	70
rect	43	71	44	72
rect	43	72	44	73
rect	43	74	44	75
rect	43	75	44	76
rect	43	77	44	78
rect	43	78	44	79
rect	43	80	44	81
rect	43	81	44	82
rect	43	83	44	84
rect	43	84	44	85
rect	43	86	44	87
rect	43	87	44	88
rect	43	89	44	90
rect	43	90	44	91
rect	43	92	44	93
rect	43	93	44	94
rect	43	95	44	96
rect	43	96	44	97
rect	43	98	44	99
rect	43	99	44	100
rect	43	101	44	102
rect	43	102	44	103
rect	43	104	44	105
rect	43	105	44	106
rect	43	107	44	108
rect	43	108	44	109
rect	43	110	44	111
rect	43	111	44	112
rect	43	113	44	114
rect	43	114	44	115
rect	43	116	44	117
rect	43	117	44	118
rect	43	119	44	120
rect	43	120	44	121
rect	43	122	44	123
rect	43	123	44	124
rect	43	125	44	126
rect	43	126	44	127
rect	43	128	44	129
rect	43	129	44	130
rect	43	131	44	132
rect	43	132	44	133
rect	43	134	44	135
rect	43	135	44	136
rect	43	137	44	138
rect	43	138	44	139
rect	43	140	44	141
rect	43	141	44	142
rect	43	143	44	144
rect	43	144	44	145
rect	43	146	44	147
rect	43	147	44	148
rect	43	149	44	150
rect	43	150	44	151
rect	43	152	44	153
rect	43	153	44	154
rect	43	155	44	156
rect	43	156	44	157
rect	43	158	44	159
rect	43	159	44	160
rect	43	161	44	162
rect	43	162	44	163
rect	43	164	44	165
rect	43	165	44	166
rect	43	167	44	168
rect	43	168	44	169
rect	43	170	44	171
rect	43	171	44	172
rect	43	173	44	174
rect	43	174	44	175
rect	43	176	44	177
rect	43	177	44	178
rect	43	179	44	180
rect	43	180	44	181
rect	43	182	44	183
rect	43	183	44	184
rect	43	185	44	186
rect	43	186	44	187
rect	43	188	44	189
rect	43	189	44	190
rect	43	191	44	192
rect	43	192	44	193
rect	43	194	44	195
rect	43	195	44	196
rect	43	197	44	198
rect	43	198	44	199
rect	43	200	44	201
rect	43	201	44	202
rect	43	203	44	204
rect	43	204	44	205
rect	43	206	44	207
rect	43	207	44	208
rect	43	209	44	210
rect	43	210	44	211
rect	43	212	44	213
rect	43	213	44	214
rect	43	215	44	216
rect	43	216	44	217
rect	43	218	44	219
rect	43	219	44	220
rect	43	221	44	222
rect	43	222	44	223
rect	43	224	44	225
rect	43	225	44	226
rect	43	227	44	228
rect	43	228	44	229
rect	43	230	44	231
rect	43	231	44	232
rect	43	233	44	234
rect	43	234	44	235
rect	43	236	44	237
rect	43	237	44	238
rect	43	239	44	240
rect	43	240	44	241
rect	43	242	44	243
rect	43	243	44	244
rect	43	245	44	246
rect	43	246	44	247
rect	43	248	44	249
rect	43	249	44	250
rect	43	251	44	252
rect	43	252	44	253
rect	43	254	44	255
rect	43	255	44	256
rect	43	257	44	258
rect	43	258	44	259
rect	43	260	44	261
rect	43	261	44	262
rect	43	263	44	264
rect	43	264	44	265
rect	43	266	44	267
rect	43	267	44	268
rect	43	269	44	270
rect	43	270	44	271
rect	43	272	44	273
rect	43	273	44	274
rect	43	275	44	276
rect	43	276	44	277
rect	43	278	44	279
rect	43	279	44	280
rect	43	281	44	282
rect	43	282	44	283
rect	43	284	44	285
rect	43	285	44	286
rect	43	287	44	288
rect	43	288	44	289
rect	43	290	44	291
rect	48	0	49	1
rect	48	2	49	3
rect	48	3	49	4
rect	48	5	49	6
rect	48	6	49	7
rect	48	8	49	9
rect	48	9	49	10
rect	48	11	49	12
rect	48	12	49	13
rect	48	14	49	15
rect	48	15	49	16
rect	48	17	49	18
rect	48	18	49	19
rect	48	20	49	21
rect	48	21	49	22
rect	48	23	49	24
rect	48	24	49	25
rect	48	26	49	27
rect	48	27	49	28
rect	48	29	49	30
rect	48	30	49	31
rect	48	32	49	33
rect	48	33	49	34
rect	48	35	49	36
rect	48	36	49	37
rect	48	38	49	39
rect	48	39	49	40
rect	48	41	49	42
rect	48	42	49	43
rect	48	44	49	45
rect	48	45	49	46
rect	48	47	49	48
rect	48	48	49	49
rect	48	50	49	51
rect	48	51	49	52
rect	48	53	49	54
rect	48	54	49	55
rect	48	56	49	57
rect	48	57	49	58
rect	48	59	49	60
rect	48	60	49	61
rect	48	62	49	63
rect	48	63	49	64
rect	48	65	49	66
rect	48	66	49	67
rect	48	68	49	69
rect	48	69	49	70
rect	48	71	49	72
rect	48	72	49	73
rect	48	74	49	75
rect	48	75	49	76
rect	48	77	49	78
rect	48	78	49	79
rect	48	80	49	81
rect	48	81	49	82
rect	48	83	49	84
rect	48	84	49	85
rect	48	86	49	87
rect	48	87	49	88
rect	48	89	49	90
rect	48	90	49	91
rect	48	92	49	93
rect	48	93	49	94
rect	48	95	49	96
rect	48	96	49	97
rect	48	98	49	99
rect	48	99	49	100
rect	48	101	49	102
rect	48	102	49	103
rect	48	104	49	105
rect	48	105	49	106
rect	48	107	49	108
rect	48	108	49	109
rect	48	110	49	111
rect	48	111	49	112
rect	48	113	49	114
rect	48	114	49	115
rect	48	116	49	117
rect	48	117	49	118
rect	48	119	49	120
rect	48	120	49	121
rect	48	122	49	123
rect	48	123	49	124
rect	48	125	49	126
rect	48	126	49	127
rect	48	128	49	129
rect	48	129	49	130
rect	48	131	49	132
rect	48	132	49	133
rect	48	134	49	135
rect	48	135	49	136
rect	48	137	49	138
rect	48	138	49	139
rect	48	140	49	141
rect	48	141	49	142
rect	48	143	49	144
rect	48	144	49	145
rect	48	146	49	147
rect	48	147	49	148
rect	48	149	49	150
rect	48	150	49	151
rect	48	152	49	153
rect	48	153	49	154
rect	48	155	49	156
rect	48	156	49	157
rect	48	158	49	159
rect	48	159	49	160
rect	48	161	49	162
rect	48	162	49	163
rect	48	164	49	165
rect	48	165	49	166
rect	48	167	49	168
rect	48	168	49	169
rect	48	170	49	171
rect	48	171	49	172
rect	48	173	49	174
rect	48	174	49	175
rect	48	176	49	177
rect	48	177	49	178
rect	48	179	49	180
rect	48	180	49	181
rect	48	182	49	183
rect	48	183	49	184
rect	48	185	49	186
rect	48	186	49	187
rect	48	188	49	189
rect	48	189	49	190
rect	48	191	49	192
rect	48	192	49	193
rect	48	194	49	195
rect	48	195	49	196
rect	48	197	49	198
rect	48	198	49	199
rect	48	200	49	201
rect	48	201	49	202
rect	48	203	49	204
rect	48	204	49	205
rect	48	206	49	207
rect	48	207	49	208
rect	48	209	49	210
rect	48	210	49	211
rect	48	212	49	213
rect	48	213	49	214
rect	48	215	49	216
rect	48	216	49	217
rect	48	218	49	219
rect	48	219	49	220
rect	48	221	49	222
rect	48	222	49	223
rect	48	224	49	225
rect	48	225	49	226
rect	48	227	49	228
rect	48	228	49	229
rect	48	230	49	231
rect	48	231	49	232
rect	48	233	49	234
rect	48	234	49	235
rect	48	236	49	237
rect	48	237	49	238
rect	48	239	49	240
rect	48	240	49	241
rect	48	242	49	243
rect	48	243	49	244
rect	48	245	49	246
rect	48	246	49	247
rect	48	248	49	249
rect	48	249	49	250
rect	48	251	49	252
rect	48	252	49	253
rect	48	254	49	255
rect	48	255	49	256
rect	48	257	49	258
rect	48	258	49	259
rect	48	260	49	261
rect	48	261	49	262
rect	48	263	49	264
rect	48	264	49	265
rect	48	266	49	267
rect	48	267	49	268
rect	48	269	49	270
rect	48	270	49	271
rect	48	272	49	273
rect	48	273	49	274
rect	48	275	49	276
rect	48	276	49	277
rect	48	278	49	279
rect	48	279	49	280
rect	48	281	49	282
rect	48	282	49	283
rect	48	284	49	285
rect	48	285	49	286
rect	48	287	49	288
rect	48	288	49	289
rect	48	290	49	291
rect	50	0	51	1
rect	50	2	51	3
rect	50	3	51	4
rect	50	5	51	6
rect	50	6	51	7
rect	50	8	51	9
rect	50	9	51	10
rect	50	11	51	12
rect	50	12	51	13
rect	50	14	51	15
rect	50	15	51	16
rect	50	17	51	18
rect	50	18	51	19
rect	50	20	51	21
rect	50	21	51	22
rect	50	23	51	24
rect	50	24	51	25
rect	50	26	51	27
rect	50	27	51	28
rect	50	29	51	30
rect	50	30	51	31
rect	50	32	51	33
rect	50	33	51	34
rect	50	35	51	36
rect	50	36	51	37
rect	50	38	51	39
rect	50	39	51	40
rect	50	41	51	42
rect	50	42	51	43
rect	50	44	51	45
rect	50	45	51	46
rect	50	47	51	48
rect	50	48	51	49
rect	50	50	51	51
rect	50	51	51	52
rect	50	53	51	54
rect	50	54	51	55
rect	50	56	51	57
rect	50	57	51	58
rect	50	59	51	60
rect	50	60	51	61
rect	50	62	51	63
rect	50	63	51	64
rect	50	65	51	66
rect	50	66	51	67
rect	50	68	51	69
rect	50	69	51	70
rect	50	71	51	72
rect	50	72	51	73
rect	50	74	51	75
rect	50	75	51	76
rect	50	77	51	78
rect	50	78	51	79
rect	50	80	51	81
rect	50	81	51	82
rect	50	83	51	84
rect	50	84	51	85
rect	50	86	51	87
rect	50	87	51	88
rect	50	89	51	90
rect	50	90	51	91
rect	50	92	51	93
rect	50	93	51	94
rect	50	95	51	96
rect	50	96	51	97
rect	50	98	51	99
rect	50	99	51	100
rect	50	101	51	102
rect	50	102	51	103
rect	50	104	51	105
rect	50	105	51	106
rect	50	107	51	108
rect	50	108	51	109
rect	50	110	51	111
rect	50	111	51	112
rect	50	113	51	114
rect	50	114	51	115
rect	50	116	51	117
rect	50	117	51	118
rect	50	119	51	120
rect	50	120	51	121
rect	50	122	51	123
rect	50	123	51	124
rect	50	125	51	126
rect	50	126	51	127
rect	50	128	51	129
rect	50	129	51	130
rect	50	131	51	132
rect	50	132	51	133
rect	50	134	51	135
rect	50	135	51	136
rect	50	137	51	138
rect	50	138	51	139
rect	50	140	51	141
rect	50	141	51	142
rect	50	143	51	144
rect	50	144	51	145
rect	50	146	51	147
rect	50	147	51	148
rect	50	149	51	150
rect	50	150	51	151
rect	50	152	51	153
rect	50	153	51	154
rect	50	155	51	156
rect	50	156	51	157
rect	50	158	51	159
rect	50	159	51	160
rect	50	161	51	162
rect	50	162	51	163
rect	50	164	51	165
rect	50	165	51	166
rect	50	167	51	168
rect	50	168	51	169
rect	50	170	51	171
rect	50	171	51	172
rect	50	173	51	174
rect	50	174	51	175
rect	50	176	51	177
rect	50	177	51	178
rect	50	179	51	180
rect	50	180	51	181
rect	50	182	51	183
rect	50	183	51	184
rect	50	185	51	186
rect	50	186	51	187
rect	50	188	51	189
rect	50	189	51	190
rect	50	191	51	192
rect	50	192	51	193
rect	50	194	51	195
rect	50	195	51	196
rect	50	197	51	198
rect	50	198	51	199
rect	50	200	51	201
rect	50	201	51	202
rect	50	203	51	204
rect	50	204	51	205
rect	50	206	51	207
rect	50	207	51	208
rect	50	209	51	210
rect	50	210	51	211
rect	50	212	51	213
rect	50	213	51	214
rect	50	215	51	216
rect	50	216	51	217
rect	50	218	51	219
rect	50	219	51	220
rect	50	221	51	222
rect	50	222	51	223
rect	50	224	51	225
rect	50	225	51	226
rect	50	227	51	228
rect	50	228	51	229
rect	50	230	51	231
rect	50	231	51	232
rect	50	233	51	234
rect	50	234	51	235
rect	50	236	51	237
rect	50	237	51	238
rect	50	239	51	240
rect	50	240	51	241
rect	50	242	51	243
rect	50	243	51	244
rect	50	245	51	246
rect	50	246	51	247
rect	50	248	51	249
rect	50	249	51	250
rect	50	251	51	252
rect	50	252	51	253
rect	50	254	51	255
rect	50	255	51	256
rect	50	257	51	258
rect	50	258	51	259
rect	50	260	51	261
rect	50	261	51	262
rect	50	263	51	264
rect	50	264	51	265
rect	50	266	51	267
rect	50	267	51	268
rect	50	269	51	270
rect	50	270	51	271
rect	50	272	51	273
rect	50	273	51	274
rect	50	275	51	276
rect	50	276	51	277
rect	50	278	51	279
rect	50	279	51	280
rect	50	281	51	282
rect	50	282	51	283
rect	50	284	51	285
rect	50	285	51	286
rect	50	287	51	288
rect	50	288	51	289
rect	50	290	51	291
rect	50	291	51	292
rect	50	293	51	294
rect	50	294	51	295
rect	50	296	51	297
rect	50	297	51	298
rect	50	299	51	300
rect	50	300	51	301
rect	50	302	51	303
rect	50	303	51	304
rect	50	305	51	306
rect	50	306	51	307
rect	50	308	51	309
rect	50	309	51	310
rect	50	311	51	312
rect	51	0	52	1
rect	51	2	52	3
rect	51	3	52	4
rect	51	5	52	6
rect	51	6	52	7
rect	51	8	52	9
rect	51	9	52	10
rect	51	11	52	12
rect	51	12	52	13
rect	51	14	52	15
rect	51	15	52	16
rect	51	17	52	18
rect	51	18	52	19
rect	51	20	52	21
rect	51	21	52	22
rect	51	23	52	24
rect	51	24	52	25
rect	51	26	52	27
rect	51	27	52	28
rect	51	29	52	30
rect	51	30	52	31
rect	51	32	52	33
rect	51	33	52	34
rect	51	35	52	36
rect	51	36	52	37
rect	51	38	52	39
rect	51	39	52	40
rect	51	41	52	42
rect	51	42	52	43
rect	51	44	52	45
rect	51	45	52	46
rect	51	47	52	48
rect	51	48	52	49
rect	51	50	52	51
rect	51	51	52	52
rect	51	53	52	54
rect	51	54	52	55
rect	51	56	52	57
rect	51	57	52	58
rect	51	59	52	60
rect	51	60	52	61
rect	51	62	52	63
rect	51	63	52	64
rect	51	65	52	66
rect	51	66	52	67
rect	51	68	52	69
rect	51	69	52	70
rect	51	71	52	72
rect	51	72	52	73
rect	51	74	52	75
rect	51	75	52	76
rect	51	77	52	78
rect	51	78	52	79
rect	51	80	52	81
rect	51	81	52	82
rect	51	83	52	84
rect	51	84	52	85
rect	51	86	52	87
rect	51	87	52	88
rect	51	89	52	90
rect	51	90	52	91
rect	51	92	52	93
rect	51	93	52	94
rect	51	95	52	96
rect	51	96	52	97
rect	51	98	52	99
rect	51	99	52	100
rect	51	101	52	102
rect	51	102	52	103
rect	51	104	52	105
rect	51	105	52	106
rect	51	107	52	108
rect	51	108	52	109
rect	51	110	52	111
rect	51	111	52	112
rect	51	113	52	114
rect	51	114	52	115
rect	51	116	52	117
rect	51	117	52	118
rect	51	119	52	120
rect	51	120	52	121
rect	51	122	52	123
rect	51	123	52	124
rect	51	125	52	126
rect	51	126	52	127
rect	51	128	52	129
rect	51	129	52	130
rect	51	131	52	132
rect	51	132	52	133
rect	51	134	52	135
rect	51	135	52	136
rect	51	137	52	138
rect	51	138	52	139
rect	51	140	52	141
rect	51	141	52	142
rect	51	143	52	144
rect	51	144	52	145
rect	51	146	52	147
rect	51	147	52	148
rect	51	149	52	150
rect	51	150	52	151
rect	51	152	52	153
rect	51	153	52	154
rect	51	155	52	156
rect	51	156	52	157
rect	51	158	52	159
rect	51	159	52	160
rect	51	161	52	162
rect	51	162	52	163
rect	51	164	52	165
rect	51	165	52	166
rect	51	167	52	168
rect	51	168	52	169
rect	51	170	52	171
rect	51	171	52	172
rect	51	173	52	174
rect	51	174	52	175
rect	51	176	52	177
rect	51	177	52	178
rect	51	179	52	180
rect	51	180	52	181
rect	51	182	52	183
rect	51	183	52	184
rect	51	185	52	186
rect	51	186	52	187
rect	51	188	52	189
rect	51	189	52	190
rect	51	191	52	192
rect	51	192	52	193
rect	51	194	52	195
rect	51	195	52	196
rect	51	197	52	198
rect	51	198	52	199
rect	51	200	52	201
rect	51	201	52	202
rect	51	203	52	204
rect	51	204	52	205
rect	51	206	52	207
rect	51	207	52	208
rect	51	209	52	210
rect	51	210	52	211
rect	51	212	52	213
rect	51	213	52	214
rect	51	215	52	216
rect	51	216	52	217
rect	51	218	52	219
rect	51	219	52	220
rect	51	221	52	222
rect	51	222	52	223
rect	51	224	52	225
rect	51	225	52	226
rect	51	227	52	228
rect	51	228	52	229
rect	51	230	52	231
rect	51	231	52	232
rect	51	233	52	234
rect	51	234	52	235
rect	51	236	52	237
rect	51	237	52	238
rect	51	239	52	240
rect	51	240	52	241
rect	51	242	52	243
rect	51	243	52	244
rect	51	245	52	246
rect	51	246	52	247
rect	51	248	52	249
rect	51	249	52	250
rect	51	251	52	252
rect	51	252	52	253
rect	51	254	52	255
rect	51	255	52	256
rect	51	257	52	258
rect	51	258	52	259
rect	51	260	52	261
rect	51	261	52	262
rect	51	263	52	264
rect	51	264	52	265
rect	51	266	52	267
rect	51	267	52	268
rect	51	269	52	270
rect	51	270	52	271
rect	51	272	52	273
rect	51	273	52	274
rect	51	275	52	276
rect	51	276	52	277
rect	51	278	52	279
rect	51	279	52	280
rect	51	281	52	282
rect	51	282	52	283
rect	51	284	52	285
rect	51	285	52	286
rect	51	287	52	288
rect	51	288	52	289
rect	51	290	52	291
rect	51	291	52	292
rect	51	293	52	294
rect	51	294	52	295
rect	51	296	52	297
rect	51	297	52	298
rect	51	299	52	300
rect	51	300	52	301
rect	51	302	52	303
rect	51	303	52	304
rect	51	305	52	306
rect	51	306	52	307
rect	51	308	52	309
rect	51	309	52	310
rect	51	311	52	312
rect	52	0	53	1
rect	52	2	53	3
rect	52	3	53	4
rect	52	5	53	6
rect	52	6	53	7
rect	52	8	53	9
rect	52	9	53	10
rect	52	11	53	12
rect	52	12	53	13
rect	52	14	53	15
rect	52	15	53	16
rect	52	17	53	18
rect	52	18	53	19
rect	52	20	53	21
rect	52	21	53	22
rect	52	23	53	24
rect	52	24	53	25
rect	52	26	53	27
rect	52	27	53	28
rect	52	29	53	30
rect	52	30	53	31
rect	52	32	53	33
rect	52	33	53	34
rect	52	35	53	36
rect	52	36	53	37
rect	52	38	53	39
rect	52	39	53	40
rect	52	41	53	42
rect	52	42	53	43
rect	52	44	53	45
rect	52	45	53	46
rect	52	47	53	48
rect	52	48	53	49
rect	52	50	53	51
rect	52	51	53	52
rect	52	53	53	54
rect	52	54	53	55
rect	52	56	53	57
rect	52	57	53	58
rect	52	59	53	60
rect	52	60	53	61
rect	52	62	53	63
rect	52	63	53	64
rect	52	65	53	66
rect	52	66	53	67
rect	52	68	53	69
rect	52	69	53	70
rect	52	71	53	72
rect	52	72	53	73
rect	52	74	53	75
rect	52	75	53	76
rect	52	77	53	78
rect	52	78	53	79
rect	52	80	53	81
rect	52	81	53	82
rect	52	83	53	84
rect	52	84	53	85
rect	52	86	53	87
rect	52	87	53	88
rect	52	89	53	90
rect	52	90	53	91
rect	52	92	53	93
rect	52	93	53	94
rect	52	95	53	96
rect	52	96	53	97
rect	52	98	53	99
rect	52	99	53	100
rect	52	101	53	102
rect	52	102	53	103
rect	52	104	53	105
rect	52	105	53	106
rect	52	107	53	108
rect	52	108	53	109
rect	52	110	53	111
rect	52	111	53	112
rect	52	113	53	114
rect	52	114	53	115
rect	52	116	53	117
rect	52	117	53	118
rect	52	119	53	120
rect	52	120	53	121
rect	52	122	53	123
rect	52	123	53	124
rect	52	125	53	126
rect	52	126	53	127
rect	52	128	53	129
rect	52	129	53	130
rect	52	131	53	132
rect	52	132	53	133
rect	52	134	53	135
rect	52	135	53	136
rect	52	137	53	138
rect	52	138	53	139
rect	52	140	53	141
rect	52	141	53	142
rect	52	143	53	144
rect	52	144	53	145
rect	52	146	53	147
rect	52	147	53	148
rect	52	149	53	150
rect	52	150	53	151
rect	52	152	53	153
rect	52	153	53	154
rect	52	155	53	156
rect	52	156	53	157
rect	52	158	53	159
rect	52	159	53	160
rect	52	161	53	162
rect	52	162	53	163
rect	52	164	53	165
rect	52	165	53	166
rect	52	167	53	168
rect	52	168	53	169
rect	52	170	53	171
rect	52	171	53	172
rect	52	173	53	174
rect	52	174	53	175
rect	52	176	53	177
rect	52	177	53	178
rect	52	179	53	180
rect	52	180	53	181
rect	52	182	53	183
rect	52	183	53	184
rect	52	185	53	186
rect	52	186	53	187
rect	52	188	53	189
rect	52	189	53	190
rect	52	191	53	192
rect	52	192	53	193
rect	52	194	53	195
rect	52	195	53	196
rect	52	197	53	198
rect	52	198	53	199
rect	52	200	53	201
rect	52	201	53	202
rect	52	203	53	204
rect	52	204	53	205
rect	52	206	53	207
rect	52	207	53	208
rect	52	209	53	210
rect	52	210	53	211
rect	52	212	53	213
rect	52	213	53	214
rect	52	215	53	216
rect	52	216	53	217
rect	52	218	53	219
rect	52	219	53	220
rect	52	221	53	222
rect	52	222	53	223
rect	52	224	53	225
rect	52	225	53	226
rect	52	227	53	228
rect	52	228	53	229
rect	52	230	53	231
rect	52	231	53	232
rect	52	233	53	234
rect	52	234	53	235
rect	52	236	53	237
rect	52	237	53	238
rect	52	239	53	240
rect	52	240	53	241
rect	52	242	53	243
rect	52	243	53	244
rect	52	245	53	246
rect	52	246	53	247
rect	52	248	53	249
rect	52	249	53	250
rect	52	251	53	252
rect	52	252	53	253
rect	52	254	53	255
rect	52	255	53	256
rect	52	257	53	258
rect	52	258	53	259
rect	52	260	53	261
rect	52	261	53	262
rect	52	263	53	264
rect	52	264	53	265
rect	52	266	53	267
rect	52	267	53	268
rect	52	269	53	270
rect	52	270	53	271
rect	52	272	53	273
rect	52	273	53	274
rect	52	275	53	276
rect	52	276	53	277
rect	52	278	53	279
rect	52	279	53	280
rect	52	281	53	282
rect	52	282	53	283
rect	52	284	53	285
rect	52	285	53	286
rect	52	287	53	288
rect	52	288	53	289
rect	52	290	53	291
rect	52	291	53	292
rect	52	293	53	294
rect	52	294	53	295
rect	52	296	53	297
rect	52	297	53	298
rect	52	299	53	300
rect	52	300	53	301
rect	52	302	53	303
rect	52	303	53	304
rect	52	305	53	306
rect	52	306	53	307
rect	52	308	53	309
rect	52	309	53	310
rect	52	311	53	312
rect	53	0	54	1
rect	53	2	54	3
rect	53	3	54	4
rect	53	5	54	6
rect	53	6	54	7
rect	53	8	54	9
rect	53	9	54	10
rect	53	11	54	12
rect	53	12	54	13
rect	53	14	54	15
rect	53	15	54	16
rect	53	17	54	18
rect	53	18	54	19
rect	53	20	54	21
rect	53	21	54	22
rect	53	23	54	24
rect	53	24	54	25
rect	53	26	54	27
rect	53	27	54	28
rect	53	29	54	30
rect	53	30	54	31
rect	53	32	54	33
rect	53	33	54	34
rect	53	35	54	36
rect	53	36	54	37
rect	53	38	54	39
rect	53	39	54	40
rect	53	41	54	42
rect	53	42	54	43
rect	53	44	54	45
rect	53	45	54	46
rect	53	47	54	48
rect	53	48	54	49
rect	53	50	54	51
rect	53	51	54	52
rect	53	53	54	54
rect	53	54	54	55
rect	53	56	54	57
rect	53	57	54	58
rect	53	59	54	60
rect	53	60	54	61
rect	53	62	54	63
rect	53	63	54	64
rect	53	65	54	66
rect	53	66	54	67
rect	53	68	54	69
rect	53	69	54	70
rect	53	71	54	72
rect	53	72	54	73
rect	53	74	54	75
rect	53	75	54	76
rect	53	77	54	78
rect	53	78	54	79
rect	53	80	54	81
rect	53	81	54	82
rect	53	83	54	84
rect	53	84	54	85
rect	53	86	54	87
rect	53	87	54	88
rect	53	89	54	90
rect	53	90	54	91
rect	53	92	54	93
rect	53	93	54	94
rect	53	95	54	96
rect	53	96	54	97
rect	53	98	54	99
rect	53	99	54	100
rect	53	101	54	102
rect	53	102	54	103
rect	53	104	54	105
rect	53	105	54	106
rect	53	107	54	108
rect	53	108	54	109
rect	53	110	54	111
rect	53	111	54	112
rect	53	113	54	114
rect	53	114	54	115
rect	53	116	54	117
rect	53	117	54	118
rect	53	119	54	120
rect	53	120	54	121
rect	53	122	54	123
rect	53	123	54	124
rect	53	125	54	126
rect	53	126	54	127
rect	53	128	54	129
rect	53	129	54	130
rect	53	131	54	132
rect	53	132	54	133
rect	53	134	54	135
rect	53	135	54	136
rect	53	137	54	138
rect	53	138	54	139
rect	53	140	54	141
rect	53	141	54	142
rect	53	143	54	144
rect	53	144	54	145
rect	53	146	54	147
rect	53	147	54	148
rect	53	149	54	150
rect	53	150	54	151
rect	53	152	54	153
rect	53	153	54	154
rect	53	155	54	156
rect	53	156	54	157
rect	53	158	54	159
rect	53	159	54	160
rect	53	161	54	162
rect	53	162	54	163
rect	53	164	54	165
rect	53	165	54	166
rect	53	167	54	168
rect	53	168	54	169
rect	53	170	54	171
rect	53	171	54	172
rect	53	173	54	174
rect	53	174	54	175
rect	53	176	54	177
rect	53	177	54	178
rect	53	179	54	180
rect	53	180	54	181
rect	53	182	54	183
rect	53	183	54	184
rect	53	185	54	186
rect	53	186	54	187
rect	53	188	54	189
rect	53	189	54	190
rect	53	191	54	192
rect	53	192	54	193
rect	53	194	54	195
rect	53	195	54	196
rect	53	197	54	198
rect	53	198	54	199
rect	53	200	54	201
rect	53	201	54	202
rect	53	203	54	204
rect	53	204	54	205
rect	53	206	54	207
rect	53	207	54	208
rect	53	209	54	210
rect	53	210	54	211
rect	53	212	54	213
rect	53	213	54	214
rect	53	215	54	216
rect	53	216	54	217
rect	53	218	54	219
rect	53	219	54	220
rect	53	221	54	222
rect	53	222	54	223
rect	53	224	54	225
rect	53	225	54	226
rect	53	227	54	228
rect	53	228	54	229
rect	53	230	54	231
rect	53	231	54	232
rect	53	233	54	234
rect	53	234	54	235
rect	53	236	54	237
rect	53	237	54	238
rect	53	239	54	240
rect	53	240	54	241
rect	53	242	54	243
rect	53	243	54	244
rect	53	245	54	246
rect	53	246	54	247
rect	53	248	54	249
rect	53	249	54	250
rect	53	251	54	252
rect	53	252	54	253
rect	53	254	54	255
rect	53	255	54	256
rect	53	257	54	258
rect	53	258	54	259
rect	53	260	54	261
rect	53	261	54	262
rect	53	263	54	264
rect	53	264	54	265
rect	53	266	54	267
rect	53	267	54	268
rect	53	269	54	270
rect	53	270	54	271
rect	53	272	54	273
rect	53	273	54	274
rect	53	275	54	276
rect	53	276	54	277
rect	53	278	54	279
rect	53	279	54	280
rect	53	281	54	282
rect	53	282	54	283
rect	53	284	54	285
rect	53	285	54	286
rect	53	287	54	288
rect	53	288	54	289
rect	53	290	54	291
rect	53	291	54	292
rect	53	293	54	294
rect	53	294	54	295
rect	53	296	54	297
rect	53	297	54	298
rect	53	299	54	300
rect	53	300	54	301
rect	53	302	54	303
rect	53	303	54	304
rect	53	305	54	306
rect	53	306	54	307
rect	53	308	54	309
rect	53	309	54	310
rect	53	311	54	312
rect	54	0	55	1
rect	54	2	55	3
rect	54	3	55	4
rect	54	5	55	6
rect	54	6	55	7
rect	54	8	55	9
rect	54	9	55	10
rect	54	11	55	12
rect	54	12	55	13
rect	54	14	55	15
rect	54	15	55	16
rect	54	17	55	18
rect	54	18	55	19
rect	54	20	55	21
rect	54	21	55	22
rect	54	23	55	24
rect	54	24	55	25
rect	54	26	55	27
rect	54	27	55	28
rect	54	29	55	30
rect	54	30	55	31
rect	54	32	55	33
rect	54	33	55	34
rect	54	35	55	36
rect	54	36	55	37
rect	54	38	55	39
rect	54	39	55	40
rect	54	41	55	42
rect	54	42	55	43
rect	54	44	55	45
rect	54	45	55	46
rect	54	47	55	48
rect	54	48	55	49
rect	54	50	55	51
rect	54	51	55	52
rect	54	53	55	54
rect	54	54	55	55
rect	54	56	55	57
rect	54	57	55	58
rect	54	59	55	60
rect	54	60	55	61
rect	54	62	55	63
rect	54	63	55	64
rect	54	65	55	66
rect	54	66	55	67
rect	54	68	55	69
rect	54	69	55	70
rect	54	71	55	72
rect	54	72	55	73
rect	54	74	55	75
rect	54	75	55	76
rect	54	77	55	78
rect	54	78	55	79
rect	54	80	55	81
rect	54	81	55	82
rect	54	83	55	84
rect	54	84	55	85
rect	54	86	55	87
rect	54	87	55	88
rect	54	89	55	90
rect	54	90	55	91
rect	54	92	55	93
rect	54	93	55	94
rect	54	95	55	96
rect	54	96	55	97
rect	54	98	55	99
rect	54	99	55	100
rect	54	101	55	102
rect	54	102	55	103
rect	54	104	55	105
rect	54	105	55	106
rect	54	107	55	108
rect	54	108	55	109
rect	54	110	55	111
rect	54	111	55	112
rect	54	113	55	114
rect	54	114	55	115
rect	54	116	55	117
rect	54	117	55	118
rect	54	119	55	120
rect	54	120	55	121
rect	54	122	55	123
rect	54	123	55	124
rect	54	125	55	126
rect	54	126	55	127
rect	54	128	55	129
rect	54	129	55	130
rect	54	131	55	132
rect	54	132	55	133
rect	54	134	55	135
rect	54	135	55	136
rect	54	137	55	138
rect	54	138	55	139
rect	54	140	55	141
rect	54	141	55	142
rect	54	143	55	144
rect	54	144	55	145
rect	54	146	55	147
rect	54	147	55	148
rect	54	149	55	150
rect	54	150	55	151
rect	54	152	55	153
rect	54	153	55	154
rect	54	155	55	156
rect	54	156	55	157
rect	54	158	55	159
rect	54	159	55	160
rect	54	161	55	162
rect	54	162	55	163
rect	54	164	55	165
rect	54	165	55	166
rect	54	167	55	168
rect	54	168	55	169
rect	54	170	55	171
rect	54	171	55	172
rect	54	173	55	174
rect	54	174	55	175
rect	54	176	55	177
rect	54	177	55	178
rect	54	179	55	180
rect	54	180	55	181
rect	54	182	55	183
rect	54	183	55	184
rect	54	185	55	186
rect	54	186	55	187
rect	54	188	55	189
rect	54	189	55	190
rect	54	191	55	192
rect	54	192	55	193
rect	54	194	55	195
rect	54	195	55	196
rect	54	197	55	198
rect	54	198	55	199
rect	54	200	55	201
rect	54	201	55	202
rect	54	203	55	204
rect	54	204	55	205
rect	54	206	55	207
rect	54	207	55	208
rect	54	209	55	210
rect	54	210	55	211
rect	54	212	55	213
rect	54	213	55	214
rect	54	215	55	216
rect	54	216	55	217
rect	54	218	55	219
rect	54	219	55	220
rect	54	221	55	222
rect	54	222	55	223
rect	54	224	55	225
rect	54	225	55	226
rect	54	227	55	228
rect	54	228	55	229
rect	54	230	55	231
rect	54	231	55	232
rect	54	233	55	234
rect	54	234	55	235
rect	54	236	55	237
rect	54	237	55	238
rect	54	239	55	240
rect	54	240	55	241
rect	54	242	55	243
rect	54	243	55	244
rect	54	245	55	246
rect	54	246	55	247
rect	54	248	55	249
rect	54	249	55	250
rect	54	251	55	252
rect	54	252	55	253
rect	54	254	55	255
rect	54	255	55	256
rect	54	257	55	258
rect	54	258	55	259
rect	54	260	55	261
rect	54	261	55	262
rect	54	263	55	264
rect	54	264	55	265
rect	54	266	55	267
rect	54	267	55	268
rect	54	269	55	270
rect	54	270	55	271
rect	54	272	55	273
rect	54	273	55	274
rect	54	275	55	276
rect	54	276	55	277
rect	54	278	55	279
rect	54	279	55	280
rect	54	281	55	282
rect	54	282	55	283
rect	54	284	55	285
rect	54	285	55	286
rect	54	287	55	288
rect	54	288	55	289
rect	54	290	55	291
rect	54	291	55	292
rect	54	293	55	294
rect	54	294	55	295
rect	54	296	55	297
rect	54	297	55	298
rect	54	299	55	300
rect	54	300	55	301
rect	54	302	55	303
rect	54	303	55	304
rect	54	305	55	306
rect	54	306	55	307
rect	54	308	55	309
rect	54	309	55	310
rect	54	311	55	312
rect	65	0	66	1
rect	65	2	66	3
rect	65	3	66	4
rect	65	5	66	6
rect	65	6	66	7
rect	65	8	66	9
rect	65	9	66	10
rect	65	11	66	12
rect	65	12	66	13
rect	65	14	66	15
rect	65	15	66	16
rect	65	17	66	18
rect	65	18	66	19
rect	65	20	66	21
rect	65	21	66	22
rect	65	23	66	24
rect	65	24	66	25
rect	65	26	66	27
rect	65	27	66	28
rect	65	29	66	30
rect	65	30	66	31
rect	65	32	66	33
rect	65	33	66	34
rect	65	35	66	36
rect	65	36	66	37
rect	65	38	66	39
rect	65	39	66	40
rect	65	41	66	42
rect	65	42	66	43
rect	65	44	66	45
rect	65	45	66	46
rect	65	47	66	48
rect	65	48	66	49
rect	65	50	66	51
rect	65	51	66	52
rect	65	53	66	54
rect	65	54	66	55
rect	65	56	66	57
rect	65	57	66	58
rect	65	59	66	60
rect	65	60	66	61
rect	65	62	66	63
rect	65	63	66	64
rect	65	65	66	66
rect	65	66	66	67
rect	65	68	66	69
rect	65	69	66	70
rect	65	71	66	72
rect	65	72	66	73
rect	65	74	66	75
rect	65	75	66	76
rect	65	77	66	78
rect	65	78	66	79
rect	65	80	66	81
rect	65	81	66	82
rect	65	83	66	84
rect	65	84	66	85
rect	65	86	66	87
rect	65	87	66	88
rect	65	89	66	90
rect	65	90	66	91
rect	65	92	66	93
rect	65	93	66	94
rect	65	95	66	96
rect	65	96	66	97
rect	65	98	66	99
rect	65	99	66	100
rect	65	101	66	102
rect	65	102	66	103
rect	65	104	66	105
rect	65	105	66	106
rect	65	107	66	108
rect	65	108	66	109
rect	65	110	66	111
rect	65	111	66	112
rect	65	113	66	114
rect	65	114	66	115
rect	65	116	66	117
rect	65	117	66	118
rect	65	119	66	120
rect	65	120	66	121
rect	65	122	66	123
rect	65	123	66	124
rect	65	125	66	126
rect	65	126	66	127
rect	65	128	66	129
rect	65	129	66	130
rect	65	131	66	132
rect	65	132	66	133
rect	65	134	66	135
rect	65	135	66	136
rect	65	137	66	138
rect	65	138	66	139
rect	65	140	66	141
rect	65	141	66	142
rect	65	143	66	144
rect	65	144	66	145
rect	65	146	66	147
rect	65	147	66	148
rect	65	149	66	150
rect	65	150	66	151
rect	65	152	66	153
rect	65	153	66	154
rect	65	155	66	156
rect	65	156	66	157
rect	65	158	66	159
rect	65	159	66	160
rect	65	161	66	162
rect	65	162	66	163
rect	65	164	66	165
rect	65	165	66	166
rect	65	167	66	168
rect	65	168	66	169
rect	65	170	66	171
rect	65	171	66	172
rect	65	173	66	174
rect	65	174	66	175
rect	65	176	66	177
rect	65	177	66	178
rect	65	179	66	180
rect	65	180	66	181
rect	65	182	66	183
rect	65	183	66	184
rect	65	185	66	186
rect	65	186	66	187
rect	65	188	66	189
rect	65	189	66	190
rect	65	191	66	192
rect	65	192	66	193
rect	65	194	66	195
rect	65	195	66	196
rect	65	197	66	198
rect	65	198	66	199
rect	65	200	66	201
rect	65	201	66	202
rect	65	203	66	204
rect	65	204	66	205
rect	65	206	66	207
rect	65	207	66	208
rect	65	209	66	210
rect	65	210	66	211
rect	65	212	66	213
rect	65	213	66	214
rect	65	215	66	216
rect	65	216	66	217
rect	65	218	66	219
rect	65	219	66	220
rect	65	221	66	222
rect	65	222	66	223
rect	65	224	66	225
rect	65	225	66	226
rect	65	227	66	228
rect	65	228	66	229
rect	65	230	66	231
rect	65	231	66	232
rect	65	233	66	234
rect	65	234	66	235
rect	65	236	66	237
rect	65	237	66	238
rect	65	239	66	240
rect	65	240	66	241
rect	65	242	66	243
rect	65	243	66	244
rect	65	245	66	246
rect	65	246	66	247
rect	65	248	66	249
rect	65	249	66	250
rect	65	251	66	252
rect	65	252	66	253
rect	65	254	66	255
rect	65	255	66	256
rect	65	257	66	258
rect	65	258	66	259
rect	65	260	66	261
rect	65	261	66	262
rect	65	263	66	264
rect	65	264	66	265
rect	65	266	66	267
rect	65	267	66	268
rect	65	269	66	270
rect	65	270	66	271
rect	65	272	66	273
rect	65	273	66	274
rect	65	275	66	276
rect	65	276	66	277
rect	65	278	66	279
rect	65	279	66	280
rect	65	281	66	282
rect	65	282	66	283
rect	65	284	66	285
rect	65	285	66	286
rect	65	287	66	288
rect	65	288	66	289
rect	65	290	66	291
rect	65	291	66	292
rect	65	293	66	294
rect	65	294	66	295
rect	65	296	66	297
rect	65	297	66	298
rect	65	299	66	300
rect	65	300	66	301
rect	65	302	66	303
rect	65	303	66	304
rect	65	305	66	306
rect	65	306	66	307
rect	65	308	66	309
rect	65	309	66	310
rect	65	311	66	312
rect	67	0	68	1
rect	67	2	68	3
rect	67	3	68	4
rect	67	5	68	6
rect	67	6	68	7
rect	67	8	68	9
rect	67	9	68	10
rect	67	11	68	12
rect	67	12	68	13
rect	67	14	68	15
rect	67	15	68	16
rect	67	17	68	18
rect	67	18	68	19
rect	67	20	68	21
rect	67	21	68	22
rect	67	23	68	24
rect	67	24	68	25
rect	67	26	68	27
rect	67	27	68	28
rect	67	29	68	30
rect	67	30	68	31
rect	67	32	68	33
rect	67	33	68	34
rect	67	35	68	36
rect	67	36	68	37
rect	67	38	68	39
rect	67	39	68	40
rect	67	41	68	42
rect	67	42	68	43
rect	67	44	68	45
rect	67	45	68	46
rect	67	47	68	48
rect	67	48	68	49
rect	67	50	68	51
rect	67	51	68	52
rect	67	53	68	54
rect	67	54	68	55
rect	67	56	68	57
rect	67	57	68	58
rect	67	59	68	60
rect	67	60	68	61
rect	67	62	68	63
rect	67	63	68	64
rect	67	65	68	66
rect	67	66	68	67
rect	67	68	68	69
rect	67	69	68	70
rect	67	71	68	72
rect	67	72	68	73
rect	67	74	68	75
rect	67	75	68	76
rect	67	77	68	78
rect	67	78	68	79
rect	67	80	68	81
rect	67	81	68	82
rect	67	83	68	84
rect	67	84	68	85
rect	67	86	68	87
rect	67	87	68	88
rect	67	89	68	90
rect	67	90	68	91
rect	67	92	68	93
rect	67	93	68	94
rect	67	95	68	96
rect	67	96	68	97
rect	67	98	68	99
rect	67	99	68	100
rect	67	101	68	102
rect	67	102	68	103
rect	67	104	68	105
rect	67	105	68	106
rect	67	107	68	108
rect	67	108	68	109
rect	67	110	68	111
rect	67	111	68	112
rect	67	113	68	114
rect	67	114	68	115
rect	67	116	68	117
rect	67	117	68	118
rect	67	119	68	120
rect	67	120	68	121
rect	67	122	68	123
rect	67	123	68	124
rect	67	125	68	126
rect	67	126	68	127
rect	67	128	68	129
rect	67	129	68	130
rect	67	131	68	132
rect	67	132	68	133
rect	67	134	68	135
rect	67	135	68	136
rect	67	137	68	138
rect	67	138	68	139
rect	67	140	68	141
rect	67	141	68	142
rect	67	143	68	144
rect	67	144	68	145
rect	67	146	68	147
rect	67	147	68	148
rect	67	149	68	150
rect	67	150	68	151
rect	67	152	68	153
rect	67	153	68	154
rect	67	155	68	156
rect	67	156	68	157
rect	67	158	68	159
rect	67	159	68	160
rect	67	161	68	162
rect	67	162	68	163
rect	67	164	68	165
rect	67	165	68	166
rect	67	167	68	168
rect	67	168	68	169
rect	67	170	68	171
rect	67	171	68	172
rect	67	173	68	174
rect	67	174	68	175
rect	67	176	68	177
rect	67	177	68	178
rect	67	179	68	180
rect	67	180	68	181
rect	67	182	68	183
rect	67	183	68	184
rect	67	185	68	186
rect	67	186	68	187
rect	67	188	68	189
rect	67	189	68	190
rect	67	191	68	192
rect	67	192	68	193
rect	67	194	68	195
rect	67	195	68	196
rect	67	197	68	198
rect	67	198	68	199
rect	67	200	68	201
rect	67	201	68	202
rect	67	203	68	204
rect	67	204	68	205
rect	67	206	68	207
rect	67	207	68	208
rect	67	209	68	210
rect	67	210	68	211
rect	67	212	68	213
rect	67	213	68	214
rect	67	215	68	216
rect	67	216	68	217
rect	67	218	68	219
rect	67	219	68	220
rect	67	221	68	222
rect	67	222	68	223
rect	67	224	68	225
rect	67	225	68	226
rect	67	227	68	228
rect	67	228	68	229
rect	67	230	68	231
rect	67	231	68	232
rect	67	233	68	234
rect	67	234	68	235
rect	67	236	68	237
rect	67	237	68	238
rect	67	239	68	240
rect	67	240	68	241
rect	67	242	68	243
rect	67	243	68	244
rect	67	245	68	246
rect	67	246	68	247
rect	67	248	68	249
rect	67	249	68	250
rect	67	251	68	252
rect	67	252	68	253
rect	67	254	68	255
rect	67	255	68	256
rect	67	257	68	258
rect	67	258	68	259
rect	67	260	68	261
rect	67	261	68	262
rect	67	263	68	264
rect	67	264	68	265
rect	67	266	68	267
rect	67	267	68	268
rect	67	269	68	270
rect	67	270	68	271
rect	67	272	68	273
rect	67	273	68	274
rect	67	275	68	276
rect	67	276	68	277
rect	67	278	68	279
rect	67	279	68	280
rect	67	281	68	282
rect	67	282	68	283
rect	67	284	68	285
rect	67	285	68	286
rect	67	287	68	288
rect	67	288	68	289
rect	67	290	68	291
rect	67	291	68	292
rect	67	293	68	294
rect	67	294	68	295
rect	67	296	68	297
rect	67	297	68	298
rect	67	299	68	300
rect	67	300	68	301
rect	67	302	68	303
rect	67	303	68	304
rect	67	305	68	306
rect	67	306	68	307
rect	67	308	68	309
rect	67	309	68	310
rect	67	311	68	312
rect	67	312	68	313
rect	67	314	68	315
rect	67	315	68	316
rect	67	317	68	318
rect	67	318	68	319
rect	67	320	68	321
rect	67	321	68	322
rect	67	323	68	324
rect	68	0	69	1
rect	68	2	69	3
rect	68	3	69	4
rect	68	5	69	6
rect	68	6	69	7
rect	68	8	69	9
rect	68	9	69	10
rect	68	11	69	12
rect	68	12	69	13
rect	68	14	69	15
rect	68	15	69	16
rect	68	17	69	18
rect	68	18	69	19
rect	68	20	69	21
rect	68	21	69	22
rect	68	23	69	24
rect	68	24	69	25
rect	68	26	69	27
rect	68	27	69	28
rect	68	29	69	30
rect	68	30	69	31
rect	68	32	69	33
rect	68	33	69	34
rect	68	35	69	36
rect	68	36	69	37
rect	68	38	69	39
rect	68	39	69	40
rect	68	41	69	42
rect	68	42	69	43
rect	68	44	69	45
rect	68	45	69	46
rect	68	47	69	48
rect	68	48	69	49
rect	68	50	69	51
rect	68	51	69	52
rect	68	53	69	54
rect	68	54	69	55
rect	68	56	69	57
rect	68	57	69	58
rect	68	59	69	60
rect	68	60	69	61
rect	68	62	69	63
rect	68	63	69	64
rect	68	65	69	66
rect	68	66	69	67
rect	68	68	69	69
rect	68	69	69	70
rect	68	71	69	72
rect	68	72	69	73
rect	68	74	69	75
rect	68	75	69	76
rect	68	77	69	78
rect	68	78	69	79
rect	68	80	69	81
rect	68	81	69	82
rect	68	83	69	84
rect	68	84	69	85
rect	68	86	69	87
rect	68	87	69	88
rect	68	89	69	90
rect	68	90	69	91
rect	68	92	69	93
rect	68	93	69	94
rect	68	95	69	96
rect	68	96	69	97
rect	68	98	69	99
rect	68	99	69	100
rect	68	101	69	102
rect	68	102	69	103
rect	68	104	69	105
rect	68	105	69	106
rect	68	107	69	108
rect	68	108	69	109
rect	68	110	69	111
rect	68	111	69	112
rect	68	113	69	114
rect	68	114	69	115
rect	68	116	69	117
rect	68	117	69	118
rect	68	119	69	120
rect	68	120	69	121
rect	68	122	69	123
rect	68	123	69	124
rect	68	125	69	126
rect	68	126	69	127
rect	68	128	69	129
rect	68	129	69	130
rect	68	131	69	132
rect	68	132	69	133
rect	68	134	69	135
rect	68	135	69	136
rect	68	137	69	138
rect	68	138	69	139
rect	68	140	69	141
rect	68	141	69	142
rect	68	143	69	144
rect	68	144	69	145
rect	68	146	69	147
rect	68	147	69	148
rect	68	149	69	150
rect	68	150	69	151
rect	68	152	69	153
rect	68	153	69	154
rect	68	155	69	156
rect	68	156	69	157
rect	68	158	69	159
rect	68	159	69	160
rect	68	161	69	162
rect	68	162	69	163
rect	68	164	69	165
rect	68	165	69	166
rect	68	167	69	168
rect	68	168	69	169
rect	68	170	69	171
rect	68	171	69	172
rect	68	173	69	174
rect	68	174	69	175
rect	68	176	69	177
rect	68	177	69	178
rect	68	179	69	180
rect	68	180	69	181
rect	68	182	69	183
rect	68	183	69	184
rect	68	185	69	186
rect	68	186	69	187
rect	68	188	69	189
rect	68	189	69	190
rect	68	191	69	192
rect	68	192	69	193
rect	68	194	69	195
rect	68	195	69	196
rect	68	197	69	198
rect	68	198	69	199
rect	68	200	69	201
rect	68	201	69	202
rect	68	203	69	204
rect	68	204	69	205
rect	68	206	69	207
rect	68	207	69	208
rect	68	209	69	210
rect	68	210	69	211
rect	68	212	69	213
rect	68	213	69	214
rect	68	215	69	216
rect	68	216	69	217
rect	68	218	69	219
rect	68	219	69	220
rect	68	221	69	222
rect	68	222	69	223
rect	68	224	69	225
rect	68	225	69	226
rect	68	227	69	228
rect	68	228	69	229
rect	68	230	69	231
rect	68	231	69	232
rect	68	233	69	234
rect	68	234	69	235
rect	68	236	69	237
rect	68	237	69	238
rect	68	239	69	240
rect	68	240	69	241
rect	68	242	69	243
rect	68	243	69	244
rect	68	245	69	246
rect	68	246	69	247
rect	68	248	69	249
rect	68	249	69	250
rect	68	251	69	252
rect	68	252	69	253
rect	68	254	69	255
rect	68	255	69	256
rect	68	257	69	258
rect	68	258	69	259
rect	68	260	69	261
rect	68	261	69	262
rect	68	263	69	264
rect	68	264	69	265
rect	68	266	69	267
rect	68	267	69	268
rect	68	269	69	270
rect	68	270	69	271
rect	68	272	69	273
rect	68	273	69	274
rect	68	275	69	276
rect	68	276	69	277
rect	68	278	69	279
rect	68	279	69	280
rect	68	281	69	282
rect	68	282	69	283
rect	68	284	69	285
rect	68	285	69	286
rect	68	287	69	288
rect	68	288	69	289
rect	68	290	69	291
rect	68	291	69	292
rect	68	293	69	294
rect	68	294	69	295
rect	68	296	69	297
rect	68	297	69	298
rect	68	299	69	300
rect	68	300	69	301
rect	68	302	69	303
rect	68	303	69	304
rect	68	305	69	306
rect	68	306	69	307
rect	68	308	69	309
rect	68	309	69	310
rect	68	311	69	312
rect	68	312	69	313
rect	68	314	69	315
rect	68	315	69	316
rect	68	317	69	318
rect	68	318	69	319
rect	68	320	69	321
rect	68	321	69	322
rect	68	323	69	324
rect	69	0	70	1
rect	69	2	70	3
rect	69	3	70	4
rect	69	5	70	6
rect	69	6	70	7
rect	69	8	70	9
rect	69	9	70	10
rect	69	11	70	12
rect	69	12	70	13
rect	69	14	70	15
rect	69	15	70	16
rect	69	17	70	18
rect	69	18	70	19
rect	69	20	70	21
rect	69	21	70	22
rect	69	23	70	24
rect	69	24	70	25
rect	69	26	70	27
rect	69	27	70	28
rect	69	29	70	30
rect	69	30	70	31
rect	69	32	70	33
rect	69	33	70	34
rect	69	35	70	36
rect	69	36	70	37
rect	69	38	70	39
rect	69	39	70	40
rect	69	41	70	42
rect	69	42	70	43
rect	69	44	70	45
rect	69	45	70	46
rect	69	47	70	48
rect	69	48	70	49
rect	69	50	70	51
rect	69	51	70	52
rect	69	53	70	54
rect	69	54	70	55
rect	69	56	70	57
rect	69	57	70	58
rect	69	59	70	60
rect	69	60	70	61
rect	69	62	70	63
rect	69	63	70	64
rect	69	65	70	66
rect	69	66	70	67
rect	69	68	70	69
rect	69	69	70	70
rect	69	71	70	72
rect	69	72	70	73
rect	69	74	70	75
rect	69	75	70	76
rect	69	77	70	78
rect	69	78	70	79
rect	69	80	70	81
rect	69	81	70	82
rect	69	83	70	84
rect	69	84	70	85
rect	69	86	70	87
rect	69	87	70	88
rect	69	89	70	90
rect	69	90	70	91
rect	69	92	70	93
rect	69	93	70	94
rect	69	95	70	96
rect	69	96	70	97
rect	69	98	70	99
rect	69	99	70	100
rect	69	101	70	102
rect	69	102	70	103
rect	69	104	70	105
rect	69	105	70	106
rect	69	107	70	108
rect	69	108	70	109
rect	69	110	70	111
rect	69	111	70	112
rect	69	113	70	114
rect	69	114	70	115
rect	69	116	70	117
rect	69	117	70	118
rect	69	119	70	120
rect	69	120	70	121
rect	69	122	70	123
rect	69	123	70	124
rect	69	125	70	126
rect	69	126	70	127
rect	69	128	70	129
rect	69	129	70	130
rect	69	131	70	132
rect	69	132	70	133
rect	69	134	70	135
rect	69	135	70	136
rect	69	137	70	138
rect	69	138	70	139
rect	69	140	70	141
rect	69	141	70	142
rect	69	143	70	144
rect	69	144	70	145
rect	69	146	70	147
rect	69	147	70	148
rect	69	149	70	150
rect	69	150	70	151
rect	69	152	70	153
rect	69	153	70	154
rect	69	155	70	156
rect	69	156	70	157
rect	69	158	70	159
rect	69	159	70	160
rect	69	161	70	162
rect	69	162	70	163
rect	69	164	70	165
rect	69	165	70	166
rect	69	167	70	168
rect	69	168	70	169
rect	69	170	70	171
rect	69	171	70	172
rect	69	173	70	174
rect	69	174	70	175
rect	69	176	70	177
rect	69	177	70	178
rect	69	179	70	180
rect	69	180	70	181
rect	69	182	70	183
rect	69	183	70	184
rect	69	185	70	186
rect	69	186	70	187
rect	69	188	70	189
rect	69	189	70	190
rect	69	191	70	192
rect	69	192	70	193
rect	69	194	70	195
rect	69	195	70	196
rect	69	197	70	198
rect	69	198	70	199
rect	69	200	70	201
rect	69	201	70	202
rect	69	203	70	204
rect	69	204	70	205
rect	69	206	70	207
rect	69	207	70	208
rect	69	209	70	210
rect	69	210	70	211
rect	69	212	70	213
rect	69	213	70	214
rect	69	215	70	216
rect	69	216	70	217
rect	69	218	70	219
rect	69	219	70	220
rect	69	221	70	222
rect	69	222	70	223
rect	69	224	70	225
rect	69	225	70	226
rect	69	227	70	228
rect	69	228	70	229
rect	69	230	70	231
rect	69	231	70	232
rect	69	233	70	234
rect	69	234	70	235
rect	69	236	70	237
rect	69	237	70	238
rect	69	239	70	240
rect	69	240	70	241
rect	69	242	70	243
rect	69	243	70	244
rect	69	245	70	246
rect	69	246	70	247
rect	69	248	70	249
rect	69	249	70	250
rect	69	251	70	252
rect	69	252	70	253
rect	69	254	70	255
rect	69	255	70	256
rect	69	257	70	258
rect	69	258	70	259
rect	69	260	70	261
rect	69	261	70	262
rect	69	263	70	264
rect	69	264	70	265
rect	69	266	70	267
rect	69	267	70	268
rect	69	269	70	270
rect	69	270	70	271
rect	69	272	70	273
rect	69	273	70	274
rect	69	275	70	276
rect	69	276	70	277
rect	69	278	70	279
rect	69	279	70	280
rect	69	281	70	282
rect	69	282	70	283
rect	69	284	70	285
rect	69	285	70	286
rect	69	287	70	288
rect	69	288	70	289
rect	69	290	70	291
rect	69	291	70	292
rect	69	293	70	294
rect	69	294	70	295
rect	69	296	70	297
rect	69	297	70	298
rect	69	299	70	300
rect	69	300	70	301
rect	69	302	70	303
rect	69	303	70	304
rect	69	305	70	306
rect	69	306	70	307
rect	69	308	70	309
rect	69	309	70	310
rect	69	311	70	312
rect	69	312	70	313
rect	69	314	70	315
rect	69	315	70	316
rect	69	317	70	318
rect	69	318	70	319
rect	69	320	70	321
rect	69	321	70	322
rect	69	323	70	324
rect	70	0	71	1
rect	70	2	71	3
rect	70	3	71	4
rect	70	5	71	6
rect	70	6	71	7
rect	70	8	71	9
rect	70	9	71	10
rect	70	11	71	12
rect	70	12	71	13
rect	70	14	71	15
rect	70	15	71	16
rect	70	17	71	18
rect	70	18	71	19
rect	70	20	71	21
rect	70	21	71	22
rect	70	23	71	24
rect	70	24	71	25
rect	70	26	71	27
rect	70	27	71	28
rect	70	29	71	30
rect	70	30	71	31
rect	70	32	71	33
rect	70	33	71	34
rect	70	35	71	36
rect	70	36	71	37
rect	70	38	71	39
rect	70	39	71	40
rect	70	41	71	42
rect	70	42	71	43
rect	70	44	71	45
rect	70	45	71	46
rect	70	47	71	48
rect	70	48	71	49
rect	70	50	71	51
rect	70	51	71	52
rect	70	53	71	54
rect	70	54	71	55
rect	70	56	71	57
rect	70	57	71	58
rect	70	59	71	60
rect	70	60	71	61
rect	70	62	71	63
rect	70	63	71	64
rect	70	65	71	66
rect	70	66	71	67
rect	70	68	71	69
rect	70	69	71	70
rect	70	71	71	72
rect	70	72	71	73
rect	70	74	71	75
rect	70	75	71	76
rect	70	77	71	78
rect	70	78	71	79
rect	70	80	71	81
rect	70	81	71	82
rect	70	83	71	84
rect	70	84	71	85
rect	70	86	71	87
rect	70	87	71	88
rect	70	89	71	90
rect	70	90	71	91
rect	70	92	71	93
rect	70	93	71	94
rect	70	95	71	96
rect	70	96	71	97
rect	70	98	71	99
rect	70	99	71	100
rect	70	101	71	102
rect	70	102	71	103
rect	70	104	71	105
rect	70	105	71	106
rect	70	107	71	108
rect	70	108	71	109
rect	70	110	71	111
rect	70	111	71	112
rect	70	113	71	114
rect	70	114	71	115
rect	70	116	71	117
rect	70	117	71	118
rect	70	119	71	120
rect	70	120	71	121
rect	70	122	71	123
rect	70	123	71	124
rect	70	125	71	126
rect	70	126	71	127
rect	70	128	71	129
rect	70	129	71	130
rect	70	131	71	132
rect	70	132	71	133
rect	70	134	71	135
rect	70	135	71	136
rect	70	137	71	138
rect	70	138	71	139
rect	70	140	71	141
rect	70	141	71	142
rect	70	143	71	144
rect	70	144	71	145
rect	70	146	71	147
rect	70	147	71	148
rect	70	149	71	150
rect	70	150	71	151
rect	70	152	71	153
rect	70	153	71	154
rect	70	155	71	156
rect	70	156	71	157
rect	70	158	71	159
rect	70	159	71	160
rect	70	161	71	162
rect	70	162	71	163
rect	70	164	71	165
rect	70	165	71	166
rect	70	167	71	168
rect	70	168	71	169
rect	70	170	71	171
rect	70	171	71	172
rect	70	173	71	174
rect	70	174	71	175
rect	70	176	71	177
rect	70	177	71	178
rect	70	179	71	180
rect	70	180	71	181
rect	70	182	71	183
rect	70	183	71	184
rect	70	185	71	186
rect	70	186	71	187
rect	70	188	71	189
rect	70	189	71	190
rect	70	191	71	192
rect	70	192	71	193
rect	70	194	71	195
rect	70	195	71	196
rect	70	197	71	198
rect	70	198	71	199
rect	70	200	71	201
rect	70	201	71	202
rect	70	203	71	204
rect	70	204	71	205
rect	70	206	71	207
rect	70	207	71	208
rect	70	209	71	210
rect	70	210	71	211
rect	70	212	71	213
rect	70	213	71	214
rect	70	215	71	216
rect	70	216	71	217
rect	70	218	71	219
rect	70	219	71	220
rect	70	221	71	222
rect	70	222	71	223
rect	70	224	71	225
rect	70	225	71	226
rect	70	227	71	228
rect	70	228	71	229
rect	70	230	71	231
rect	70	231	71	232
rect	70	233	71	234
rect	70	234	71	235
rect	70	236	71	237
rect	70	237	71	238
rect	70	239	71	240
rect	70	240	71	241
rect	70	242	71	243
rect	70	243	71	244
rect	70	245	71	246
rect	70	246	71	247
rect	70	248	71	249
rect	70	249	71	250
rect	70	251	71	252
rect	70	252	71	253
rect	70	254	71	255
rect	70	255	71	256
rect	70	257	71	258
rect	70	258	71	259
rect	70	260	71	261
rect	70	261	71	262
rect	70	263	71	264
rect	70	264	71	265
rect	70	266	71	267
rect	70	267	71	268
rect	70	269	71	270
rect	70	270	71	271
rect	70	272	71	273
rect	70	273	71	274
rect	70	275	71	276
rect	70	276	71	277
rect	70	278	71	279
rect	70	279	71	280
rect	70	281	71	282
rect	70	282	71	283
rect	70	284	71	285
rect	70	285	71	286
rect	70	287	71	288
rect	70	288	71	289
rect	70	290	71	291
rect	70	291	71	292
rect	70	293	71	294
rect	70	294	71	295
rect	70	296	71	297
rect	70	297	71	298
rect	70	299	71	300
rect	70	300	71	301
rect	70	302	71	303
rect	70	303	71	304
rect	70	305	71	306
rect	70	306	71	307
rect	70	308	71	309
rect	70	309	71	310
rect	70	311	71	312
rect	70	312	71	313
rect	70	314	71	315
rect	70	315	71	316
rect	70	317	71	318
rect	70	318	71	319
rect	70	320	71	321
rect	70	321	71	322
rect	70	323	71	324
rect	71	0	72	1
rect	71	2	72	3
rect	71	3	72	4
rect	71	5	72	6
rect	71	6	72	7
rect	71	8	72	9
rect	71	9	72	10
rect	71	11	72	12
rect	71	12	72	13
rect	71	14	72	15
rect	71	15	72	16
rect	71	17	72	18
rect	71	18	72	19
rect	71	20	72	21
rect	71	21	72	22
rect	71	23	72	24
rect	71	24	72	25
rect	71	26	72	27
rect	71	27	72	28
rect	71	29	72	30
rect	71	30	72	31
rect	71	32	72	33
rect	71	33	72	34
rect	71	35	72	36
rect	71	36	72	37
rect	71	38	72	39
rect	71	39	72	40
rect	71	41	72	42
rect	71	42	72	43
rect	71	44	72	45
rect	71	45	72	46
rect	71	47	72	48
rect	71	48	72	49
rect	71	50	72	51
rect	71	51	72	52
rect	71	53	72	54
rect	71	54	72	55
rect	71	56	72	57
rect	71	57	72	58
rect	71	59	72	60
rect	71	60	72	61
rect	71	62	72	63
rect	71	63	72	64
rect	71	65	72	66
rect	71	66	72	67
rect	71	68	72	69
rect	71	69	72	70
rect	71	71	72	72
rect	71	72	72	73
rect	71	74	72	75
rect	71	75	72	76
rect	71	77	72	78
rect	71	78	72	79
rect	71	80	72	81
rect	71	81	72	82
rect	71	83	72	84
rect	71	84	72	85
rect	71	86	72	87
rect	71	87	72	88
rect	71	89	72	90
rect	71	90	72	91
rect	71	92	72	93
rect	71	93	72	94
rect	71	95	72	96
rect	71	96	72	97
rect	71	98	72	99
rect	71	99	72	100
rect	71	101	72	102
rect	71	102	72	103
rect	71	104	72	105
rect	71	105	72	106
rect	71	107	72	108
rect	71	108	72	109
rect	71	110	72	111
rect	71	111	72	112
rect	71	113	72	114
rect	71	114	72	115
rect	71	116	72	117
rect	71	117	72	118
rect	71	119	72	120
rect	71	120	72	121
rect	71	122	72	123
rect	71	123	72	124
rect	71	125	72	126
rect	71	126	72	127
rect	71	128	72	129
rect	71	129	72	130
rect	71	131	72	132
rect	71	132	72	133
rect	71	134	72	135
rect	71	135	72	136
rect	71	137	72	138
rect	71	138	72	139
rect	71	140	72	141
rect	71	141	72	142
rect	71	143	72	144
rect	71	144	72	145
rect	71	146	72	147
rect	71	147	72	148
rect	71	149	72	150
rect	71	150	72	151
rect	71	152	72	153
rect	71	153	72	154
rect	71	155	72	156
rect	71	156	72	157
rect	71	158	72	159
rect	71	159	72	160
rect	71	161	72	162
rect	71	162	72	163
rect	71	164	72	165
rect	71	165	72	166
rect	71	167	72	168
rect	71	168	72	169
rect	71	170	72	171
rect	71	171	72	172
rect	71	173	72	174
rect	71	174	72	175
rect	71	176	72	177
rect	71	177	72	178
rect	71	179	72	180
rect	71	180	72	181
rect	71	182	72	183
rect	71	183	72	184
rect	71	185	72	186
rect	71	186	72	187
rect	71	188	72	189
rect	71	189	72	190
rect	71	191	72	192
rect	71	192	72	193
rect	71	194	72	195
rect	71	195	72	196
rect	71	197	72	198
rect	71	198	72	199
rect	71	200	72	201
rect	71	201	72	202
rect	71	203	72	204
rect	71	204	72	205
rect	71	206	72	207
rect	71	207	72	208
rect	71	209	72	210
rect	71	210	72	211
rect	71	212	72	213
rect	71	213	72	214
rect	71	215	72	216
rect	71	216	72	217
rect	71	218	72	219
rect	71	219	72	220
rect	71	221	72	222
rect	71	222	72	223
rect	71	224	72	225
rect	71	225	72	226
rect	71	227	72	228
rect	71	228	72	229
rect	71	230	72	231
rect	71	231	72	232
rect	71	233	72	234
rect	71	234	72	235
rect	71	236	72	237
rect	71	237	72	238
rect	71	239	72	240
rect	71	240	72	241
rect	71	242	72	243
rect	71	243	72	244
rect	71	245	72	246
rect	71	246	72	247
rect	71	248	72	249
rect	71	249	72	250
rect	71	251	72	252
rect	71	252	72	253
rect	71	254	72	255
rect	71	255	72	256
rect	71	257	72	258
rect	71	258	72	259
rect	71	260	72	261
rect	71	261	72	262
rect	71	263	72	264
rect	71	264	72	265
rect	71	266	72	267
rect	71	267	72	268
rect	71	269	72	270
rect	71	270	72	271
rect	71	272	72	273
rect	71	273	72	274
rect	71	275	72	276
rect	71	276	72	277
rect	71	278	72	279
rect	71	279	72	280
rect	71	281	72	282
rect	71	282	72	283
rect	71	284	72	285
rect	71	285	72	286
rect	71	287	72	288
rect	71	288	72	289
rect	71	290	72	291
rect	71	291	72	292
rect	71	293	72	294
rect	71	294	72	295
rect	71	296	72	297
rect	71	297	72	298
rect	71	299	72	300
rect	71	300	72	301
rect	71	302	72	303
rect	71	303	72	304
rect	71	305	72	306
rect	71	306	72	307
rect	71	308	72	309
rect	71	309	72	310
rect	71	311	72	312
rect	71	312	72	313
rect	71	314	72	315
rect	71	315	72	316
rect	71	317	72	318
rect	71	318	72	319
rect	71	320	72	321
rect	71	321	72	322
rect	71	323	72	324
rect	80	0	81	1
rect	80	2	81	3
rect	80	3	81	4
rect	80	5	81	6
rect	80	6	81	7
rect	80	8	81	9
rect	80	9	81	10
rect	80	11	81	12
rect	80	12	81	13
rect	80	14	81	15
rect	80	15	81	16
rect	80	17	81	18
rect	80	18	81	19
rect	80	20	81	21
rect	80	21	81	22
rect	80	23	81	24
rect	80	24	81	25
rect	80	26	81	27
rect	80	27	81	28
rect	80	29	81	30
rect	80	30	81	31
rect	80	32	81	33
rect	80	33	81	34
rect	80	35	81	36
rect	80	36	81	37
rect	80	38	81	39
rect	80	39	81	40
rect	80	41	81	42
rect	80	42	81	43
rect	80	44	81	45
rect	80	45	81	46
rect	80	47	81	48
rect	80	48	81	49
rect	80	50	81	51
rect	80	51	81	52
rect	80	53	81	54
rect	80	54	81	55
rect	80	56	81	57
rect	80	57	81	58
rect	80	59	81	60
rect	80	60	81	61
rect	80	62	81	63
rect	80	63	81	64
rect	80	65	81	66
rect	80	66	81	67
rect	80	68	81	69
rect	80	69	81	70
rect	80	71	81	72
rect	80	72	81	73
rect	80	74	81	75
rect	80	75	81	76
rect	80	77	81	78
rect	80	78	81	79
rect	80	80	81	81
rect	80	81	81	82
rect	80	83	81	84
rect	80	84	81	85
rect	80	86	81	87
rect	80	87	81	88
rect	80	89	81	90
rect	80	90	81	91
rect	80	92	81	93
rect	80	93	81	94
rect	80	95	81	96
rect	80	96	81	97
rect	80	98	81	99
rect	80	99	81	100
rect	80	101	81	102
rect	80	102	81	103
rect	80	104	81	105
rect	80	105	81	106
rect	80	107	81	108
rect	80	108	81	109
rect	80	110	81	111
rect	80	111	81	112
rect	80	113	81	114
rect	80	114	81	115
rect	80	116	81	117
rect	80	117	81	118
rect	80	119	81	120
rect	80	120	81	121
rect	80	122	81	123
rect	80	123	81	124
rect	80	125	81	126
rect	80	126	81	127
rect	80	128	81	129
rect	80	129	81	130
rect	80	131	81	132
rect	80	132	81	133
rect	80	134	81	135
rect	80	135	81	136
rect	80	137	81	138
rect	80	138	81	139
rect	80	140	81	141
rect	80	141	81	142
rect	80	143	81	144
rect	80	144	81	145
rect	80	146	81	147
rect	80	147	81	148
rect	80	149	81	150
rect	80	150	81	151
rect	80	152	81	153
rect	80	153	81	154
rect	80	155	81	156
rect	80	156	81	157
rect	80	158	81	159
rect	80	159	81	160
rect	80	161	81	162
rect	80	162	81	163
rect	80	164	81	165
rect	80	165	81	166
rect	80	167	81	168
rect	80	168	81	169
rect	80	170	81	171
rect	80	171	81	172
rect	80	173	81	174
rect	80	174	81	175
rect	80	176	81	177
rect	80	177	81	178
rect	80	179	81	180
rect	80	180	81	181
rect	80	182	81	183
rect	80	183	81	184
rect	80	185	81	186
rect	80	186	81	187
rect	80	188	81	189
rect	80	189	81	190
rect	80	191	81	192
rect	80	192	81	193
rect	80	194	81	195
rect	80	195	81	196
rect	80	197	81	198
rect	80	198	81	199
rect	80	200	81	201
rect	80	201	81	202
rect	80	203	81	204
rect	80	204	81	205
rect	80	206	81	207
rect	80	207	81	208
rect	80	209	81	210
rect	80	210	81	211
rect	80	212	81	213
rect	80	213	81	214
rect	80	215	81	216
rect	80	216	81	217
rect	80	218	81	219
rect	80	219	81	220
rect	80	221	81	222
rect	80	222	81	223
rect	80	224	81	225
rect	80	225	81	226
rect	80	227	81	228
rect	80	228	81	229
rect	80	230	81	231
rect	80	231	81	232
rect	80	233	81	234
rect	80	234	81	235
rect	80	236	81	237
rect	80	237	81	238
rect	80	239	81	240
rect	80	240	81	241
rect	80	242	81	243
rect	80	243	81	244
rect	80	245	81	246
rect	80	246	81	247
rect	80	248	81	249
rect	80	249	81	250
rect	80	251	81	252
rect	80	252	81	253
rect	80	254	81	255
rect	80	255	81	256
rect	80	257	81	258
rect	80	258	81	259
rect	80	260	81	261
rect	80	261	81	262
rect	80	263	81	264
rect	80	264	81	265
rect	80	266	81	267
rect	80	267	81	268
rect	80	269	81	270
rect	80	270	81	271
rect	80	272	81	273
rect	80	273	81	274
rect	80	275	81	276
rect	80	276	81	277
rect	80	278	81	279
rect	80	279	81	280
rect	80	281	81	282
rect	80	282	81	283
rect	80	284	81	285
rect	80	285	81	286
rect	80	287	81	288
rect	80	288	81	289
rect	80	290	81	291
rect	80	291	81	292
rect	80	293	81	294
rect	80	294	81	295
rect	80	296	81	297
rect	80	297	81	298
rect	80	299	81	300
rect	80	300	81	301
rect	80	302	81	303
rect	80	303	81	304
rect	80	305	81	306
rect	80	306	81	307
rect	80	308	81	309
rect	80	309	81	310
rect	80	311	81	312
rect	80	312	81	313
rect	80	314	81	315
rect	80	315	81	316
rect	80	317	81	318
rect	80	318	81	319
rect	80	320	81	321
rect	80	321	81	322
rect	80	323	81	324
rect	82	0	83	1
rect	82	2	83	3
rect	82	3	83	4
rect	82	5	83	6
rect	82	6	83	7
rect	82	8	83	9
rect	82	9	83	10
rect	82	11	83	12
rect	82	12	83	13
rect	82	14	83	15
rect	82	15	83	16
rect	82	17	83	18
rect	82	18	83	19
rect	82	20	83	21
rect	82	21	83	22
rect	82	23	83	24
rect	82	24	83	25
rect	82	26	83	27
rect	82	27	83	28
rect	82	29	83	30
rect	82	30	83	31
rect	82	32	83	33
rect	82	33	83	34
rect	82	35	83	36
rect	82	36	83	37
rect	82	38	83	39
rect	82	39	83	40
rect	82	41	83	42
rect	82	42	83	43
rect	82	44	83	45
rect	82	45	83	46
rect	82	47	83	48
rect	82	48	83	49
rect	82	50	83	51
rect	82	51	83	52
rect	82	53	83	54
rect	82	54	83	55
rect	82	56	83	57
rect	82	57	83	58
rect	82	59	83	60
rect	82	60	83	61
rect	82	62	83	63
rect	82	63	83	64
rect	82	65	83	66
rect	82	66	83	67
rect	82	68	83	69
rect	82	69	83	70
rect	82	71	83	72
rect	82	72	83	73
rect	82	74	83	75
rect	82	75	83	76
rect	82	77	83	78
rect	82	78	83	79
rect	82	80	83	81
rect	82	81	83	82
rect	82	83	83	84
rect	82	84	83	85
rect	82	86	83	87
rect	82	87	83	88
rect	82	89	83	90
rect	82	90	83	91
rect	82	92	83	93
rect	82	93	83	94
rect	82	95	83	96
rect	82	96	83	97
rect	82	98	83	99
rect	82	99	83	100
rect	82	101	83	102
rect	82	102	83	103
rect	82	104	83	105
rect	82	105	83	106
rect	82	107	83	108
rect	82	108	83	109
rect	82	110	83	111
rect	82	111	83	112
rect	82	113	83	114
rect	82	114	83	115
rect	82	116	83	117
rect	82	117	83	118
rect	82	119	83	120
rect	82	120	83	121
rect	82	122	83	123
rect	82	123	83	124
rect	82	125	83	126
rect	82	126	83	127
rect	82	128	83	129
rect	82	129	83	130
rect	82	131	83	132
rect	82	132	83	133
rect	82	134	83	135
rect	82	135	83	136
rect	82	137	83	138
rect	82	138	83	139
rect	82	140	83	141
rect	82	141	83	142
rect	82	143	83	144
rect	82	144	83	145
rect	82	146	83	147
rect	82	147	83	148
rect	82	149	83	150
rect	82	150	83	151
rect	82	152	83	153
rect	82	153	83	154
rect	82	155	83	156
rect	82	156	83	157
rect	82	158	83	159
rect	82	159	83	160
rect	82	161	83	162
rect	82	162	83	163
rect	82	164	83	165
rect	82	165	83	166
rect	82	167	83	168
rect	82	168	83	169
rect	82	170	83	171
rect	82	171	83	172
rect	82	173	83	174
rect	82	174	83	175
rect	82	176	83	177
rect	82	177	83	178
rect	82	179	83	180
rect	82	180	83	181
rect	82	182	83	183
rect	82	183	83	184
rect	82	185	83	186
rect	82	186	83	187
rect	82	188	83	189
rect	82	189	83	190
rect	82	191	83	192
rect	82	192	83	193
rect	82	194	83	195
rect	82	195	83	196
rect	82	197	83	198
rect	82	198	83	199
rect	82	200	83	201
rect	82	201	83	202
rect	82	203	83	204
rect	82	204	83	205
rect	82	206	83	207
rect	82	207	83	208
rect	82	209	83	210
rect	82	210	83	211
rect	82	212	83	213
rect	82	213	83	214
rect	82	215	83	216
rect	82	216	83	217
rect	82	218	83	219
rect	82	219	83	220
rect	82	221	83	222
rect	82	222	83	223
rect	82	224	83	225
rect	82	225	83	226
rect	82	227	83	228
rect	82	228	83	229
rect	82	230	83	231
rect	82	231	83	232
rect	82	233	83	234
rect	82	234	83	235
rect	82	236	83	237
rect	82	237	83	238
rect	82	239	83	240
rect	82	240	83	241
rect	82	242	83	243
rect	82	243	83	244
rect	82	245	83	246
rect	82	246	83	247
rect	82	248	83	249
rect	82	249	83	250
rect	82	251	83	252
rect	82	252	83	253
rect	82	254	83	255
rect	82	255	83	256
rect	82	257	83	258
rect	82	258	83	259
rect	82	260	83	261
rect	82	261	83	262
rect	82	263	83	264
rect	82	264	83	265
rect	82	266	83	267
rect	82	267	83	268
rect	82	269	83	270
rect	82	270	83	271
rect	82	272	83	273
rect	82	273	83	274
rect	82	275	83	276
rect	82	276	83	277
rect	82	278	83	279
rect	82	279	83	280
rect	82	281	83	282
rect	82	282	83	283
rect	82	284	83	285
rect	82	285	83	286
rect	82	287	83	288
rect	82	288	83	289
rect	82	290	83	291
rect	82	291	83	292
rect	82	293	83	294
rect	82	294	83	295
rect	82	296	83	297
rect	82	297	83	298
rect	82	299	83	300
rect	82	300	83	301
rect	82	302	83	303
rect	82	303	83	304
rect	82	305	83	306
rect	82	306	83	307
rect	82	308	83	309
rect	82	309	83	310
rect	82	311	83	312
rect	82	312	83	313
rect	82	314	83	315
rect	82	315	83	316
rect	82	317	83	318
rect	82	318	83	319
rect	82	320	83	321
rect	82	321	83	322
rect	82	323	83	324
rect	82	324	83	325
rect	82	326	83	327
rect	82	327	83	328
rect	82	329	83	330
rect	83	0	84	1
rect	83	2	84	3
rect	83	3	84	4
rect	83	5	84	6
rect	83	6	84	7
rect	83	8	84	9
rect	83	9	84	10
rect	83	11	84	12
rect	83	12	84	13
rect	83	14	84	15
rect	83	15	84	16
rect	83	17	84	18
rect	83	18	84	19
rect	83	20	84	21
rect	83	21	84	22
rect	83	23	84	24
rect	83	24	84	25
rect	83	26	84	27
rect	83	27	84	28
rect	83	29	84	30
rect	83	30	84	31
rect	83	32	84	33
rect	83	33	84	34
rect	83	35	84	36
rect	83	36	84	37
rect	83	38	84	39
rect	83	39	84	40
rect	83	41	84	42
rect	83	42	84	43
rect	83	44	84	45
rect	83	45	84	46
rect	83	47	84	48
rect	83	48	84	49
rect	83	50	84	51
rect	83	51	84	52
rect	83	53	84	54
rect	83	54	84	55
rect	83	56	84	57
rect	83	57	84	58
rect	83	59	84	60
rect	83	60	84	61
rect	83	62	84	63
rect	83	63	84	64
rect	83	65	84	66
rect	83	66	84	67
rect	83	68	84	69
rect	83	69	84	70
rect	83	71	84	72
rect	83	72	84	73
rect	83	74	84	75
rect	83	75	84	76
rect	83	77	84	78
rect	83	78	84	79
rect	83	80	84	81
rect	83	81	84	82
rect	83	83	84	84
rect	83	84	84	85
rect	83	86	84	87
rect	83	87	84	88
rect	83	89	84	90
rect	83	90	84	91
rect	83	92	84	93
rect	83	93	84	94
rect	83	95	84	96
rect	83	96	84	97
rect	83	98	84	99
rect	83	99	84	100
rect	83	101	84	102
rect	83	102	84	103
rect	83	104	84	105
rect	83	105	84	106
rect	83	107	84	108
rect	83	108	84	109
rect	83	110	84	111
rect	83	111	84	112
rect	83	113	84	114
rect	83	114	84	115
rect	83	116	84	117
rect	83	117	84	118
rect	83	119	84	120
rect	83	120	84	121
rect	83	122	84	123
rect	83	123	84	124
rect	83	125	84	126
rect	83	126	84	127
rect	83	128	84	129
rect	83	129	84	130
rect	83	131	84	132
rect	83	132	84	133
rect	83	134	84	135
rect	83	135	84	136
rect	83	137	84	138
rect	83	138	84	139
rect	83	140	84	141
rect	83	141	84	142
rect	83	143	84	144
rect	83	144	84	145
rect	83	146	84	147
rect	83	147	84	148
rect	83	149	84	150
rect	83	150	84	151
rect	83	152	84	153
rect	83	153	84	154
rect	83	155	84	156
rect	83	156	84	157
rect	83	158	84	159
rect	83	159	84	160
rect	83	161	84	162
rect	83	162	84	163
rect	83	164	84	165
rect	83	165	84	166
rect	83	167	84	168
rect	83	168	84	169
rect	83	170	84	171
rect	83	171	84	172
rect	83	173	84	174
rect	83	174	84	175
rect	83	176	84	177
rect	83	177	84	178
rect	83	179	84	180
rect	83	180	84	181
rect	83	182	84	183
rect	83	183	84	184
rect	83	185	84	186
rect	83	186	84	187
rect	83	188	84	189
rect	83	189	84	190
rect	83	191	84	192
rect	83	192	84	193
rect	83	194	84	195
rect	83	195	84	196
rect	83	197	84	198
rect	83	198	84	199
rect	83	200	84	201
rect	83	201	84	202
rect	83	203	84	204
rect	83	204	84	205
rect	83	206	84	207
rect	83	207	84	208
rect	83	209	84	210
rect	83	210	84	211
rect	83	212	84	213
rect	83	213	84	214
rect	83	215	84	216
rect	83	216	84	217
rect	83	218	84	219
rect	83	219	84	220
rect	83	221	84	222
rect	83	222	84	223
rect	83	224	84	225
rect	83	225	84	226
rect	83	227	84	228
rect	83	228	84	229
rect	83	230	84	231
rect	83	231	84	232
rect	83	233	84	234
rect	83	234	84	235
rect	83	236	84	237
rect	83	237	84	238
rect	83	239	84	240
rect	83	240	84	241
rect	83	242	84	243
rect	83	243	84	244
rect	83	245	84	246
rect	83	246	84	247
rect	83	248	84	249
rect	83	249	84	250
rect	83	251	84	252
rect	83	252	84	253
rect	83	254	84	255
rect	83	255	84	256
rect	83	257	84	258
rect	83	258	84	259
rect	83	260	84	261
rect	83	261	84	262
rect	83	263	84	264
rect	83	264	84	265
rect	83	266	84	267
rect	83	267	84	268
rect	83	269	84	270
rect	83	270	84	271
rect	83	272	84	273
rect	83	273	84	274
rect	83	275	84	276
rect	83	276	84	277
rect	83	278	84	279
rect	83	279	84	280
rect	83	281	84	282
rect	83	282	84	283
rect	83	284	84	285
rect	83	285	84	286
rect	83	287	84	288
rect	83	288	84	289
rect	83	290	84	291
rect	83	291	84	292
rect	83	293	84	294
rect	83	294	84	295
rect	83	296	84	297
rect	83	297	84	298
rect	83	299	84	300
rect	83	300	84	301
rect	83	302	84	303
rect	83	303	84	304
rect	83	305	84	306
rect	83	306	84	307
rect	83	308	84	309
rect	83	309	84	310
rect	83	311	84	312
rect	83	312	84	313
rect	83	314	84	315
rect	83	315	84	316
rect	83	317	84	318
rect	83	318	84	319
rect	83	320	84	321
rect	83	321	84	322
rect	83	323	84	324
rect	83	324	84	325
rect	83	326	84	327
rect	83	327	84	328
rect	83	329	84	330
rect	84	0	85	1
rect	84	2	85	3
rect	84	3	85	4
rect	84	5	85	6
rect	84	6	85	7
rect	84	8	85	9
rect	84	9	85	10
rect	84	11	85	12
rect	84	12	85	13
rect	84	14	85	15
rect	84	15	85	16
rect	84	17	85	18
rect	84	18	85	19
rect	84	20	85	21
rect	84	21	85	22
rect	84	23	85	24
rect	84	24	85	25
rect	84	26	85	27
rect	84	27	85	28
rect	84	29	85	30
rect	84	30	85	31
rect	84	32	85	33
rect	84	33	85	34
rect	84	35	85	36
rect	84	36	85	37
rect	84	38	85	39
rect	84	39	85	40
rect	84	41	85	42
rect	84	42	85	43
rect	84	44	85	45
rect	84	45	85	46
rect	84	47	85	48
rect	84	48	85	49
rect	84	50	85	51
rect	84	51	85	52
rect	84	53	85	54
rect	84	54	85	55
rect	84	56	85	57
rect	84	57	85	58
rect	84	59	85	60
rect	84	60	85	61
rect	84	62	85	63
rect	84	63	85	64
rect	84	65	85	66
rect	84	66	85	67
rect	84	68	85	69
rect	84	69	85	70
rect	84	71	85	72
rect	84	72	85	73
rect	84	74	85	75
rect	84	75	85	76
rect	84	77	85	78
rect	84	78	85	79
rect	84	80	85	81
rect	84	81	85	82
rect	84	83	85	84
rect	84	84	85	85
rect	84	86	85	87
rect	84	87	85	88
rect	84	89	85	90
rect	84	90	85	91
rect	84	92	85	93
rect	84	93	85	94
rect	84	95	85	96
rect	84	96	85	97
rect	84	98	85	99
rect	84	99	85	100
rect	84	101	85	102
rect	84	102	85	103
rect	84	104	85	105
rect	84	105	85	106
rect	84	107	85	108
rect	84	108	85	109
rect	84	110	85	111
rect	84	111	85	112
rect	84	113	85	114
rect	84	114	85	115
rect	84	116	85	117
rect	84	117	85	118
rect	84	119	85	120
rect	84	120	85	121
rect	84	122	85	123
rect	84	123	85	124
rect	84	125	85	126
rect	84	126	85	127
rect	84	128	85	129
rect	84	129	85	130
rect	84	131	85	132
rect	84	132	85	133
rect	84	134	85	135
rect	84	135	85	136
rect	84	137	85	138
rect	84	138	85	139
rect	84	140	85	141
rect	84	141	85	142
rect	84	143	85	144
rect	84	144	85	145
rect	84	146	85	147
rect	84	147	85	148
rect	84	149	85	150
rect	84	150	85	151
rect	84	152	85	153
rect	84	153	85	154
rect	84	155	85	156
rect	84	156	85	157
rect	84	158	85	159
rect	84	159	85	160
rect	84	161	85	162
rect	84	162	85	163
rect	84	164	85	165
rect	84	165	85	166
rect	84	167	85	168
rect	84	168	85	169
rect	84	170	85	171
rect	84	171	85	172
rect	84	173	85	174
rect	84	174	85	175
rect	84	176	85	177
rect	84	177	85	178
rect	84	179	85	180
rect	84	180	85	181
rect	84	182	85	183
rect	84	183	85	184
rect	84	185	85	186
rect	84	186	85	187
rect	84	188	85	189
rect	84	189	85	190
rect	84	191	85	192
rect	84	192	85	193
rect	84	194	85	195
rect	84	195	85	196
rect	84	197	85	198
rect	84	198	85	199
rect	84	200	85	201
rect	84	201	85	202
rect	84	203	85	204
rect	84	204	85	205
rect	84	206	85	207
rect	84	207	85	208
rect	84	209	85	210
rect	84	210	85	211
rect	84	212	85	213
rect	84	213	85	214
rect	84	215	85	216
rect	84	216	85	217
rect	84	218	85	219
rect	84	219	85	220
rect	84	221	85	222
rect	84	222	85	223
rect	84	224	85	225
rect	84	225	85	226
rect	84	227	85	228
rect	84	228	85	229
rect	84	230	85	231
rect	84	231	85	232
rect	84	233	85	234
rect	84	234	85	235
rect	84	236	85	237
rect	84	237	85	238
rect	84	239	85	240
rect	84	240	85	241
rect	84	242	85	243
rect	84	243	85	244
rect	84	245	85	246
rect	84	246	85	247
rect	84	248	85	249
rect	84	249	85	250
rect	84	251	85	252
rect	84	252	85	253
rect	84	254	85	255
rect	84	255	85	256
rect	84	257	85	258
rect	84	258	85	259
rect	84	260	85	261
rect	84	261	85	262
rect	84	263	85	264
rect	84	264	85	265
rect	84	266	85	267
rect	84	267	85	268
rect	84	269	85	270
rect	84	270	85	271
rect	84	272	85	273
rect	84	273	85	274
rect	84	275	85	276
rect	84	276	85	277
rect	84	278	85	279
rect	84	279	85	280
rect	84	281	85	282
rect	84	282	85	283
rect	84	284	85	285
rect	84	285	85	286
rect	84	287	85	288
rect	84	288	85	289
rect	84	290	85	291
rect	84	291	85	292
rect	84	293	85	294
rect	84	294	85	295
rect	84	296	85	297
rect	84	297	85	298
rect	84	299	85	300
rect	84	300	85	301
rect	84	302	85	303
rect	84	303	85	304
rect	84	305	85	306
rect	84	306	85	307
rect	84	308	85	309
rect	84	309	85	310
rect	84	311	85	312
rect	84	312	85	313
rect	84	314	85	315
rect	84	315	85	316
rect	84	317	85	318
rect	84	318	85	319
rect	84	320	85	321
rect	84	321	85	322
rect	84	323	85	324
rect	84	324	85	325
rect	84	326	85	327
rect	84	327	85	328
rect	84	329	85	330
rect	85	0	86	1
rect	85	2	86	3
rect	85	3	86	4
rect	85	5	86	6
rect	85	6	86	7
rect	85	8	86	9
rect	85	9	86	10
rect	85	11	86	12
rect	85	12	86	13
rect	85	14	86	15
rect	85	15	86	16
rect	85	17	86	18
rect	85	18	86	19
rect	85	20	86	21
rect	85	21	86	22
rect	85	23	86	24
rect	85	24	86	25
rect	85	26	86	27
rect	85	27	86	28
rect	85	29	86	30
rect	85	30	86	31
rect	85	32	86	33
rect	85	33	86	34
rect	85	35	86	36
rect	85	36	86	37
rect	85	38	86	39
rect	85	39	86	40
rect	85	41	86	42
rect	85	42	86	43
rect	85	44	86	45
rect	85	45	86	46
rect	85	47	86	48
rect	85	48	86	49
rect	85	50	86	51
rect	85	51	86	52
rect	85	53	86	54
rect	85	54	86	55
rect	85	56	86	57
rect	85	57	86	58
rect	85	59	86	60
rect	85	60	86	61
rect	85	62	86	63
rect	85	63	86	64
rect	85	65	86	66
rect	85	66	86	67
rect	85	68	86	69
rect	85	69	86	70
rect	85	71	86	72
rect	85	72	86	73
rect	85	74	86	75
rect	85	75	86	76
rect	85	77	86	78
rect	85	78	86	79
rect	85	80	86	81
rect	85	81	86	82
rect	85	83	86	84
rect	85	84	86	85
rect	85	86	86	87
rect	85	87	86	88
rect	85	89	86	90
rect	85	90	86	91
rect	85	92	86	93
rect	85	93	86	94
rect	85	95	86	96
rect	85	96	86	97
rect	85	98	86	99
rect	85	99	86	100
rect	85	101	86	102
rect	85	102	86	103
rect	85	104	86	105
rect	85	105	86	106
rect	85	107	86	108
rect	85	108	86	109
rect	85	110	86	111
rect	85	111	86	112
rect	85	113	86	114
rect	85	114	86	115
rect	85	116	86	117
rect	85	117	86	118
rect	85	119	86	120
rect	85	120	86	121
rect	85	122	86	123
rect	85	123	86	124
rect	85	125	86	126
rect	85	126	86	127
rect	85	128	86	129
rect	85	129	86	130
rect	85	131	86	132
rect	85	132	86	133
rect	85	134	86	135
rect	85	135	86	136
rect	85	137	86	138
rect	85	138	86	139
rect	85	140	86	141
rect	85	141	86	142
rect	85	143	86	144
rect	85	144	86	145
rect	85	146	86	147
rect	85	147	86	148
rect	85	149	86	150
rect	85	150	86	151
rect	85	152	86	153
rect	85	153	86	154
rect	85	155	86	156
rect	85	156	86	157
rect	85	158	86	159
rect	85	159	86	160
rect	85	161	86	162
rect	85	162	86	163
rect	85	164	86	165
rect	85	165	86	166
rect	85	167	86	168
rect	85	168	86	169
rect	85	170	86	171
rect	85	171	86	172
rect	85	173	86	174
rect	85	174	86	175
rect	85	176	86	177
rect	85	177	86	178
rect	85	179	86	180
rect	85	180	86	181
rect	85	182	86	183
rect	85	183	86	184
rect	85	185	86	186
rect	85	186	86	187
rect	85	188	86	189
rect	85	189	86	190
rect	85	191	86	192
rect	85	192	86	193
rect	85	194	86	195
rect	85	195	86	196
rect	85	197	86	198
rect	85	198	86	199
rect	85	200	86	201
rect	85	201	86	202
rect	85	203	86	204
rect	85	204	86	205
rect	85	206	86	207
rect	85	207	86	208
rect	85	209	86	210
rect	85	210	86	211
rect	85	212	86	213
rect	85	213	86	214
rect	85	215	86	216
rect	85	216	86	217
rect	85	218	86	219
rect	85	219	86	220
rect	85	221	86	222
rect	85	222	86	223
rect	85	224	86	225
rect	85	225	86	226
rect	85	227	86	228
rect	85	228	86	229
rect	85	230	86	231
rect	85	231	86	232
rect	85	233	86	234
rect	85	234	86	235
rect	85	236	86	237
rect	85	237	86	238
rect	85	239	86	240
rect	85	240	86	241
rect	85	242	86	243
rect	85	243	86	244
rect	85	245	86	246
rect	85	246	86	247
rect	85	248	86	249
rect	85	249	86	250
rect	85	251	86	252
rect	85	252	86	253
rect	85	254	86	255
rect	85	255	86	256
rect	85	257	86	258
rect	85	258	86	259
rect	85	260	86	261
rect	85	261	86	262
rect	85	263	86	264
rect	85	264	86	265
rect	85	266	86	267
rect	85	267	86	268
rect	85	269	86	270
rect	85	270	86	271
rect	85	272	86	273
rect	85	273	86	274
rect	85	275	86	276
rect	85	276	86	277
rect	85	278	86	279
rect	85	279	86	280
rect	85	281	86	282
rect	85	282	86	283
rect	85	284	86	285
rect	85	285	86	286
rect	85	287	86	288
rect	85	288	86	289
rect	85	290	86	291
rect	85	291	86	292
rect	85	293	86	294
rect	85	294	86	295
rect	85	296	86	297
rect	85	297	86	298
rect	85	299	86	300
rect	85	300	86	301
rect	85	302	86	303
rect	85	303	86	304
rect	85	305	86	306
rect	85	306	86	307
rect	85	308	86	309
rect	85	309	86	310
rect	85	311	86	312
rect	85	312	86	313
rect	85	314	86	315
rect	85	315	86	316
rect	85	317	86	318
rect	85	318	86	319
rect	85	320	86	321
rect	85	321	86	322
rect	85	323	86	324
rect	85	324	86	325
rect	85	326	86	327
rect	85	327	86	328
rect	85	329	86	330
rect	86	0	87	1
rect	86	2	87	3
rect	86	3	87	4
rect	86	5	87	6
rect	86	6	87	7
rect	86	8	87	9
rect	86	9	87	10
rect	86	11	87	12
rect	86	12	87	13
rect	86	14	87	15
rect	86	15	87	16
rect	86	17	87	18
rect	86	18	87	19
rect	86	20	87	21
rect	86	21	87	22
rect	86	23	87	24
rect	86	24	87	25
rect	86	26	87	27
rect	86	27	87	28
rect	86	29	87	30
rect	86	30	87	31
rect	86	32	87	33
rect	86	33	87	34
rect	86	35	87	36
rect	86	36	87	37
rect	86	38	87	39
rect	86	39	87	40
rect	86	41	87	42
rect	86	42	87	43
rect	86	44	87	45
rect	86	45	87	46
rect	86	47	87	48
rect	86	48	87	49
rect	86	50	87	51
rect	86	51	87	52
rect	86	53	87	54
rect	86	54	87	55
rect	86	56	87	57
rect	86	57	87	58
rect	86	59	87	60
rect	86	60	87	61
rect	86	62	87	63
rect	86	63	87	64
rect	86	65	87	66
rect	86	66	87	67
rect	86	68	87	69
rect	86	69	87	70
rect	86	71	87	72
rect	86	72	87	73
rect	86	74	87	75
rect	86	75	87	76
rect	86	77	87	78
rect	86	78	87	79
rect	86	80	87	81
rect	86	81	87	82
rect	86	83	87	84
rect	86	84	87	85
rect	86	86	87	87
rect	86	87	87	88
rect	86	89	87	90
rect	86	90	87	91
rect	86	92	87	93
rect	86	93	87	94
rect	86	95	87	96
rect	86	96	87	97
rect	86	98	87	99
rect	86	99	87	100
rect	86	101	87	102
rect	86	102	87	103
rect	86	104	87	105
rect	86	105	87	106
rect	86	107	87	108
rect	86	108	87	109
rect	86	110	87	111
rect	86	111	87	112
rect	86	113	87	114
rect	86	114	87	115
rect	86	116	87	117
rect	86	117	87	118
rect	86	119	87	120
rect	86	120	87	121
rect	86	122	87	123
rect	86	123	87	124
rect	86	125	87	126
rect	86	126	87	127
rect	86	128	87	129
rect	86	129	87	130
rect	86	131	87	132
rect	86	132	87	133
rect	86	134	87	135
rect	86	135	87	136
rect	86	137	87	138
rect	86	138	87	139
rect	86	140	87	141
rect	86	141	87	142
rect	86	143	87	144
rect	86	144	87	145
rect	86	146	87	147
rect	86	147	87	148
rect	86	149	87	150
rect	86	150	87	151
rect	86	152	87	153
rect	86	153	87	154
rect	86	155	87	156
rect	86	156	87	157
rect	86	158	87	159
rect	86	159	87	160
rect	86	161	87	162
rect	86	162	87	163
rect	86	164	87	165
rect	86	165	87	166
rect	86	167	87	168
rect	86	168	87	169
rect	86	170	87	171
rect	86	171	87	172
rect	86	173	87	174
rect	86	174	87	175
rect	86	176	87	177
rect	86	177	87	178
rect	86	179	87	180
rect	86	180	87	181
rect	86	182	87	183
rect	86	183	87	184
rect	86	185	87	186
rect	86	186	87	187
rect	86	188	87	189
rect	86	189	87	190
rect	86	191	87	192
rect	86	192	87	193
rect	86	194	87	195
rect	86	195	87	196
rect	86	197	87	198
rect	86	198	87	199
rect	86	200	87	201
rect	86	201	87	202
rect	86	203	87	204
rect	86	204	87	205
rect	86	206	87	207
rect	86	207	87	208
rect	86	209	87	210
rect	86	210	87	211
rect	86	212	87	213
rect	86	213	87	214
rect	86	215	87	216
rect	86	216	87	217
rect	86	218	87	219
rect	86	219	87	220
rect	86	221	87	222
rect	86	222	87	223
rect	86	224	87	225
rect	86	225	87	226
rect	86	227	87	228
rect	86	228	87	229
rect	86	230	87	231
rect	86	231	87	232
rect	86	233	87	234
rect	86	234	87	235
rect	86	236	87	237
rect	86	237	87	238
rect	86	239	87	240
rect	86	240	87	241
rect	86	242	87	243
rect	86	243	87	244
rect	86	245	87	246
rect	86	246	87	247
rect	86	248	87	249
rect	86	249	87	250
rect	86	251	87	252
rect	86	252	87	253
rect	86	254	87	255
rect	86	255	87	256
rect	86	257	87	258
rect	86	258	87	259
rect	86	260	87	261
rect	86	261	87	262
rect	86	263	87	264
rect	86	264	87	265
rect	86	266	87	267
rect	86	267	87	268
rect	86	269	87	270
rect	86	270	87	271
rect	86	272	87	273
rect	86	273	87	274
rect	86	275	87	276
rect	86	276	87	277
rect	86	278	87	279
rect	86	279	87	280
rect	86	281	87	282
rect	86	282	87	283
rect	86	284	87	285
rect	86	285	87	286
rect	86	287	87	288
rect	86	288	87	289
rect	86	290	87	291
rect	86	291	87	292
rect	86	293	87	294
rect	86	294	87	295
rect	86	296	87	297
rect	86	297	87	298
rect	86	299	87	300
rect	86	300	87	301
rect	86	302	87	303
rect	86	303	87	304
rect	86	305	87	306
rect	86	306	87	307
rect	86	308	87	309
rect	86	309	87	310
rect	86	311	87	312
rect	86	312	87	313
rect	86	314	87	315
rect	86	315	87	316
rect	86	317	87	318
rect	86	318	87	319
rect	86	320	87	321
rect	86	321	87	322
rect	86	323	87	324
rect	86	324	87	325
rect	86	326	87	327
rect	86	327	87	328
rect	86	329	87	330
rect	93	0	94	1
rect	93	2	94	3
rect	93	3	94	4
rect	93	5	94	6
rect	93	6	94	7
rect	93	8	94	9
rect	93	9	94	10
rect	93	11	94	12
rect	93	12	94	13
rect	93	14	94	15
rect	93	15	94	16
rect	93	17	94	18
rect	93	18	94	19
rect	93	20	94	21
rect	93	21	94	22
rect	93	23	94	24
rect	93	24	94	25
rect	93	26	94	27
rect	93	27	94	28
rect	93	29	94	30
rect	93	30	94	31
rect	93	32	94	33
rect	93	33	94	34
rect	93	35	94	36
rect	93	36	94	37
rect	93	38	94	39
rect	93	39	94	40
rect	93	41	94	42
rect	93	42	94	43
rect	93	44	94	45
rect	93	45	94	46
rect	93	47	94	48
rect	93	48	94	49
rect	93	50	94	51
rect	93	51	94	52
rect	93	53	94	54
rect	93	54	94	55
rect	93	56	94	57
rect	93	57	94	58
rect	93	59	94	60
rect	93	60	94	61
rect	93	62	94	63
rect	93	63	94	64
rect	93	65	94	66
rect	93	66	94	67
rect	93	68	94	69
rect	93	69	94	70
rect	93	71	94	72
rect	93	72	94	73
rect	93	74	94	75
rect	93	75	94	76
rect	93	77	94	78
rect	93	78	94	79
rect	93	80	94	81
rect	93	81	94	82
rect	93	83	94	84
rect	93	84	94	85
rect	93	86	94	87
rect	93	87	94	88
rect	93	89	94	90
rect	93	90	94	91
rect	93	92	94	93
rect	93	93	94	94
rect	93	95	94	96
rect	93	96	94	97
rect	93	98	94	99
rect	93	99	94	100
rect	93	101	94	102
rect	93	102	94	103
rect	93	104	94	105
rect	93	105	94	106
rect	93	107	94	108
rect	93	108	94	109
rect	93	110	94	111
rect	93	111	94	112
rect	93	113	94	114
rect	93	114	94	115
rect	93	116	94	117
rect	93	117	94	118
rect	93	119	94	120
rect	93	120	94	121
rect	93	122	94	123
rect	93	123	94	124
rect	93	125	94	126
rect	93	126	94	127
rect	93	128	94	129
rect	93	129	94	130
rect	93	131	94	132
rect	93	132	94	133
rect	93	134	94	135
rect	93	135	94	136
rect	93	137	94	138
rect	93	138	94	139
rect	93	140	94	141
rect	93	141	94	142
rect	93	143	94	144
rect	93	144	94	145
rect	93	146	94	147
rect	93	147	94	148
rect	93	149	94	150
rect	93	150	94	151
rect	93	152	94	153
rect	93	153	94	154
rect	93	155	94	156
rect	93	156	94	157
rect	93	158	94	159
rect	93	159	94	160
rect	93	161	94	162
rect	93	162	94	163
rect	93	164	94	165
rect	93	165	94	166
rect	93	167	94	168
rect	93	168	94	169
rect	93	170	94	171
rect	93	171	94	172
rect	93	173	94	174
rect	93	174	94	175
rect	93	176	94	177
rect	93	177	94	178
rect	93	179	94	180
rect	93	180	94	181
rect	93	182	94	183
rect	93	183	94	184
rect	93	185	94	186
rect	93	186	94	187
rect	93	188	94	189
rect	93	189	94	190
rect	93	191	94	192
rect	93	192	94	193
rect	93	194	94	195
rect	93	195	94	196
rect	93	197	94	198
rect	93	198	94	199
rect	93	200	94	201
rect	93	201	94	202
rect	93	203	94	204
rect	93	204	94	205
rect	93	206	94	207
rect	93	207	94	208
rect	93	209	94	210
rect	93	210	94	211
rect	93	212	94	213
rect	93	213	94	214
rect	93	215	94	216
rect	93	216	94	217
rect	93	218	94	219
rect	93	219	94	220
rect	93	221	94	222
rect	93	222	94	223
rect	93	224	94	225
rect	93	225	94	226
rect	93	227	94	228
rect	93	228	94	229
rect	93	230	94	231
rect	93	231	94	232
rect	93	233	94	234
rect	93	234	94	235
rect	93	236	94	237
rect	93	237	94	238
rect	93	239	94	240
rect	93	240	94	241
rect	93	242	94	243
rect	93	243	94	244
rect	93	245	94	246
rect	93	246	94	247
rect	93	248	94	249
rect	93	249	94	250
rect	93	251	94	252
rect	93	252	94	253
rect	93	254	94	255
rect	93	255	94	256
rect	93	257	94	258
rect	93	258	94	259
rect	93	260	94	261
rect	93	261	94	262
rect	93	263	94	264
rect	93	264	94	265
rect	93	266	94	267
rect	93	267	94	268
rect	93	269	94	270
rect	93	270	94	271
rect	93	272	94	273
rect	93	273	94	274
rect	93	275	94	276
rect	93	276	94	277
rect	93	278	94	279
rect	93	279	94	280
rect	93	281	94	282
rect	93	282	94	283
rect	93	284	94	285
rect	93	285	94	286
rect	93	287	94	288
rect	93	288	94	289
rect	93	290	94	291
rect	93	291	94	292
rect	93	293	94	294
rect	93	294	94	295
rect	93	296	94	297
rect	93	297	94	298
rect	93	299	94	300
rect	93	300	94	301
rect	93	302	94	303
rect	93	303	94	304
rect	93	305	94	306
rect	93	306	94	307
rect	93	308	94	309
rect	93	309	94	310
rect	93	311	94	312
rect	93	312	94	313
rect	93	314	94	315
rect	93	315	94	316
rect	93	317	94	318
rect	93	318	94	319
rect	93	320	94	321
rect	93	321	94	322
rect	93	323	94	324
rect	93	324	94	325
rect	93	326	94	327
rect	93	327	94	328
rect	93	329	94	330
rect	95	0	96	1
rect	95	2	96	3
rect	95	3	96	4
rect	95	5	96	6
rect	95	6	96	7
rect	95	8	96	9
rect	95	9	96	10
rect	95	11	96	12
rect	95	12	96	13
rect	95	14	96	15
rect	95	15	96	16
rect	95	17	96	18
rect	95	18	96	19
rect	95	20	96	21
rect	95	21	96	22
rect	95	23	96	24
rect	95	24	96	25
rect	95	26	96	27
rect	95	27	96	28
rect	95	29	96	30
rect	95	30	96	31
rect	95	32	96	33
rect	95	33	96	34
rect	95	35	96	36
rect	95	36	96	37
rect	95	38	96	39
rect	95	39	96	40
rect	95	41	96	42
rect	95	42	96	43
rect	95	44	96	45
rect	95	45	96	46
rect	95	47	96	48
rect	95	48	96	49
rect	95	50	96	51
rect	95	51	96	52
rect	95	53	96	54
rect	95	54	96	55
rect	95	56	96	57
rect	95	57	96	58
rect	95	59	96	60
rect	95	60	96	61
rect	95	62	96	63
rect	95	63	96	64
rect	95	65	96	66
rect	95	66	96	67
rect	95	68	96	69
rect	95	69	96	70
rect	95	71	96	72
rect	95	72	96	73
rect	95	74	96	75
rect	95	75	96	76
rect	95	77	96	78
rect	95	78	96	79
rect	95	80	96	81
rect	95	81	96	82
rect	95	83	96	84
rect	95	84	96	85
rect	95	86	96	87
rect	95	87	96	88
rect	95	89	96	90
rect	95	90	96	91
rect	95	92	96	93
rect	95	93	96	94
rect	95	95	96	96
rect	95	96	96	97
rect	95	98	96	99
rect	95	99	96	100
rect	95	101	96	102
rect	95	102	96	103
rect	95	104	96	105
rect	95	105	96	106
rect	95	107	96	108
rect	95	108	96	109
rect	95	110	96	111
rect	95	111	96	112
rect	95	113	96	114
rect	95	114	96	115
rect	95	116	96	117
rect	95	117	96	118
rect	95	119	96	120
rect	95	120	96	121
rect	95	122	96	123
rect	95	123	96	124
rect	95	125	96	126
rect	95	126	96	127
rect	95	128	96	129
rect	95	129	96	130
rect	95	131	96	132
rect	95	132	96	133
rect	95	134	96	135
rect	95	135	96	136
rect	95	137	96	138
rect	95	138	96	139
rect	95	140	96	141
rect	95	141	96	142
rect	95	143	96	144
rect	95	144	96	145
rect	95	146	96	147
rect	95	147	96	148
rect	95	149	96	150
rect	95	150	96	151
rect	95	152	96	153
rect	95	153	96	154
rect	95	155	96	156
rect	95	156	96	157
rect	95	158	96	159
rect	95	159	96	160
rect	95	161	96	162
rect	95	162	96	163
rect	95	164	96	165
rect	95	165	96	166
rect	95	167	96	168
rect	95	168	96	169
rect	95	170	96	171
rect	95	171	96	172
rect	95	173	96	174
rect	95	174	96	175
rect	95	176	96	177
rect	95	177	96	178
rect	95	179	96	180
rect	95	180	96	181
rect	95	182	96	183
rect	95	183	96	184
rect	95	185	96	186
rect	95	186	96	187
rect	95	188	96	189
rect	95	189	96	190
rect	95	191	96	192
rect	95	192	96	193
rect	95	194	96	195
rect	95	195	96	196
rect	95	197	96	198
rect	95	198	96	199
rect	95	200	96	201
rect	95	201	96	202
rect	95	203	96	204
rect	95	204	96	205
rect	95	206	96	207
rect	95	207	96	208
rect	95	209	96	210
rect	95	210	96	211
rect	95	212	96	213
rect	95	213	96	214
rect	95	215	96	216
rect	95	216	96	217
rect	95	218	96	219
rect	95	219	96	220
rect	95	221	96	222
rect	95	222	96	223
rect	95	224	96	225
rect	95	225	96	226
rect	95	227	96	228
rect	95	228	96	229
rect	95	230	96	231
rect	95	231	96	232
rect	95	233	96	234
rect	95	234	96	235
rect	95	236	96	237
rect	95	237	96	238
rect	95	239	96	240
rect	95	240	96	241
rect	95	242	96	243
rect	95	243	96	244
rect	95	245	96	246
rect	95	246	96	247
rect	95	248	96	249
rect	95	249	96	250
rect	95	251	96	252
rect	95	252	96	253
rect	95	254	96	255
rect	95	255	96	256
rect	95	257	96	258
rect	95	258	96	259
rect	95	260	96	261
rect	95	261	96	262
rect	95	263	96	264
rect	95	264	96	265
rect	95	266	96	267
rect	95	267	96	268
rect	95	269	96	270
rect	95	270	96	271
rect	95	272	96	273
rect	95	273	96	274
rect	95	275	96	276
rect	95	276	96	277
rect	95	278	96	279
rect	95	279	96	280
rect	95	281	96	282
rect	95	282	96	283
rect	95	284	96	285
rect	95	285	96	286
rect	95	287	96	288
rect	95	288	96	289
rect	95	290	96	291
rect	95	291	96	292
rect	95	293	96	294
rect	95	294	96	295
rect	95	296	96	297
rect	95	297	96	298
rect	95	299	96	300
rect	95	300	96	301
rect	95	302	96	303
rect	95	303	96	304
rect	95	305	96	306
rect	95	306	96	307
rect	95	308	96	309
rect	95	309	96	310
rect	95	311	96	312
rect	95	312	96	313
rect	95	314	96	315
rect	95	315	96	316
rect	95	317	96	318
rect	95	318	96	319
rect	95	320	96	321
rect	95	321	96	322
rect	95	323	96	324
rect	95	324	96	325
rect	95	326	96	327
rect	95	327	96	328
rect	95	329	96	330
rect	95	330	96	331
rect	95	332	96	333
rect	95	333	96	334
rect	95	335	96	336
rect	96	0	97	1
rect	96	2	97	3
rect	96	3	97	4
rect	96	5	97	6
rect	96	6	97	7
rect	96	8	97	9
rect	96	9	97	10
rect	96	11	97	12
rect	96	12	97	13
rect	96	14	97	15
rect	96	15	97	16
rect	96	17	97	18
rect	96	18	97	19
rect	96	20	97	21
rect	96	21	97	22
rect	96	23	97	24
rect	96	24	97	25
rect	96	26	97	27
rect	96	27	97	28
rect	96	29	97	30
rect	96	30	97	31
rect	96	32	97	33
rect	96	33	97	34
rect	96	35	97	36
rect	96	36	97	37
rect	96	38	97	39
rect	96	39	97	40
rect	96	41	97	42
rect	96	42	97	43
rect	96	44	97	45
rect	96	45	97	46
rect	96	47	97	48
rect	96	48	97	49
rect	96	50	97	51
rect	96	51	97	52
rect	96	53	97	54
rect	96	54	97	55
rect	96	56	97	57
rect	96	57	97	58
rect	96	59	97	60
rect	96	60	97	61
rect	96	62	97	63
rect	96	63	97	64
rect	96	65	97	66
rect	96	66	97	67
rect	96	68	97	69
rect	96	69	97	70
rect	96	71	97	72
rect	96	72	97	73
rect	96	74	97	75
rect	96	75	97	76
rect	96	77	97	78
rect	96	78	97	79
rect	96	80	97	81
rect	96	81	97	82
rect	96	83	97	84
rect	96	84	97	85
rect	96	86	97	87
rect	96	87	97	88
rect	96	89	97	90
rect	96	90	97	91
rect	96	92	97	93
rect	96	93	97	94
rect	96	95	97	96
rect	96	96	97	97
rect	96	98	97	99
rect	96	99	97	100
rect	96	101	97	102
rect	96	102	97	103
rect	96	104	97	105
rect	96	105	97	106
rect	96	107	97	108
rect	96	108	97	109
rect	96	110	97	111
rect	96	111	97	112
rect	96	113	97	114
rect	96	114	97	115
rect	96	116	97	117
rect	96	117	97	118
rect	96	119	97	120
rect	96	120	97	121
rect	96	122	97	123
rect	96	123	97	124
rect	96	125	97	126
rect	96	126	97	127
rect	96	128	97	129
rect	96	129	97	130
rect	96	131	97	132
rect	96	132	97	133
rect	96	134	97	135
rect	96	135	97	136
rect	96	137	97	138
rect	96	138	97	139
rect	96	140	97	141
rect	96	141	97	142
rect	96	143	97	144
rect	96	144	97	145
rect	96	146	97	147
rect	96	147	97	148
rect	96	149	97	150
rect	96	150	97	151
rect	96	152	97	153
rect	96	153	97	154
rect	96	155	97	156
rect	96	156	97	157
rect	96	158	97	159
rect	96	159	97	160
rect	96	161	97	162
rect	96	162	97	163
rect	96	164	97	165
rect	96	165	97	166
rect	96	167	97	168
rect	96	168	97	169
rect	96	170	97	171
rect	96	171	97	172
rect	96	173	97	174
rect	96	174	97	175
rect	96	176	97	177
rect	96	177	97	178
rect	96	179	97	180
rect	96	180	97	181
rect	96	182	97	183
rect	96	183	97	184
rect	96	185	97	186
rect	96	186	97	187
rect	96	188	97	189
rect	96	189	97	190
rect	96	191	97	192
rect	96	192	97	193
rect	96	194	97	195
rect	96	195	97	196
rect	96	197	97	198
rect	96	198	97	199
rect	96	200	97	201
rect	96	201	97	202
rect	96	203	97	204
rect	96	204	97	205
rect	96	206	97	207
rect	96	207	97	208
rect	96	209	97	210
rect	96	210	97	211
rect	96	212	97	213
rect	96	213	97	214
rect	96	215	97	216
rect	96	216	97	217
rect	96	218	97	219
rect	96	219	97	220
rect	96	221	97	222
rect	96	222	97	223
rect	96	224	97	225
rect	96	225	97	226
rect	96	227	97	228
rect	96	228	97	229
rect	96	230	97	231
rect	96	231	97	232
rect	96	233	97	234
rect	96	234	97	235
rect	96	236	97	237
rect	96	237	97	238
rect	96	239	97	240
rect	96	240	97	241
rect	96	242	97	243
rect	96	243	97	244
rect	96	245	97	246
rect	96	246	97	247
rect	96	248	97	249
rect	96	249	97	250
rect	96	251	97	252
rect	96	252	97	253
rect	96	254	97	255
rect	96	255	97	256
rect	96	257	97	258
rect	96	258	97	259
rect	96	260	97	261
rect	96	261	97	262
rect	96	263	97	264
rect	96	264	97	265
rect	96	266	97	267
rect	96	267	97	268
rect	96	269	97	270
rect	96	270	97	271
rect	96	272	97	273
rect	96	273	97	274
rect	96	275	97	276
rect	96	276	97	277
rect	96	278	97	279
rect	96	279	97	280
rect	96	281	97	282
rect	96	282	97	283
rect	96	284	97	285
rect	96	285	97	286
rect	96	287	97	288
rect	96	288	97	289
rect	96	290	97	291
rect	96	291	97	292
rect	96	293	97	294
rect	96	294	97	295
rect	96	296	97	297
rect	96	297	97	298
rect	96	299	97	300
rect	96	300	97	301
rect	96	302	97	303
rect	96	303	97	304
rect	96	305	97	306
rect	96	306	97	307
rect	96	308	97	309
rect	96	309	97	310
rect	96	311	97	312
rect	96	312	97	313
rect	96	314	97	315
rect	96	315	97	316
rect	96	317	97	318
rect	96	318	97	319
rect	96	320	97	321
rect	96	321	97	322
rect	96	323	97	324
rect	96	324	97	325
rect	96	326	97	327
rect	96	327	97	328
rect	96	329	97	330
rect	96	330	97	331
rect	96	332	97	333
rect	96	333	97	334
rect	96	335	97	336
rect	97	0	98	1
rect	97	2	98	3
rect	97	3	98	4
rect	97	5	98	6
rect	97	6	98	7
rect	97	8	98	9
rect	97	9	98	10
rect	97	11	98	12
rect	97	12	98	13
rect	97	14	98	15
rect	97	15	98	16
rect	97	17	98	18
rect	97	18	98	19
rect	97	20	98	21
rect	97	21	98	22
rect	97	23	98	24
rect	97	24	98	25
rect	97	26	98	27
rect	97	27	98	28
rect	97	29	98	30
rect	97	30	98	31
rect	97	32	98	33
rect	97	33	98	34
rect	97	35	98	36
rect	97	36	98	37
rect	97	38	98	39
rect	97	39	98	40
rect	97	41	98	42
rect	97	42	98	43
rect	97	44	98	45
rect	97	45	98	46
rect	97	47	98	48
rect	97	48	98	49
rect	97	50	98	51
rect	97	51	98	52
rect	97	53	98	54
rect	97	54	98	55
rect	97	56	98	57
rect	97	57	98	58
rect	97	59	98	60
rect	97	60	98	61
rect	97	62	98	63
rect	97	63	98	64
rect	97	65	98	66
rect	97	66	98	67
rect	97	68	98	69
rect	97	69	98	70
rect	97	71	98	72
rect	97	72	98	73
rect	97	74	98	75
rect	97	75	98	76
rect	97	77	98	78
rect	97	78	98	79
rect	97	80	98	81
rect	97	81	98	82
rect	97	83	98	84
rect	97	84	98	85
rect	97	86	98	87
rect	97	87	98	88
rect	97	89	98	90
rect	97	90	98	91
rect	97	92	98	93
rect	97	93	98	94
rect	97	95	98	96
rect	97	96	98	97
rect	97	98	98	99
rect	97	99	98	100
rect	97	101	98	102
rect	97	102	98	103
rect	97	104	98	105
rect	97	105	98	106
rect	97	107	98	108
rect	97	108	98	109
rect	97	110	98	111
rect	97	111	98	112
rect	97	113	98	114
rect	97	114	98	115
rect	97	116	98	117
rect	97	117	98	118
rect	97	119	98	120
rect	97	120	98	121
rect	97	122	98	123
rect	97	123	98	124
rect	97	125	98	126
rect	97	126	98	127
rect	97	128	98	129
rect	97	129	98	130
rect	97	131	98	132
rect	97	132	98	133
rect	97	134	98	135
rect	97	135	98	136
rect	97	137	98	138
rect	97	138	98	139
rect	97	140	98	141
rect	97	141	98	142
rect	97	143	98	144
rect	97	144	98	145
rect	97	146	98	147
rect	97	147	98	148
rect	97	149	98	150
rect	97	150	98	151
rect	97	152	98	153
rect	97	153	98	154
rect	97	155	98	156
rect	97	156	98	157
rect	97	158	98	159
rect	97	159	98	160
rect	97	161	98	162
rect	97	162	98	163
rect	97	164	98	165
rect	97	165	98	166
rect	97	167	98	168
rect	97	168	98	169
rect	97	170	98	171
rect	97	171	98	172
rect	97	173	98	174
rect	97	174	98	175
rect	97	176	98	177
rect	97	177	98	178
rect	97	179	98	180
rect	97	180	98	181
rect	97	182	98	183
rect	97	183	98	184
rect	97	185	98	186
rect	97	186	98	187
rect	97	188	98	189
rect	97	189	98	190
rect	97	191	98	192
rect	97	192	98	193
rect	97	194	98	195
rect	97	195	98	196
rect	97	197	98	198
rect	97	198	98	199
rect	97	200	98	201
rect	97	201	98	202
rect	97	203	98	204
rect	97	204	98	205
rect	97	206	98	207
rect	97	207	98	208
rect	97	209	98	210
rect	97	210	98	211
rect	97	212	98	213
rect	97	213	98	214
rect	97	215	98	216
rect	97	216	98	217
rect	97	218	98	219
rect	97	219	98	220
rect	97	221	98	222
rect	97	222	98	223
rect	97	224	98	225
rect	97	225	98	226
rect	97	227	98	228
rect	97	228	98	229
rect	97	230	98	231
rect	97	231	98	232
rect	97	233	98	234
rect	97	234	98	235
rect	97	236	98	237
rect	97	237	98	238
rect	97	239	98	240
rect	97	240	98	241
rect	97	242	98	243
rect	97	243	98	244
rect	97	245	98	246
rect	97	246	98	247
rect	97	248	98	249
rect	97	249	98	250
rect	97	251	98	252
rect	97	252	98	253
rect	97	254	98	255
rect	97	255	98	256
rect	97	257	98	258
rect	97	258	98	259
rect	97	260	98	261
rect	97	261	98	262
rect	97	263	98	264
rect	97	264	98	265
rect	97	266	98	267
rect	97	267	98	268
rect	97	269	98	270
rect	97	270	98	271
rect	97	272	98	273
rect	97	273	98	274
rect	97	275	98	276
rect	97	276	98	277
rect	97	278	98	279
rect	97	279	98	280
rect	97	281	98	282
rect	97	282	98	283
rect	97	284	98	285
rect	97	285	98	286
rect	97	287	98	288
rect	97	288	98	289
rect	97	290	98	291
rect	97	291	98	292
rect	97	293	98	294
rect	97	294	98	295
rect	97	296	98	297
rect	97	297	98	298
rect	97	299	98	300
rect	97	300	98	301
rect	97	302	98	303
rect	97	303	98	304
rect	97	305	98	306
rect	97	306	98	307
rect	97	308	98	309
rect	97	309	98	310
rect	97	311	98	312
rect	97	312	98	313
rect	97	314	98	315
rect	97	315	98	316
rect	97	317	98	318
rect	97	318	98	319
rect	97	320	98	321
rect	97	321	98	322
rect	97	323	98	324
rect	97	324	98	325
rect	97	326	98	327
rect	97	327	98	328
rect	97	329	98	330
rect	97	330	98	331
rect	97	332	98	333
rect	97	333	98	334
rect	97	335	98	336
rect	98	0	99	1
rect	98	2	99	3
rect	98	3	99	4
rect	98	5	99	6
rect	98	6	99	7
rect	98	8	99	9
rect	98	9	99	10
rect	98	11	99	12
rect	98	12	99	13
rect	98	14	99	15
rect	98	15	99	16
rect	98	17	99	18
rect	98	18	99	19
rect	98	20	99	21
rect	98	21	99	22
rect	98	23	99	24
rect	98	24	99	25
rect	98	26	99	27
rect	98	27	99	28
rect	98	29	99	30
rect	98	30	99	31
rect	98	32	99	33
rect	98	33	99	34
rect	98	35	99	36
rect	98	36	99	37
rect	98	38	99	39
rect	98	39	99	40
rect	98	41	99	42
rect	98	42	99	43
rect	98	44	99	45
rect	98	45	99	46
rect	98	47	99	48
rect	98	48	99	49
rect	98	50	99	51
rect	98	51	99	52
rect	98	53	99	54
rect	98	54	99	55
rect	98	56	99	57
rect	98	57	99	58
rect	98	59	99	60
rect	98	60	99	61
rect	98	62	99	63
rect	98	63	99	64
rect	98	65	99	66
rect	98	66	99	67
rect	98	68	99	69
rect	98	69	99	70
rect	98	71	99	72
rect	98	72	99	73
rect	98	74	99	75
rect	98	75	99	76
rect	98	77	99	78
rect	98	78	99	79
rect	98	80	99	81
rect	98	81	99	82
rect	98	83	99	84
rect	98	84	99	85
rect	98	86	99	87
rect	98	87	99	88
rect	98	89	99	90
rect	98	90	99	91
rect	98	92	99	93
rect	98	93	99	94
rect	98	95	99	96
rect	98	96	99	97
rect	98	98	99	99
rect	98	99	99	100
rect	98	101	99	102
rect	98	102	99	103
rect	98	104	99	105
rect	98	105	99	106
rect	98	107	99	108
rect	98	108	99	109
rect	98	110	99	111
rect	98	111	99	112
rect	98	113	99	114
rect	98	114	99	115
rect	98	116	99	117
rect	98	117	99	118
rect	98	119	99	120
rect	98	120	99	121
rect	98	122	99	123
rect	98	123	99	124
rect	98	125	99	126
rect	98	126	99	127
rect	98	128	99	129
rect	98	129	99	130
rect	98	131	99	132
rect	98	132	99	133
rect	98	134	99	135
rect	98	135	99	136
rect	98	137	99	138
rect	98	138	99	139
rect	98	140	99	141
rect	98	141	99	142
rect	98	143	99	144
rect	98	144	99	145
rect	98	146	99	147
rect	98	147	99	148
rect	98	149	99	150
rect	98	150	99	151
rect	98	152	99	153
rect	98	153	99	154
rect	98	155	99	156
rect	98	156	99	157
rect	98	158	99	159
rect	98	159	99	160
rect	98	161	99	162
rect	98	162	99	163
rect	98	164	99	165
rect	98	165	99	166
rect	98	167	99	168
rect	98	168	99	169
rect	98	170	99	171
rect	98	171	99	172
rect	98	173	99	174
rect	98	174	99	175
rect	98	176	99	177
rect	98	177	99	178
rect	98	179	99	180
rect	98	180	99	181
rect	98	182	99	183
rect	98	183	99	184
rect	98	185	99	186
rect	98	186	99	187
rect	98	188	99	189
rect	98	189	99	190
rect	98	191	99	192
rect	98	192	99	193
rect	98	194	99	195
rect	98	195	99	196
rect	98	197	99	198
rect	98	198	99	199
rect	98	200	99	201
rect	98	201	99	202
rect	98	203	99	204
rect	98	204	99	205
rect	98	206	99	207
rect	98	207	99	208
rect	98	209	99	210
rect	98	210	99	211
rect	98	212	99	213
rect	98	213	99	214
rect	98	215	99	216
rect	98	216	99	217
rect	98	218	99	219
rect	98	219	99	220
rect	98	221	99	222
rect	98	222	99	223
rect	98	224	99	225
rect	98	225	99	226
rect	98	227	99	228
rect	98	228	99	229
rect	98	230	99	231
rect	98	231	99	232
rect	98	233	99	234
rect	98	234	99	235
rect	98	236	99	237
rect	98	237	99	238
rect	98	239	99	240
rect	98	240	99	241
rect	98	242	99	243
rect	98	243	99	244
rect	98	245	99	246
rect	98	246	99	247
rect	98	248	99	249
rect	98	249	99	250
rect	98	251	99	252
rect	98	252	99	253
rect	98	254	99	255
rect	98	255	99	256
rect	98	257	99	258
rect	98	258	99	259
rect	98	260	99	261
rect	98	261	99	262
rect	98	263	99	264
rect	98	264	99	265
rect	98	266	99	267
rect	98	267	99	268
rect	98	269	99	270
rect	98	270	99	271
rect	98	272	99	273
rect	98	273	99	274
rect	98	275	99	276
rect	98	276	99	277
rect	98	278	99	279
rect	98	279	99	280
rect	98	281	99	282
rect	98	282	99	283
rect	98	284	99	285
rect	98	285	99	286
rect	98	287	99	288
rect	98	288	99	289
rect	98	290	99	291
rect	98	291	99	292
rect	98	293	99	294
rect	98	294	99	295
rect	98	296	99	297
rect	98	297	99	298
rect	98	299	99	300
rect	98	300	99	301
rect	98	302	99	303
rect	98	303	99	304
rect	98	305	99	306
rect	98	306	99	307
rect	98	308	99	309
rect	98	309	99	310
rect	98	311	99	312
rect	98	312	99	313
rect	98	314	99	315
rect	98	315	99	316
rect	98	317	99	318
rect	98	318	99	319
rect	98	320	99	321
rect	98	321	99	322
rect	98	323	99	324
rect	98	324	99	325
rect	98	326	99	327
rect	98	327	99	328
rect	98	329	99	330
rect	98	330	99	331
rect	98	332	99	333
rect	98	333	99	334
rect	98	335	99	336
rect	99	0	100	1
rect	99	2	100	3
rect	99	3	100	4
rect	99	5	100	6
rect	99	6	100	7
rect	99	8	100	9
rect	99	9	100	10
rect	99	11	100	12
rect	99	12	100	13
rect	99	14	100	15
rect	99	15	100	16
rect	99	17	100	18
rect	99	18	100	19
rect	99	20	100	21
rect	99	21	100	22
rect	99	23	100	24
rect	99	24	100	25
rect	99	26	100	27
rect	99	27	100	28
rect	99	29	100	30
rect	99	30	100	31
rect	99	32	100	33
rect	99	33	100	34
rect	99	35	100	36
rect	99	36	100	37
rect	99	38	100	39
rect	99	39	100	40
rect	99	41	100	42
rect	99	42	100	43
rect	99	44	100	45
rect	99	45	100	46
rect	99	47	100	48
rect	99	48	100	49
rect	99	50	100	51
rect	99	51	100	52
rect	99	53	100	54
rect	99	54	100	55
rect	99	56	100	57
rect	99	57	100	58
rect	99	59	100	60
rect	99	60	100	61
rect	99	62	100	63
rect	99	63	100	64
rect	99	65	100	66
rect	99	66	100	67
rect	99	68	100	69
rect	99	69	100	70
rect	99	71	100	72
rect	99	72	100	73
rect	99	74	100	75
rect	99	75	100	76
rect	99	77	100	78
rect	99	78	100	79
rect	99	80	100	81
rect	99	81	100	82
rect	99	83	100	84
rect	99	84	100	85
rect	99	86	100	87
rect	99	87	100	88
rect	99	89	100	90
rect	99	90	100	91
rect	99	92	100	93
rect	99	93	100	94
rect	99	95	100	96
rect	99	96	100	97
rect	99	98	100	99
rect	99	99	100	100
rect	99	101	100	102
rect	99	102	100	103
rect	99	104	100	105
rect	99	105	100	106
rect	99	107	100	108
rect	99	108	100	109
rect	99	110	100	111
rect	99	111	100	112
rect	99	113	100	114
rect	99	114	100	115
rect	99	116	100	117
rect	99	117	100	118
rect	99	119	100	120
rect	99	120	100	121
rect	99	122	100	123
rect	99	123	100	124
rect	99	125	100	126
rect	99	126	100	127
rect	99	128	100	129
rect	99	129	100	130
rect	99	131	100	132
rect	99	132	100	133
rect	99	134	100	135
rect	99	135	100	136
rect	99	137	100	138
rect	99	138	100	139
rect	99	140	100	141
rect	99	141	100	142
rect	99	143	100	144
rect	99	144	100	145
rect	99	146	100	147
rect	99	147	100	148
rect	99	149	100	150
rect	99	150	100	151
rect	99	152	100	153
rect	99	153	100	154
rect	99	155	100	156
rect	99	156	100	157
rect	99	158	100	159
rect	99	159	100	160
rect	99	161	100	162
rect	99	162	100	163
rect	99	164	100	165
rect	99	165	100	166
rect	99	167	100	168
rect	99	168	100	169
rect	99	170	100	171
rect	99	171	100	172
rect	99	173	100	174
rect	99	174	100	175
rect	99	176	100	177
rect	99	177	100	178
rect	99	179	100	180
rect	99	180	100	181
rect	99	182	100	183
rect	99	183	100	184
rect	99	185	100	186
rect	99	186	100	187
rect	99	188	100	189
rect	99	189	100	190
rect	99	191	100	192
rect	99	192	100	193
rect	99	194	100	195
rect	99	195	100	196
rect	99	197	100	198
rect	99	198	100	199
rect	99	200	100	201
rect	99	201	100	202
rect	99	203	100	204
rect	99	204	100	205
rect	99	206	100	207
rect	99	207	100	208
rect	99	209	100	210
rect	99	210	100	211
rect	99	212	100	213
rect	99	213	100	214
rect	99	215	100	216
rect	99	216	100	217
rect	99	218	100	219
rect	99	219	100	220
rect	99	221	100	222
rect	99	222	100	223
rect	99	224	100	225
rect	99	225	100	226
rect	99	227	100	228
rect	99	228	100	229
rect	99	230	100	231
rect	99	231	100	232
rect	99	233	100	234
rect	99	234	100	235
rect	99	236	100	237
rect	99	237	100	238
rect	99	239	100	240
rect	99	240	100	241
rect	99	242	100	243
rect	99	243	100	244
rect	99	245	100	246
rect	99	246	100	247
rect	99	248	100	249
rect	99	249	100	250
rect	99	251	100	252
rect	99	252	100	253
rect	99	254	100	255
rect	99	255	100	256
rect	99	257	100	258
rect	99	258	100	259
rect	99	260	100	261
rect	99	261	100	262
rect	99	263	100	264
rect	99	264	100	265
rect	99	266	100	267
rect	99	267	100	268
rect	99	269	100	270
rect	99	270	100	271
rect	99	272	100	273
rect	99	273	100	274
rect	99	275	100	276
rect	99	276	100	277
rect	99	278	100	279
rect	99	279	100	280
rect	99	281	100	282
rect	99	282	100	283
rect	99	284	100	285
rect	99	285	100	286
rect	99	287	100	288
rect	99	288	100	289
rect	99	290	100	291
rect	99	291	100	292
rect	99	293	100	294
rect	99	294	100	295
rect	99	296	100	297
rect	99	297	100	298
rect	99	299	100	300
rect	99	300	100	301
rect	99	302	100	303
rect	99	303	100	304
rect	99	305	100	306
rect	99	306	100	307
rect	99	308	100	309
rect	99	309	100	310
rect	99	311	100	312
rect	99	312	100	313
rect	99	314	100	315
rect	99	315	100	316
rect	99	317	100	318
rect	99	318	100	319
rect	99	320	100	321
rect	99	321	100	322
rect	99	323	100	324
rect	99	324	100	325
rect	99	326	100	327
rect	99	327	100	328
rect	99	329	100	330
rect	99	330	100	331
rect	99	332	100	333
rect	99	333	100	334
rect	99	335	100	336
rect	108	0	109	1
rect	108	2	109	3
rect	108	3	109	4
rect	108	5	109	6
rect	108	6	109	7
rect	108	8	109	9
rect	108	9	109	10
rect	108	11	109	12
rect	108	12	109	13
rect	108	14	109	15
rect	108	15	109	16
rect	108	17	109	18
rect	108	18	109	19
rect	108	20	109	21
rect	108	21	109	22
rect	108	23	109	24
rect	108	24	109	25
rect	108	26	109	27
rect	108	27	109	28
rect	108	29	109	30
rect	108	30	109	31
rect	108	32	109	33
rect	108	33	109	34
rect	108	35	109	36
rect	108	36	109	37
rect	108	38	109	39
rect	108	39	109	40
rect	108	41	109	42
rect	108	42	109	43
rect	108	44	109	45
rect	108	45	109	46
rect	108	47	109	48
rect	108	48	109	49
rect	108	50	109	51
rect	108	51	109	52
rect	108	53	109	54
rect	108	54	109	55
rect	108	56	109	57
rect	108	57	109	58
rect	108	59	109	60
rect	108	60	109	61
rect	108	62	109	63
rect	108	63	109	64
rect	108	65	109	66
rect	108	66	109	67
rect	108	68	109	69
rect	108	69	109	70
rect	108	71	109	72
rect	108	72	109	73
rect	108	74	109	75
rect	108	75	109	76
rect	108	77	109	78
rect	108	78	109	79
rect	108	80	109	81
rect	108	81	109	82
rect	108	83	109	84
rect	108	84	109	85
rect	108	86	109	87
rect	108	87	109	88
rect	108	89	109	90
rect	108	90	109	91
rect	108	92	109	93
rect	108	93	109	94
rect	108	95	109	96
rect	108	96	109	97
rect	108	98	109	99
rect	108	99	109	100
rect	108	101	109	102
rect	108	102	109	103
rect	108	104	109	105
rect	108	105	109	106
rect	108	107	109	108
rect	108	108	109	109
rect	108	110	109	111
rect	108	111	109	112
rect	108	113	109	114
rect	108	114	109	115
rect	108	116	109	117
rect	108	117	109	118
rect	108	119	109	120
rect	108	120	109	121
rect	108	122	109	123
rect	108	123	109	124
rect	108	125	109	126
rect	108	126	109	127
rect	108	128	109	129
rect	108	129	109	130
rect	108	131	109	132
rect	108	132	109	133
rect	108	134	109	135
rect	108	135	109	136
rect	108	137	109	138
rect	108	138	109	139
rect	108	140	109	141
rect	108	141	109	142
rect	108	143	109	144
rect	108	144	109	145
rect	108	146	109	147
rect	108	147	109	148
rect	108	149	109	150
rect	108	150	109	151
rect	108	152	109	153
rect	108	153	109	154
rect	108	155	109	156
rect	108	156	109	157
rect	108	158	109	159
rect	108	159	109	160
rect	108	161	109	162
rect	108	162	109	163
rect	108	164	109	165
rect	108	165	109	166
rect	108	167	109	168
rect	108	168	109	169
rect	108	170	109	171
rect	108	171	109	172
rect	108	173	109	174
rect	108	174	109	175
rect	108	176	109	177
rect	108	177	109	178
rect	108	179	109	180
rect	108	180	109	181
rect	108	182	109	183
rect	108	183	109	184
rect	108	185	109	186
rect	108	186	109	187
rect	108	188	109	189
rect	108	189	109	190
rect	108	191	109	192
rect	108	192	109	193
rect	108	194	109	195
rect	108	195	109	196
rect	108	197	109	198
rect	108	198	109	199
rect	108	200	109	201
rect	108	201	109	202
rect	108	203	109	204
rect	108	204	109	205
rect	108	206	109	207
rect	108	207	109	208
rect	108	209	109	210
rect	108	210	109	211
rect	108	212	109	213
rect	108	213	109	214
rect	108	215	109	216
rect	108	216	109	217
rect	108	218	109	219
rect	108	219	109	220
rect	108	221	109	222
rect	108	222	109	223
rect	108	224	109	225
rect	108	225	109	226
rect	108	227	109	228
rect	108	228	109	229
rect	108	230	109	231
rect	108	231	109	232
rect	108	233	109	234
rect	108	234	109	235
rect	108	236	109	237
rect	108	237	109	238
rect	108	239	109	240
rect	108	240	109	241
rect	108	242	109	243
rect	108	243	109	244
rect	108	245	109	246
rect	108	246	109	247
rect	108	248	109	249
rect	108	249	109	250
rect	108	251	109	252
rect	108	252	109	253
rect	108	254	109	255
rect	108	255	109	256
rect	108	257	109	258
rect	108	258	109	259
rect	108	260	109	261
rect	108	261	109	262
rect	108	263	109	264
rect	108	264	109	265
rect	108	266	109	267
rect	108	267	109	268
rect	108	269	109	270
rect	108	270	109	271
rect	108	272	109	273
rect	108	273	109	274
rect	108	275	109	276
rect	108	276	109	277
rect	108	278	109	279
rect	108	279	109	280
rect	108	281	109	282
rect	108	282	109	283
rect	108	284	109	285
rect	108	285	109	286
rect	108	287	109	288
rect	108	288	109	289
rect	108	290	109	291
rect	108	291	109	292
rect	108	293	109	294
rect	108	294	109	295
rect	108	296	109	297
rect	108	297	109	298
rect	108	299	109	300
rect	108	300	109	301
rect	108	302	109	303
rect	108	303	109	304
rect	108	305	109	306
rect	108	306	109	307
rect	108	308	109	309
rect	108	309	109	310
rect	108	311	109	312
rect	108	312	109	313
rect	108	314	109	315
rect	108	315	109	316
rect	108	317	109	318
rect	108	318	109	319
rect	108	320	109	321
rect	108	321	109	322
rect	108	323	109	324
rect	108	324	109	325
rect	108	326	109	327
rect	108	327	109	328
rect	108	329	109	330
rect	108	330	109	331
rect	108	332	109	333
rect	108	333	109	334
rect	108	335	109	336
rect	110	0	111	1
rect	110	2	111	3
rect	110	3	111	4
rect	110	5	111	6
rect	110	6	111	7
rect	110	8	111	9
rect	110	9	111	10
rect	110	11	111	12
rect	110	12	111	13
rect	110	14	111	15
rect	110	15	111	16
rect	110	17	111	18
rect	110	18	111	19
rect	110	20	111	21
rect	110	21	111	22
rect	110	23	111	24
rect	110	24	111	25
rect	110	26	111	27
rect	110	27	111	28
rect	110	29	111	30
rect	110	30	111	31
rect	110	32	111	33
rect	110	33	111	34
rect	110	35	111	36
rect	110	36	111	37
rect	110	38	111	39
rect	110	39	111	40
rect	110	41	111	42
rect	110	42	111	43
rect	110	44	111	45
rect	110	45	111	46
rect	110	47	111	48
rect	110	48	111	49
rect	110	50	111	51
rect	110	51	111	52
rect	110	53	111	54
rect	110	54	111	55
rect	110	56	111	57
rect	110	57	111	58
rect	110	59	111	60
rect	110	60	111	61
rect	110	62	111	63
rect	110	63	111	64
rect	110	65	111	66
rect	110	66	111	67
rect	110	68	111	69
rect	110	69	111	70
rect	110	71	111	72
rect	110	72	111	73
rect	110	74	111	75
rect	110	75	111	76
rect	110	77	111	78
rect	110	78	111	79
rect	110	80	111	81
rect	110	81	111	82
rect	110	83	111	84
rect	110	84	111	85
rect	110	86	111	87
rect	110	87	111	88
rect	110	89	111	90
rect	110	90	111	91
rect	110	92	111	93
rect	110	93	111	94
rect	110	95	111	96
rect	110	96	111	97
rect	110	98	111	99
rect	110	99	111	100
rect	110	101	111	102
rect	110	102	111	103
rect	110	104	111	105
rect	110	105	111	106
rect	110	107	111	108
rect	110	108	111	109
rect	110	110	111	111
rect	110	111	111	112
rect	110	113	111	114
rect	110	114	111	115
rect	110	116	111	117
rect	110	117	111	118
rect	110	119	111	120
rect	110	120	111	121
rect	110	122	111	123
rect	110	123	111	124
rect	110	125	111	126
rect	110	126	111	127
rect	110	128	111	129
rect	110	129	111	130
rect	110	131	111	132
rect	110	132	111	133
rect	110	134	111	135
rect	110	135	111	136
rect	110	137	111	138
rect	110	138	111	139
rect	110	140	111	141
rect	110	141	111	142
rect	110	143	111	144
rect	110	144	111	145
rect	110	146	111	147
rect	110	147	111	148
rect	110	149	111	150
rect	110	150	111	151
rect	110	152	111	153
rect	110	153	111	154
rect	110	155	111	156
rect	110	156	111	157
rect	110	158	111	159
rect	110	159	111	160
rect	110	161	111	162
rect	110	162	111	163
rect	110	164	111	165
rect	110	165	111	166
rect	110	167	111	168
rect	110	168	111	169
rect	110	170	111	171
rect	110	171	111	172
rect	110	173	111	174
rect	110	174	111	175
rect	110	176	111	177
rect	110	177	111	178
rect	110	179	111	180
rect	110	180	111	181
rect	110	182	111	183
rect	110	183	111	184
rect	110	185	111	186
rect	110	186	111	187
rect	110	188	111	189
rect	110	189	111	190
rect	110	191	111	192
rect	110	192	111	193
rect	110	194	111	195
rect	110	195	111	196
rect	110	197	111	198
rect	110	198	111	199
rect	110	200	111	201
rect	110	201	111	202
rect	110	203	111	204
rect	110	204	111	205
rect	110	206	111	207
rect	110	207	111	208
rect	110	209	111	210
rect	110	210	111	211
rect	110	212	111	213
rect	110	213	111	214
rect	110	215	111	216
rect	110	216	111	217
rect	110	218	111	219
rect	110	219	111	220
rect	110	221	111	222
rect	110	222	111	223
rect	110	224	111	225
rect	110	225	111	226
rect	110	227	111	228
rect	110	228	111	229
rect	110	230	111	231
rect	110	231	111	232
rect	110	233	111	234
rect	110	234	111	235
rect	110	236	111	237
rect	110	237	111	238
rect	110	239	111	240
rect	110	240	111	241
rect	110	242	111	243
rect	110	243	111	244
rect	110	245	111	246
rect	110	246	111	247
rect	110	248	111	249
rect	110	249	111	250
rect	110	251	111	252
rect	110	252	111	253
rect	110	254	111	255
rect	110	255	111	256
rect	110	257	111	258
rect	110	258	111	259
rect	110	260	111	261
rect	110	261	111	262
rect	110	263	111	264
rect	110	264	111	265
rect	110	266	111	267
rect	110	267	111	268
rect	110	269	111	270
rect	110	270	111	271
rect	110	272	111	273
rect	110	273	111	274
rect	110	275	111	276
rect	110	276	111	277
rect	110	278	111	279
rect	110	279	111	280
rect	110	281	111	282
rect	110	282	111	283
rect	110	284	111	285
rect	110	285	111	286
rect	110	287	111	288
rect	110	288	111	289
rect	110	290	111	291
rect	110	291	111	292
rect	110	293	111	294
rect	110	294	111	295
rect	110	296	111	297
rect	110	297	111	298
rect	110	299	111	300
rect	110	300	111	301
rect	110	302	111	303
rect	110	303	111	304
rect	110	305	111	306
rect	110	306	111	307
rect	110	308	111	309
rect	110	309	111	310
rect	110	311	111	312
rect	110	312	111	313
rect	110	314	111	315
rect	110	315	111	316
rect	110	317	111	318
rect	110	318	111	319
rect	110	320	111	321
rect	110	321	111	322
rect	110	323	111	324
rect	110	324	111	325
rect	110	326	111	327
rect	110	327	111	328
rect	110	329	111	330
rect	110	330	111	331
rect	110	332	111	333
rect	110	333	111	334
rect	110	335	111	336
rect	111	0	112	1
rect	111	2	112	3
rect	111	3	112	4
rect	111	5	112	6
rect	111	6	112	7
rect	111	8	112	9
rect	111	9	112	10
rect	111	11	112	12
rect	111	12	112	13
rect	111	14	112	15
rect	111	15	112	16
rect	111	17	112	18
rect	111	18	112	19
rect	111	20	112	21
rect	111	21	112	22
rect	111	23	112	24
rect	111	24	112	25
rect	111	26	112	27
rect	111	27	112	28
rect	111	29	112	30
rect	111	30	112	31
rect	111	32	112	33
rect	111	33	112	34
rect	111	35	112	36
rect	111	36	112	37
rect	111	38	112	39
rect	111	39	112	40
rect	111	41	112	42
rect	111	42	112	43
rect	111	44	112	45
rect	111	45	112	46
rect	111	47	112	48
rect	111	48	112	49
rect	111	50	112	51
rect	111	51	112	52
rect	111	53	112	54
rect	111	54	112	55
rect	111	56	112	57
rect	111	57	112	58
rect	111	59	112	60
rect	111	60	112	61
rect	111	62	112	63
rect	111	63	112	64
rect	111	65	112	66
rect	111	66	112	67
rect	111	68	112	69
rect	111	69	112	70
rect	111	71	112	72
rect	111	72	112	73
rect	111	74	112	75
rect	111	75	112	76
rect	111	77	112	78
rect	111	78	112	79
rect	111	80	112	81
rect	111	81	112	82
rect	111	83	112	84
rect	111	84	112	85
rect	111	86	112	87
rect	111	87	112	88
rect	111	89	112	90
rect	111	90	112	91
rect	111	92	112	93
rect	111	93	112	94
rect	111	95	112	96
rect	111	96	112	97
rect	111	98	112	99
rect	111	99	112	100
rect	111	101	112	102
rect	111	102	112	103
rect	111	104	112	105
rect	111	105	112	106
rect	111	107	112	108
rect	111	108	112	109
rect	111	110	112	111
rect	111	111	112	112
rect	111	113	112	114
rect	111	114	112	115
rect	111	116	112	117
rect	111	117	112	118
rect	111	119	112	120
rect	111	120	112	121
rect	111	122	112	123
rect	111	123	112	124
rect	111	125	112	126
rect	111	126	112	127
rect	111	128	112	129
rect	111	129	112	130
rect	111	131	112	132
rect	111	132	112	133
rect	111	134	112	135
rect	111	135	112	136
rect	111	137	112	138
rect	111	138	112	139
rect	111	140	112	141
rect	111	141	112	142
rect	111	143	112	144
rect	111	144	112	145
rect	111	146	112	147
rect	111	147	112	148
rect	111	149	112	150
rect	111	150	112	151
rect	111	152	112	153
rect	111	153	112	154
rect	111	155	112	156
rect	111	156	112	157
rect	111	158	112	159
rect	111	159	112	160
rect	111	161	112	162
rect	111	162	112	163
rect	111	164	112	165
rect	111	165	112	166
rect	111	167	112	168
rect	111	168	112	169
rect	111	170	112	171
rect	111	171	112	172
rect	111	173	112	174
rect	111	174	112	175
rect	111	176	112	177
rect	111	177	112	178
rect	111	179	112	180
rect	111	180	112	181
rect	111	182	112	183
rect	111	183	112	184
rect	111	185	112	186
rect	111	186	112	187
rect	111	188	112	189
rect	111	189	112	190
rect	111	191	112	192
rect	111	192	112	193
rect	111	194	112	195
rect	111	195	112	196
rect	111	197	112	198
rect	111	198	112	199
rect	111	200	112	201
rect	111	201	112	202
rect	111	203	112	204
rect	111	204	112	205
rect	111	206	112	207
rect	111	207	112	208
rect	111	209	112	210
rect	111	210	112	211
rect	111	212	112	213
rect	111	213	112	214
rect	111	215	112	216
rect	111	216	112	217
rect	111	218	112	219
rect	111	219	112	220
rect	111	221	112	222
rect	111	222	112	223
rect	111	224	112	225
rect	111	225	112	226
rect	111	227	112	228
rect	111	228	112	229
rect	111	230	112	231
rect	111	231	112	232
rect	111	233	112	234
rect	111	234	112	235
rect	111	236	112	237
rect	111	237	112	238
rect	111	239	112	240
rect	111	240	112	241
rect	111	242	112	243
rect	111	243	112	244
rect	111	245	112	246
rect	111	246	112	247
rect	111	248	112	249
rect	111	249	112	250
rect	111	251	112	252
rect	111	252	112	253
rect	111	254	112	255
rect	111	255	112	256
rect	111	257	112	258
rect	111	258	112	259
rect	111	260	112	261
rect	111	261	112	262
rect	111	263	112	264
rect	111	264	112	265
rect	111	266	112	267
rect	111	267	112	268
rect	111	269	112	270
rect	111	270	112	271
rect	111	272	112	273
rect	111	273	112	274
rect	111	275	112	276
rect	111	276	112	277
rect	111	278	112	279
rect	111	279	112	280
rect	111	281	112	282
rect	111	282	112	283
rect	111	284	112	285
rect	111	285	112	286
rect	111	287	112	288
rect	111	288	112	289
rect	111	290	112	291
rect	111	291	112	292
rect	111	293	112	294
rect	111	294	112	295
rect	111	296	112	297
rect	111	297	112	298
rect	111	299	112	300
rect	111	300	112	301
rect	111	302	112	303
rect	111	303	112	304
rect	111	305	112	306
rect	111	306	112	307
rect	111	308	112	309
rect	111	309	112	310
rect	111	311	112	312
rect	111	312	112	313
rect	111	314	112	315
rect	111	315	112	316
rect	111	317	112	318
rect	111	318	112	319
rect	111	320	112	321
rect	111	321	112	322
rect	111	323	112	324
rect	111	324	112	325
rect	111	326	112	327
rect	111	327	112	328
rect	111	329	112	330
rect	111	330	112	331
rect	111	332	112	333
rect	111	333	112	334
rect	111	335	112	336
rect	112	0	113	1
rect	112	2	113	3
rect	112	3	113	4
rect	112	5	113	6
rect	112	6	113	7
rect	112	8	113	9
rect	112	9	113	10
rect	112	11	113	12
rect	112	12	113	13
rect	112	14	113	15
rect	112	15	113	16
rect	112	17	113	18
rect	112	18	113	19
rect	112	20	113	21
rect	112	21	113	22
rect	112	23	113	24
rect	112	24	113	25
rect	112	26	113	27
rect	112	27	113	28
rect	112	29	113	30
rect	112	30	113	31
rect	112	32	113	33
rect	112	33	113	34
rect	112	35	113	36
rect	112	36	113	37
rect	112	38	113	39
rect	112	39	113	40
rect	112	41	113	42
rect	112	42	113	43
rect	112	44	113	45
rect	112	45	113	46
rect	112	47	113	48
rect	112	48	113	49
rect	112	50	113	51
rect	112	51	113	52
rect	112	53	113	54
rect	112	54	113	55
rect	112	56	113	57
rect	112	57	113	58
rect	112	59	113	60
rect	112	60	113	61
rect	112	62	113	63
rect	112	63	113	64
rect	112	65	113	66
rect	112	66	113	67
rect	112	68	113	69
rect	112	69	113	70
rect	112	71	113	72
rect	112	72	113	73
rect	112	74	113	75
rect	112	75	113	76
rect	112	77	113	78
rect	112	78	113	79
rect	112	80	113	81
rect	112	81	113	82
rect	112	83	113	84
rect	112	84	113	85
rect	112	86	113	87
rect	112	87	113	88
rect	112	89	113	90
rect	112	90	113	91
rect	112	92	113	93
rect	112	93	113	94
rect	112	95	113	96
rect	112	96	113	97
rect	112	98	113	99
rect	112	99	113	100
rect	112	101	113	102
rect	112	102	113	103
rect	112	104	113	105
rect	112	105	113	106
rect	112	107	113	108
rect	112	108	113	109
rect	112	110	113	111
rect	112	111	113	112
rect	112	113	113	114
rect	112	114	113	115
rect	112	116	113	117
rect	112	117	113	118
rect	112	119	113	120
rect	112	120	113	121
rect	112	122	113	123
rect	112	123	113	124
rect	112	125	113	126
rect	112	126	113	127
rect	112	128	113	129
rect	112	129	113	130
rect	112	131	113	132
rect	112	132	113	133
rect	112	134	113	135
rect	112	135	113	136
rect	112	137	113	138
rect	112	138	113	139
rect	112	140	113	141
rect	112	141	113	142
rect	112	143	113	144
rect	112	144	113	145
rect	112	146	113	147
rect	112	147	113	148
rect	112	149	113	150
rect	112	150	113	151
rect	112	152	113	153
rect	112	153	113	154
rect	112	155	113	156
rect	112	156	113	157
rect	112	158	113	159
rect	112	159	113	160
rect	112	161	113	162
rect	112	162	113	163
rect	112	164	113	165
rect	112	165	113	166
rect	112	167	113	168
rect	112	168	113	169
rect	112	170	113	171
rect	112	171	113	172
rect	112	173	113	174
rect	112	174	113	175
rect	112	176	113	177
rect	112	177	113	178
rect	112	179	113	180
rect	112	180	113	181
rect	112	182	113	183
rect	112	183	113	184
rect	112	185	113	186
rect	112	186	113	187
rect	112	188	113	189
rect	112	189	113	190
rect	112	191	113	192
rect	112	192	113	193
rect	112	194	113	195
rect	112	195	113	196
rect	112	197	113	198
rect	112	198	113	199
rect	112	200	113	201
rect	112	201	113	202
rect	112	203	113	204
rect	112	204	113	205
rect	112	206	113	207
rect	112	207	113	208
rect	112	209	113	210
rect	112	210	113	211
rect	112	212	113	213
rect	112	213	113	214
rect	112	215	113	216
rect	112	216	113	217
rect	112	218	113	219
rect	112	219	113	220
rect	112	221	113	222
rect	112	222	113	223
rect	112	224	113	225
rect	112	225	113	226
rect	112	227	113	228
rect	112	228	113	229
rect	112	230	113	231
rect	112	231	113	232
rect	112	233	113	234
rect	112	234	113	235
rect	112	236	113	237
rect	112	237	113	238
rect	112	239	113	240
rect	112	240	113	241
rect	112	242	113	243
rect	112	243	113	244
rect	112	245	113	246
rect	112	246	113	247
rect	112	248	113	249
rect	112	249	113	250
rect	112	251	113	252
rect	112	252	113	253
rect	112	254	113	255
rect	112	255	113	256
rect	112	257	113	258
rect	112	258	113	259
rect	112	260	113	261
rect	112	261	113	262
rect	112	263	113	264
rect	112	264	113	265
rect	112	266	113	267
rect	112	267	113	268
rect	112	269	113	270
rect	112	270	113	271
rect	112	272	113	273
rect	112	273	113	274
rect	112	275	113	276
rect	112	276	113	277
rect	112	278	113	279
rect	112	279	113	280
rect	112	281	113	282
rect	112	282	113	283
rect	112	284	113	285
rect	112	285	113	286
rect	112	287	113	288
rect	112	288	113	289
rect	112	290	113	291
rect	112	291	113	292
rect	112	293	113	294
rect	112	294	113	295
rect	112	296	113	297
rect	112	297	113	298
rect	112	299	113	300
rect	112	300	113	301
rect	112	302	113	303
rect	112	303	113	304
rect	112	305	113	306
rect	112	306	113	307
rect	112	308	113	309
rect	112	309	113	310
rect	112	311	113	312
rect	112	312	113	313
rect	112	314	113	315
rect	112	315	113	316
rect	112	317	113	318
rect	112	318	113	319
rect	112	320	113	321
rect	112	321	113	322
rect	112	323	113	324
rect	112	324	113	325
rect	112	326	113	327
rect	112	327	113	328
rect	112	329	113	330
rect	112	330	113	331
rect	112	332	113	333
rect	112	333	113	334
rect	112	335	113	336
rect	113	0	114	1
rect	113	2	114	3
rect	113	3	114	4
rect	113	5	114	6
rect	113	6	114	7
rect	113	8	114	9
rect	113	9	114	10
rect	113	11	114	12
rect	113	12	114	13
rect	113	14	114	15
rect	113	15	114	16
rect	113	17	114	18
rect	113	18	114	19
rect	113	20	114	21
rect	113	21	114	22
rect	113	23	114	24
rect	113	24	114	25
rect	113	26	114	27
rect	113	27	114	28
rect	113	29	114	30
rect	113	30	114	31
rect	113	32	114	33
rect	113	33	114	34
rect	113	35	114	36
rect	113	36	114	37
rect	113	38	114	39
rect	113	39	114	40
rect	113	41	114	42
rect	113	42	114	43
rect	113	44	114	45
rect	113	45	114	46
rect	113	47	114	48
rect	113	48	114	49
rect	113	50	114	51
rect	113	51	114	52
rect	113	53	114	54
rect	113	54	114	55
rect	113	56	114	57
rect	113	57	114	58
rect	113	59	114	60
rect	113	60	114	61
rect	113	62	114	63
rect	113	63	114	64
rect	113	65	114	66
rect	113	66	114	67
rect	113	68	114	69
rect	113	69	114	70
rect	113	71	114	72
rect	113	72	114	73
rect	113	74	114	75
rect	113	75	114	76
rect	113	77	114	78
rect	113	78	114	79
rect	113	80	114	81
rect	113	81	114	82
rect	113	83	114	84
rect	113	84	114	85
rect	113	86	114	87
rect	113	87	114	88
rect	113	89	114	90
rect	113	90	114	91
rect	113	92	114	93
rect	113	93	114	94
rect	113	95	114	96
rect	113	96	114	97
rect	113	98	114	99
rect	113	99	114	100
rect	113	101	114	102
rect	113	102	114	103
rect	113	104	114	105
rect	113	105	114	106
rect	113	107	114	108
rect	113	108	114	109
rect	113	110	114	111
rect	113	111	114	112
rect	113	113	114	114
rect	113	114	114	115
rect	113	116	114	117
rect	113	117	114	118
rect	113	119	114	120
rect	113	120	114	121
rect	113	122	114	123
rect	113	123	114	124
rect	113	125	114	126
rect	113	126	114	127
rect	113	128	114	129
rect	113	129	114	130
rect	113	131	114	132
rect	113	132	114	133
rect	113	134	114	135
rect	113	135	114	136
rect	113	137	114	138
rect	113	138	114	139
rect	113	140	114	141
rect	113	141	114	142
rect	113	143	114	144
rect	113	144	114	145
rect	113	146	114	147
rect	113	147	114	148
rect	113	149	114	150
rect	113	150	114	151
rect	113	152	114	153
rect	113	153	114	154
rect	113	155	114	156
rect	113	156	114	157
rect	113	158	114	159
rect	113	159	114	160
rect	113	161	114	162
rect	113	162	114	163
rect	113	164	114	165
rect	113	165	114	166
rect	113	167	114	168
rect	113	168	114	169
rect	113	170	114	171
rect	113	171	114	172
rect	113	173	114	174
rect	113	174	114	175
rect	113	176	114	177
rect	113	177	114	178
rect	113	179	114	180
rect	113	180	114	181
rect	113	182	114	183
rect	113	183	114	184
rect	113	185	114	186
rect	113	186	114	187
rect	113	188	114	189
rect	113	189	114	190
rect	113	191	114	192
rect	113	192	114	193
rect	113	194	114	195
rect	113	195	114	196
rect	113	197	114	198
rect	113	198	114	199
rect	113	200	114	201
rect	113	201	114	202
rect	113	203	114	204
rect	113	204	114	205
rect	113	206	114	207
rect	113	207	114	208
rect	113	209	114	210
rect	113	210	114	211
rect	113	212	114	213
rect	113	213	114	214
rect	113	215	114	216
rect	113	216	114	217
rect	113	218	114	219
rect	113	219	114	220
rect	113	221	114	222
rect	113	222	114	223
rect	113	224	114	225
rect	113	225	114	226
rect	113	227	114	228
rect	113	228	114	229
rect	113	230	114	231
rect	113	231	114	232
rect	113	233	114	234
rect	113	234	114	235
rect	113	236	114	237
rect	113	237	114	238
rect	113	239	114	240
rect	113	240	114	241
rect	113	242	114	243
rect	113	243	114	244
rect	113	245	114	246
rect	113	246	114	247
rect	113	248	114	249
rect	113	249	114	250
rect	113	251	114	252
rect	113	252	114	253
rect	113	254	114	255
rect	113	255	114	256
rect	113	257	114	258
rect	113	258	114	259
rect	113	260	114	261
rect	113	261	114	262
rect	113	263	114	264
rect	113	264	114	265
rect	113	266	114	267
rect	113	267	114	268
rect	113	269	114	270
rect	113	270	114	271
rect	113	272	114	273
rect	113	273	114	274
rect	113	275	114	276
rect	113	276	114	277
rect	113	278	114	279
rect	113	279	114	280
rect	113	281	114	282
rect	113	282	114	283
rect	113	284	114	285
rect	113	285	114	286
rect	113	287	114	288
rect	113	288	114	289
rect	113	290	114	291
rect	113	291	114	292
rect	113	293	114	294
rect	113	294	114	295
rect	113	296	114	297
rect	113	297	114	298
rect	113	299	114	300
rect	113	300	114	301
rect	113	302	114	303
rect	113	303	114	304
rect	113	305	114	306
rect	113	306	114	307
rect	113	308	114	309
rect	113	309	114	310
rect	113	311	114	312
rect	113	312	114	313
rect	113	314	114	315
rect	113	315	114	316
rect	113	317	114	318
rect	113	318	114	319
rect	113	320	114	321
rect	113	321	114	322
rect	113	323	114	324
rect	113	324	114	325
rect	113	326	114	327
rect	113	327	114	328
rect	113	329	114	330
rect	113	330	114	331
rect	113	332	114	333
rect	113	333	114	334
rect	113	335	114	336
rect	114	0	115	1
rect	114	2	115	3
rect	114	3	115	4
rect	114	5	115	6
rect	114	6	115	7
rect	114	8	115	9
rect	114	9	115	10
rect	114	11	115	12
rect	114	12	115	13
rect	114	14	115	15
rect	114	15	115	16
rect	114	17	115	18
rect	114	18	115	19
rect	114	20	115	21
rect	114	21	115	22
rect	114	23	115	24
rect	114	24	115	25
rect	114	26	115	27
rect	114	27	115	28
rect	114	29	115	30
rect	114	30	115	31
rect	114	32	115	33
rect	114	33	115	34
rect	114	35	115	36
rect	114	36	115	37
rect	114	38	115	39
rect	114	39	115	40
rect	114	41	115	42
rect	114	42	115	43
rect	114	44	115	45
rect	114	45	115	46
rect	114	47	115	48
rect	114	48	115	49
rect	114	50	115	51
rect	114	51	115	52
rect	114	53	115	54
rect	114	54	115	55
rect	114	56	115	57
rect	114	57	115	58
rect	114	59	115	60
rect	114	60	115	61
rect	114	62	115	63
rect	114	63	115	64
rect	114	65	115	66
rect	114	66	115	67
rect	114	68	115	69
rect	114	69	115	70
rect	114	71	115	72
rect	114	72	115	73
rect	114	74	115	75
rect	114	75	115	76
rect	114	77	115	78
rect	114	78	115	79
rect	114	80	115	81
rect	114	81	115	82
rect	114	83	115	84
rect	114	84	115	85
rect	114	86	115	87
rect	114	87	115	88
rect	114	89	115	90
rect	114	90	115	91
rect	114	92	115	93
rect	114	93	115	94
rect	114	95	115	96
rect	114	96	115	97
rect	114	98	115	99
rect	114	99	115	100
rect	114	101	115	102
rect	114	102	115	103
rect	114	104	115	105
rect	114	105	115	106
rect	114	107	115	108
rect	114	108	115	109
rect	114	110	115	111
rect	114	111	115	112
rect	114	113	115	114
rect	114	114	115	115
rect	114	116	115	117
rect	114	117	115	118
rect	114	119	115	120
rect	114	120	115	121
rect	114	122	115	123
rect	114	123	115	124
rect	114	125	115	126
rect	114	126	115	127
rect	114	128	115	129
rect	114	129	115	130
rect	114	131	115	132
rect	114	132	115	133
rect	114	134	115	135
rect	114	135	115	136
rect	114	137	115	138
rect	114	138	115	139
rect	114	140	115	141
rect	114	141	115	142
rect	114	143	115	144
rect	114	144	115	145
rect	114	146	115	147
rect	114	147	115	148
rect	114	149	115	150
rect	114	150	115	151
rect	114	152	115	153
rect	114	153	115	154
rect	114	155	115	156
rect	114	156	115	157
rect	114	158	115	159
rect	114	159	115	160
rect	114	161	115	162
rect	114	162	115	163
rect	114	164	115	165
rect	114	165	115	166
rect	114	167	115	168
rect	114	168	115	169
rect	114	170	115	171
rect	114	171	115	172
rect	114	173	115	174
rect	114	174	115	175
rect	114	176	115	177
rect	114	177	115	178
rect	114	179	115	180
rect	114	180	115	181
rect	114	182	115	183
rect	114	183	115	184
rect	114	185	115	186
rect	114	186	115	187
rect	114	188	115	189
rect	114	189	115	190
rect	114	191	115	192
rect	114	192	115	193
rect	114	194	115	195
rect	114	195	115	196
rect	114	197	115	198
rect	114	198	115	199
rect	114	200	115	201
rect	114	201	115	202
rect	114	203	115	204
rect	114	204	115	205
rect	114	206	115	207
rect	114	207	115	208
rect	114	209	115	210
rect	114	210	115	211
rect	114	212	115	213
rect	114	213	115	214
rect	114	215	115	216
rect	114	216	115	217
rect	114	218	115	219
rect	114	219	115	220
rect	114	221	115	222
rect	114	222	115	223
rect	114	224	115	225
rect	114	225	115	226
rect	114	227	115	228
rect	114	228	115	229
rect	114	230	115	231
rect	114	231	115	232
rect	114	233	115	234
rect	114	234	115	235
rect	114	236	115	237
rect	114	237	115	238
rect	114	239	115	240
rect	114	240	115	241
rect	114	242	115	243
rect	114	243	115	244
rect	114	245	115	246
rect	114	246	115	247
rect	114	248	115	249
rect	114	249	115	250
rect	114	251	115	252
rect	114	252	115	253
rect	114	254	115	255
rect	114	255	115	256
rect	114	257	115	258
rect	114	258	115	259
rect	114	260	115	261
rect	114	261	115	262
rect	114	263	115	264
rect	114	264	115	265
rect	114	266	115	267
rect	114	267	115	268
rect	114	269	115	270
rect	114	270	115	271
rect	114	272	115	273
rect	114	273	115	274
rect	114	275	115	276
rect	114	276	115	277
rect	114	278	115	279
rect	114	279	115	280
rect	114	281	115	282
rect	114	282	115	283
rect	114	284	115	285
rect	114	285	115	286
rect	114	287	115	288
rect	114	288	115	289
rect	114	290	115	291
rect	114	291	115	292
rect	114	293	115	294
rect	114	294	115	295
rect	114	296	115	297
rect	114	297	115	298
rect	114	299	115	300
rect	114	300	115	301
rect	114	302	115	303
rect	114	303	115	304
rect	114	305	115	306
rect	114	306	115	307
rect	114	308	115	309
rect	114	309	115	310
rect	114	311	115	312
rect	114	312	115	313
rect	114	314	115	315
rect	114	315	115	316
rect	114	317	115	318
rect	114	318	115	319
rect	114	320	115	321
rect	114	321	115	322
rect	114	323	115	324
rect	114	324	115	325
rect	114	326	115	327
rect	114	327	115	328
rect	114	329	115	330
rect	114	330	115	331
rect	114	332	115	333
rect	114	333	115	334
rect	114	335	115	336
rect	119	0	120	1
rect	119	2	120	3
rect	119	3	120	4
rect	119	5	120	6
rect	119	6	120	7
rect	119	8	120	9
rect	119	9	120	10
rect	119	11	120	12
rect	119	12	120	13
rect	119	14	120	15
rect	119	15	120	16
rect	119	17	120	18
rect	119	18	120	19
rect	119	20	120	21
rect	119	21	120	22
rect	119	23	120	24
rect	119	24	120	25
rect	119	26	120	27
rect	119	27	120	28
rect	119	29	120	30
rect	119	30	120	31
rect	119	32	120	33
rect	119	33	120	34
rect	119	35	120	36
rect	119	36	120	37
rect	119	38	120	39
rect	119	39	120	40
rect	119	41	120	42
rect	119	42	120	43
rect	119	44	120	45
rect	119	45	120	46
rect	119	47	120	48
rect	119	48	120	49
rect	119	50	120	51
rect	119	51	120	52
rect	119	53	120	54
rect	119	54	120	55
rect	119	56	120	57
rect	119	57	120	58
rect	119	59	120	60
rect	119	60	120	61
rect	119	62	120	63
rect	119	63	120	64
rect	119	65	120	66
rect	119	66	120	67
rect	119	68	120	69
rect	119	69	120	70
rect	119	71	120	72
rect	119	72	120	73
rect	119	74	120	75
rect	119	75	120	76
rect	119	77	120	78
rect	119	78	120	79
rect	119	80	120	81
rect	119	81	120	82
rect	119	83	120	84
rect	119	84	120	85
rect	119	86	120	87
rect	119	87	120	88
rect	119	89	120	90
rect	119	90	120	91
rect	119	92	120	93
rect	119	93	120	94
rect	119	95	120	96
rect	119	96	120	97
rect	119	98	120	99
rect	119	99	120	100
rect	119	101	120	102
rect	119	102	120	103
rect	119	104	120	105
rect	119	105	120	106
rect	119	107	120	108
rect	119	108	120	109
rect	119	110	120	111
rect	119	111	120	112
rect	119	113	120	114
rect	119	114	120	115
rect	119	116	120	117
rect	119	117	120	118
rect	119	119	120	120
rect	119	120	120	121
rect	119	122	120	123
rect	119	123	120	124
rect	119	125	120	126
rect	119	126	120	127
rect	119	128	120	129
rect	119	129	120	130
rect	119	131	120	132
rect	119	132	120	133
rect	119	134	120	135
rect	119	135	120	136
rect	119	137	120	138
rect	119	138	120	139
rect	119	140	120	141
rect	119	141	120	142
rect	119	143	120	144
rect	119	144	120	145
rect	119	146	120	147
rect	119	147	120	148
rect	119	149	120	150
rect	119	150	120	151
rect	119	152	120	153
rect	119	153	120	154
rect	119	155	120	156
rect	119	156	120	157
rect	119	158	120	159
rect	119	159	120	160
rect	119	161	120	162
rect	119	162	120	163
rect	119	164	120	165
rect	119	165	120	166
rect	119	167	120	168
rect	119	168	120	169
rect	119	170	120	171
rect	119	171	120	172
rect	119	173	120	174
rect	119	174	120	175
rect	119	176	120	177
rect	119	177	120	178
rect	119	179	120	180
rect	119	180	120	181
rect	119	182	120	183
rect	119	183	120	184
rect	119	185	120	186
rect	119	186	120	187
rect	119	188	120	189
rect	119	189	120	190
rect	119	191	120	192
rect	119	192	120	193
rect	119	194	120	195
rect	119	195	120	196
rect	119	197	120	198
rect	119	198	120	199
rect	119	200	120	201
rect	119	201	120	202
rect	119	203	120	204
rect	119	204	120	205
rect	119	206	120	207
rect	119	207	120	208
rect	119	209	120	210
rect	119	210	120	211
rect	119	212	120	213
rect	119	213	120	214
rect	119	215	120	216
rect	119	216	120	217
rect	119	218	120	219
rect	119	219	120	220
rect	119	221	120	222
rect	119	222	120	223
rect	119	224	120	225
rect	119	225	120	226
rect	119	227	120	228
rect	119	228	120	229
rect	119	230	120	231
rect	119	231	120	232
rect	119	233	120	234
rect	119	234	120	235
rect	119	236	120	237
rect	119	237	120	238
rect	119	239	120	240
rect	119	240	120	241
rect	119	242	120	243
rect	119	243	120	244
rect	119	245	120	246
rect	119	246	120	247
rect	119	248	120	249
rect	119	249	120	250
rect	119	251	120	252
rect	119	252	120	253
rect	119	254	120	255
rect	119	255	120	256
rect	119	257	120	258
rect	119	258	120	259
rect	119	260	120	261
rect	119	261	120	262
rect	119	263	120	264
rect	119	264	120	265
rect	119	266	120	267
rect	119	267	120	268
rect	119	269	120	270
rect	119	270	120	271
rect	119	272	120	273
rect	119	273	120	274
rect	119	275	120	276
rect	119	276	120	277
rect	119	278	120	279
rect	119	279	120	280
rect	119	281	120	282
rect	119	282	120	283
rect	119	284	120	285
rect	119	285	120	286
rect	119	287	120	288
rect	119	288	120	289
rect	119	290	120	291
rect	119	291	120	292
rect	119	293	120	294
rect	119	294	120	295
rect	119	296	120	297
rect	119	297	120	298
rect	119	299	120	300
rect	119	300	120	301
rect	119	302	120	303
rect	119	303	120	304
rect	119	305	120	306
rect	119	306	120	307
rect	119	308	120	309
rect	119	309	120	310
rect	119	311	120	312
rect	119	312	120	313
rect	119	314	120	315
rect	119	315	120	316
rect	119	317	120	318
rect	119	318	120	319
rect	119	320	120	321
rect	119	321	120	322
rect	119	323	120	324
rect	119	324	120	325
rect	119	326	120	327
rect	119	327	120	328
rect	119	329	120	330
rect	119	330	120	331
rect	119	332	120	333
rect	119	333	120	334
rect	119	335	120	336
rect	121	0	122	1
rect	121	2	122	3
rect	121	3	122	4
rect	121	5	122	6
rect	121	6	122	7
rect	121	8	122	9
rect	121	9	122	10
rect	121	11	122	12
rect	121	12	122	13
rect	121	14	122	15
rect	121	15	122	16
rect	121	17	122	18
rect	121	18	122	19
rect	121	20	122	21
rect	121	21	122	22
rect	121	23	122	24
rect	121	24	122	25
rect	121	26	122	27
rect	121	27	122	28
rect	121	29	122	30
rect	121	30	122	31
rect	121	32	122	33
rect	121	33	122	34
rect	121	35	122	36
rect	121	36	122	37
rect	121	38	122	39
rect	121	39	122	40
rect	121	41	122	42
rect	121	42	122	43
rect	121	44	122	45
rect	121	45	122	46
rect	121	47	122	48
rect	121	48	122	49
rect	121	50	122	51
rect	121	51	122	52
rect	121	53	122	54
rect	121	54	122	55
rect	121	56	122	57
rect	121	57	122	58
rect	121	59	122	60
rect	121	60	122	61
rect	121	62	122	63
rect	121	63	122	64
rect	121	65	122	66
rect	121	66	122	67
rect	121	68	122	69
rect	121	69	122	70
rect	121	71	122	72
rect	121	72	122	73
rect	121	74	122	75
rect	121	75	122	76
rect	121	77	122	78
rect	121	78	122	79
rect	121	80	122	81
rect	121	81	122	82
rect	121	83	122	84
rect	121	84	122	85
rect	121	86	122	87
rect	121	87	122	88
rect	121	89	122	90
rect	121	90	122	91
rect	121	92	122	93
rect	121	93	122	94
rect	121	95	122	96
rect	121	96	122	97
rect	121	98	122	99
rect	121	99	122	100
rect	121	101	122	102
rect	121	102	122	103
rect	121	104	122	105
rect	121	105	122	106
rect	121	107	122	108
rect	121	108	122	109
rect	121	110	122	111
rect	121	111	122	112
rect	121	113	122	114
rect	121	114	122	115
rect	121	116	122	117
rect	121	117	122	118
rect	121	119	122	120
rect	121	120	122	121
rect	121	122	122	123
rect	121	123	122	124
rect	121	125	122	126
rect	121	126	122	127
rect	121	128	122	129
rect	121	129	122	130
rect	121	131	122	132
rect	121	132	122	133
rect	121	134	122	135
rect	121	135	122	136
rect	121	137	122	138
rect	121	138	122	139
rect	121	140	122	141
rect	121	141	122	142
rect	121	143	122	144
rect	121	144	122	145
rect	121	146	122	147
rect	121	147	122	148
rect	121	149	122	150
rect	121	150	122	151
rect	121	152	122	153
rect	121	153	122	154
rect	121	155	122	156
rect	121	156	122	157
rect	121	158	122	159
rect	121	159	122	160
rect	121	161	122	162
rect	121	162	122	163
rect	121	164	122	165
rect	121	165	122	166
rect	121	167	122	168
rect	121	168	122	169
rect	121	170	122	171
rect	121	171	122	172
rect	121	173	122	174
rect	121	174	122	175
rect	121	176	122	177
rect	121	177	122	178
rect	121	179	122	180
rect	121	180	122	181
rect	121	182	122	183
rect	121	183	122	184
rect	121	185	122	186
rect	121	186	122	187
rect	121	188	122	189
rect	121	189	122	190
rect	121	191	122	192
rect	121	192	122	193
rect	121	194	122	195
rect	121	195	122	196
rect	121	197	122	198
rect	121	198	122	199
rect	121	200	122	201
rect	121	201	122	202
rect	121	203	122	204
rect	121	204	122	205
rect	121	206	122	207
rect	121	207	122	208
rect	121	209	122	210
rect	121	210	122	211
rect	121	212	122	213
rect	121	213	122	214
rect	121	215	122	216
rect	121	216	122	217
rect	121	218	122	219
rect	121	219	122	220
rect	121	221	122	222
rect	121	222	122	223
rect	121	224	122	225
rect	121	225	122	226
rect	121	227	122	228
rect	121	228	122	229
rect	121	230	122	231
rect	121	231	122	232
rect	121	233	122	234
rect	121	234	122	235
rect	121	236	122	237
rect	121	237	122	238
rect	121	239	122	240
rect	121	240	122	241
rect	121	242	122	243
rect	121	243	122	244
rect	121	245	122	246
rect	121	246	122	247
rect	121	248	122	249
rect	121	249	122	250
rect	121	251	122	252
rect	121	252	122	253
rect	121	254	122	255
rect	121	255	122	256
rect	121	257	122	258
rect	121	258	122	259
rect	121	260	122	261
rect	121	261	122	262
rect	121	263	122	264
rect	121	264	122	265
rect	121	266	122	267
rect	121	267	122	268
rect	121	269	122	270
rect	121	270	122	271
rect	121	272	122	273
rect	121	273	122	274
rect	121	275	122	276
rect	121	276	122	277
rect	121	278	122	279
rect	121	279	122	280
rect	121	281	122	282
rect	121	282	122	283
rect	121	284	122	285
rect	121	285	122	286
rect	121	287	122	288
rect	121	288	122	289
rect	121	290	122	291
rect	121	291	122	292
rect	121	293	122	294
rect	121	294	122	295
rect	121	296	122	297
rect	121	297	122	298
rect	121	299	122	300
rect	121	300	122	301
rect	121	302	122	303
rect	121	303	122	304
rect	121	305	122	306
rect	121	306	122	307
rect	121	308	122	309
rect	121	309	122	310
rect	121	311	122	312
rect	121	312	122	313
rect	121	314	122	315
rect	121	315	122	316
rect	121	317	122	318
rect	121	318	122	319
rect	121	320	122	321
rect	121	321	122	322
rect	121	323	122	324
rect	121	324	122	325
rect	121	326	122	327
rect	121	327	122	328
rect	121	329	122	330
rect	121	330	122	331
rect	121	332	122	333
rect	121	333	122	334
rect	121	335	122	336
rect	121	336	122	337
rect	121	338	122	339
rect	121	339	122	340
rect	121	341	122	342
rect	121	342	122	343
rect	121	344	122	345
rect	121	345	122	346
rect	121	347	122	348
rect	121	348	122	349
rect	121	350	122	351
rect	121	351	122	352
rect	121	353	122	354
rect	121	354	122	355
rect	121	356	122	357
rect	121	357	122	358
rect	121	359	122	360
rect	121	360	122	361
rect	121	362	122	363
rect	121	363	122	364
rect	121	365	122	366
rect	122	0	123	1
rect	122	2	123	3
rect	122	3	123	4
rect	122	5	123	6
rect	122	6	123	7
rect	122	8	123	9
rect	122	9	123	10
rect	122	11	123	12
rect	122	12	123	13
rect	122	14	123	15
rect	122	15	123	16
rect	122	17	123	18
rect	122	18	123	19
rect	122	20	123	21
rect	122	21	123	22
rect	122	23	123	24
rect	122	24	123	25
rect	122	26	123	27
rect	122	27	123	28
rect	122	29	123	30
rect	122	30	123	31
rect	122	32	123	33
rect	122	33	123	34
rect	122	35	123	36
rect	122	36	123	37
rect	122	38	123	39
rect	122	39	123	40
rect	122	41	123	42
rect	122	42	123	43
rect	122	44	123	45
rect	122	45	123	46
rect	122	47	123	48
rect	122	48	123	49
rect	122	50	123	51
rect	122	51	123	52
rect	122	53	123	54
rect	122	54	123	55
rect	122	56	123	57
rect	122	57	123	58
rect	122	59	123	60
rect	122	60	123	61
rect	122	62	123	63
rect	122	63	123	64
rect	122	65	123	66
rect	122	66	123	67
rect	122	68	123	69
rect	122	69	123	70
rect	122	71	123	72
rect	122	72	123	73
rect	122	74	123	75
rect	122	75	123	76
rect	122	77	123	78
rect	122	78	123	79
rect	122	80	123	81
rect	122	81	123	82
rect	122	83	123	84
rect	122	84	123	85
rect	122	86	123	87
rect	122	87	123	88
rect	122	89	123	90
rect	122	90	123	91
rect	122	92	123	93
rect	122	93	123	94
rect	122	95	123	96
rect	122	96	123	97
rect	122	98	123	99
rect	122	99	123	100
rect	122	101	123	102
rect	122	102	123	103
rect	122	104	123	105
rect	122	105	123	106
rect	122	107	123	108
rect	122	108	123	109
rect	122	110	123	111
rect	122	111	123	112
rect	122	113	123	114
rect	122	114	123	115
rect	122	116	123	117
rect	122	117	123	118
rect	122	119	123	120
rect	122	120	123	121
rect	122	122	123	123
rect	122	123	123	124
rect	122	125	123	126
rect	122	126	123	127
rect	122	128	123	129
rect	122	129	123	130
rect	122	131	123	132
rect	122	132	123	133
rect	122	134	123	135
rect	122	135	123	136
rect	122	137	123	138
rect	122	138	123	139
rect	122	140	123	141
rect	122	141	123	142
rect	122	143	123	144
rect	122	144	123	145
rect	122	146	123	147
rect	122	147	123	148
rect	122	149	123	150
rect	122	150	123	151
rect	122	152	123	153
rect	122	153	123	154
rect	122	155	123	156
rect	122	156	123	157
rect	122	158	123	159
rect	122	159	123	160
rect	122	161	123	162
rect	122	162	123	163
rect	122	164	123	165
rect	122	165	123	166
rect	122	167	123	168
rect	122	168	123	169
rect	122	170	123	171
rect	122	171	123	172
rect	122	173	123	174
rect	122	174	123	175
rect	122	176	123	177
rect	122	177	123	178
rect	122	179	123	180
rect	122	180	123	181
rect	122	182	123	183
rect	122	183	123	184
rect	122	185	123	186
rect	122	186	123	187
rect	122	188	123	189
rect	122	189	123	190
rect	122	191	123	192
rect	122	192	123	193
rect	122	194	123	195
rect	122	195	123	196
rect	122	197	123	198
rect	122	198	123	199
rect	122	200	123	201
rect	122	201	123	202
rect	122	203	123	204
rect	122	204	123	205
rect	122	206	123	207
rect	122	207	123	208
rect	122	209	123	210
rect	122	210	123	211
rect	122	212	123	213
rect	122	213	123	214
rect	122	215	123	216
rect	122	216	123	217
rect	122	218	123	219
rect	122	219	123	220
rect	122	221	123	222
rect	122	222	123	223
rect	122	224	123	225
rect	122	225	123	226
rect	122	227	123	228
rect	122	228	123	229
rect	122	230	123	231
rect	122	231	123	232
rect	122	233	123	234
rect	122	234	123	235
rect	122	236	123	237
rect	122	237	123	238
rect	122	239	123	240
rect	122	240	123	241
rect	122	242	123	243
rect	122	243	123	244
rect	122	245	123	246
rect	122	246	123	247
rect	122	248	123	249
rect	122	249	123	250
rect	122	251	123	252
rect	122	252	123	253
rect	122	254	123	255
rect	122	255	123	256
rect	122	257	123	258
rect	122	258	123	259
rect	122	260	123	261
rect	122	261	123	262
rect	122	263	123	264
rect	122	264	123	265
rect	122	266	123	267
rect	122	267	123	268
rect	122	269	123	270
rect	122	270	123	271
rect	122	272	123	273
rect	122	273	123	274
rect	122	275	123	276
rect	122	276	123	277
rect	122	278	123	279
rect	122	279	123	280
rect	122	281	123	282
rect	122	282	123	283
rect	122	284	123	285
rect	122	285	123	286
rect	122	287	123	288
rect	122	288	123	289
rect	122	290	123	291
rect	122	291	123	292
rect	122	293	123	294
rect	122	294	123	295
rect	122	296	123	297
rect	122	297	123	298
rect	122	299	123	300
rect	122	300	123	301
rect	122	302	123	303
rect	122	303	123	304
rect	122	305	123	306
rect	122	306	123	307
rect	122	308	123	309
rect	122	309	123	310
rect	122	311	123	312
rect	122	312	123	313
rect	122	314	123	315
rect	122	315	123	316
rect	122	317	123	318
rect	122	318	123	319
rect	122	320	123	321
rect	122	321	123	322
rect	122	323	123	324
rect	122	324	123	325
rect	122	326	123	327
rect	122	327	123	328
rect	122	329	123	330
rect	122	330	123	331
rect	122	332	123	333
rect	122	333	123	334
rect	122	335	123	336
rect	122	336	123	337
rect	122	338	123	339
rect	122	339	123	340
rect	122	341	123	342
rect	122	342	123	343
rect	122	344	123	345
rect	122	345	123	346
rect	122	347	123	348
rect	122	348	123	349
rect	122	350	123	351
rect	122	351	123	352
rect	122	353	123	354
rect	122	354	123	355
rect	122	356	123	357
rect	122	357	123	358
rect	122	359	123	360
rect	122	360	123	361
rect	122	362	123	363
rect	122	363	123	364
rect	122	365	123	366
rect	123	0	124	1
rect	123	2	124	3
rect	123	3	124	4
rect	123	5	124	6
rect	123	6	124	7
rect	123	8	124	9
rect	123	9	124	10
rect	123	11	124	12
rect	123	12	124	13
rect	123	14	124	15
rect	123	15	124	16
rect	123	17	124	18
rect	123	18	124	19
rect	123	20	124	21
rect	123	21	124	22
rect	123	23	124	24
rect	123	24	124	25
rect	123	26	124	27
rect	123	27	124	28
rect	123	29	124	30
rect	123	30	124	31
rect	123	32	124	33
rect	123	33	124	34
rect	123	35	124	36
rect	123	36	124	37
rect	123	38	124	39
rect	123	39	124	40
rect	123	41	124	42
rect	123	42	124	43
rect	123	44	124	45
rect	123	45	124	46
rect	123	47	124	48
rect	123	48	124	49
rect	123	50	124	51
rect	123	51	124	52
rect	123	53	124	54
rect	123	54	124	55
rect	123	56	124	57
rect	123	57	124	58
rect	123	59	124	60
rect	123	60	124	61
rect	123	62	124	63
rect	123	63	124	64
rect	123	65	124	66
rect	123	66	124	67
rect	123	68	124	69
rect	123	69	124	70
rect	123	71	124	72
rect	123	72	124	73
rect	123	74	124	75
rect	123	75	124	76
rect	123	77	124	78
rect	123	78	124	79
rect	123	80	124	81
rect	123	81	124	82
rect	123	83	124	84
rect	123	84	124	85
rect	123	86	124	87
rect	123	87	124	88
rect	123	89	124	90
rect	123	90	124	91
rect	123	92	124	93
rect	123	93	124	94
rect	123	95	124	96
rect	123	96	124	97
rect	123	98	124	99
rect	123	99	124	100
rect	123	101	124	102
rect	123	102	124	103
rect	123	104	124	105
rect	123	105	124	106
rect	123	107	124	108
rect	123	108	124	109
rect	123	110	124	111
rect	123	111	124	112
rect	123	113	124	114
rect	123	114	124	115
rect	123	116	124	117
rect	123	117	124	118
rect	123	119	124	120
rect	123	120	124	121
rect	123	122	124	123
rect	123	123	124	124
rect	123	125	124	126
rect	123	126	124	127
rect	123	128	124	129
rect	123	129	124	130
rect	123	131	124	132
rect	123	132	124	133
rect	123	134	124	135
rect	123	135	124	136
rect	123	137	124	138
rect	123	138	124	139
rect	123	140	124	141
rect	123	141	124	142
rect	123	143	124	144
rect	123	144	124	145
rect	123	146	124	147
rect	123	147	124	148
rect	123	149	124	150
rect	123	150	124	151
rect	123	152	124	153
rect	123	153	124	154
rect	123	155	124	156
rect	123	156	124	157
rect	123	158	124	159
rect	123	159	124	160
rect	123	161	124	162
rect	123	162	124	163
rect	123	164	124	165
rect	123	165	124	166
rect	123	167	124	168
rect	123	168	124	169
rect	123	170	124	171
rect	123	171	124	172
rect	123	173	124	174
rect	123	174	124	175
rect	123	176	124	177
rect	123	177	124	178
rect	123	179	124	180
rect	123	180	124	181
rect	123	182	124	183
rect	123	183	124	184
rect	123	185	124	186
rect	123	186	124	187
rect	123	188	124	189
rect	123	189	124	190
rect	123	191	124	192
rect	123	192	124	193
rect	123	194	124	195
rect	123	195	124	196
rect	123	197	124	198
rect	123	198	124	199
rect	123	200	124	201
rect	123	201	124	202
rect	123	203	124	204
rect	123	204	124	205
rect	123	206	124	207
rect	123	207	124	208
rect	123	209	124	210
rect	123	210	124	211
rect	123	212	124	213
rect	123	213	124	214
rect	123	215	124	216
rect	123	216	124	217
rect	123	218	124	219
rect	123	219	124	220
rect	123	221	124	222
rect	123	222	124	223
rect	123	224	124	225
rect	123	225	124	226
rect	123	227	124	228
rect	123	228	124	229
rect	123	230	124	231
rect	123	231	124	232
rect	123	233	124	234
rect	123	234	124	235
rect	123	236	124	237
rect	123	237	124	238
rect	123	239	124	240
rect	123	240	124	241
rect	123	242	124	243
rect	123	243	124	244
rect	123	245	124	246
rect	123	246	124	247
rect	123	248	124	249
rect	123	249	124	250
rect	123	251	124	252
rect	123	252	124	253
rect	123	254	124	255
rect	123	255	124	256
rect	123	257	124	258
rect	123	258	124	259
rect	123	260	124	261
rect	123	261	124	262
rect	123	263	124	264
rect	123	264	124	265
rect	123	266	124	267
rect	123	267	124	268
rect	123	269	124	270
rect	123	270	124	271
rect	123	272	124	273
rect	123	273	124	274
rect	123	275	124	276
rect	123	276	124	277
rect	123	278	124	279
rect	123	279	124	280
rect	123	281	124	282
rect	123	282	124	283
rect	123	284	124	285
rect	123	285	124	286
rect	123	287	124	288
rect	123	288	124	289
rect	123	290	124	291
rect	123	291	124	292
rect	123	293	124	294
rect	123	294	124	295
rect	123	296	124	297
rect	123	297	124	298
rect	123	299	124	300
rect	123	300	124	301
rect	123	302	124	303
rect	123	303	124	304
rect	123	305	124	306
rect	123	306	124	307
rect	123	308	124	309
rect	123	309	124	310
rect	123	311	124	312
rect	123	312	124	313
rect	123	314	124	315
rect	123	315	124	316
rect	123	317	124	318
rect	123	318	124	319
rect	123	320	124	321
rect	123	321	124	322
rect	123	323	124	324
rect	123	324	124	325
rect	123	326	124	327
rect	123	327	124	328
rect	123	329	124	330
rect	123	330	124	331
rect	123	332	124	333
rect	123	333	124	334
rect	123	335	124	336
rect	123	336	124	337
rect	123	338	124	339
rect	123	339	124	340
rect	123	341	124	342
rect	123	342	124	343
rect	123	344	124	345
rect	123	345	124	346
rect	123	347	124	348
rect	123	348	124	349
rect	123	350	124	351
rect	123	351	124	352
rect	123	353	124	354
rect	123	354	124	355
rect	123	356	124	357
rect	123	357	124	358
rect	123	359	124	360
rect	123	360	124	361
rect	123	362	124	363
rect	123	363	124	364
rect	123	365	124	366
rect	124	0	125	1
rect	124	2	125	3
rect	124	3	125	4
rect	124	5	125	6
rect	124	6	125	7
rect	124	8	125	9
rect	124	9	125	10
rect	124	11	125	12
rect	124	12	125	13
rect	124	14	125	15
rect	124	15	125	16
rect	124	17	125	18
rect	124	18	125	19
rect	124	20	125	21
rect	124	21	125	22
rect	124	23	125	24
rect	124	24	125	25
rect	124	26	125	27
rect	124	27	125	28
rect	124	29	125	30
rect	124	30	125	31
rect	124	32	125	33
rect	124	33	125	34
rect	124	35	125	36
rect	124	36	125	37
rect	124	38	125	39
rect	124	39	125	40
rect	124	41	125	42
rect	124	42	125	43
rect	124	44	125	45
rect	124	45	125	46
rect	124	47	125	48
rect	124	48	125	49
rect	124	50	125	51
rect	124	51	125	52
rect	124	53	125	54
rect	124	54	125	55
rect	124	56	125	57
rect	124	57	125	58
rect	124	59	125	60
rect	124	60	125	61
rect	124	62	125	63
rect	124	63	125	64
rect	124	65	125	66
rect	124	66	125	67
rect	124	68	125	69
rect	124	69	125	70
rect	124	71	125	72
rect	124	72	125	73
rect	124	74	125	75
rect	124	75	125	76
rect	124	77	125	78
rect	124	78	125	79
rect	124	80	125	81
rect	124	81	125	82
rect	124	83	125	84
rect	124	84	125	85
rect	124	86	125	87
rect	124	87	125	88
rect	124	89	125	90
rect	124	90	125	91
rect	124	92	125	93
rect	124	93	125	94
rect	124	95	125	96
rect	124	96	125	97
rect	124	98	125	99
rect	124	99	125	100
rect	124	101	125	102
rect	124	102	125	103
rect	124	104	125	105
rect	124	105	125	106
rect	124	107	125	108
rect	124	108	125	109
rect	124	110	125	111
rect	124	111	125	112
rect	124	113	125	114
rect	124	114	125	115
rect	124	116	125	117
rect	124	117	125	118
rect	124	119	125	120
rect	124	120	125	121
rect	124	122	125	123
rect	124	123	125	124
rect	124	125	125	126
rect	124	126	125	127
rect	124	128	125	129
rect	124	129	125	130
rect	124	131	125	132
rect	124	132	125	133
rect	124	134	125	135
rect	124	135	125	136
rect	124	137	125	138
rect	124	138	125	139
rect	124	140	125	141
rect	124	141	125	142
rect	124	143	125	144
rect	124	144	125	145
rect	124	146	125	147
rect	124	147	125	148
rect	124	149	125	150
rect	124	150	125	151
rect	124	152	125	153
rect	124	153	125	154
rect	124	155	125	156
rect	124	156	125	157
rect	124	158	125	159
rect	124	159	125	160
rect	124	161	125	162
rect	124	162	125	163
rect	124	164	125	165
rect	124	165	125	166
rect	124	167	125	168
rect	124	168	125	169
rect	124	170	125	171
rect	124	171	125	172
rect	124	173	125	174
rect	124	174	125	175
rect	124	176	125	177
rect	124	177	125	178
rect	124	179	125	180
rect	124	180	125	181
rect	124	182	125	183
rect	124	183	125	184
rect	124	185	125	186
rect	124	186	125	187
rect	124	188	125	189
rect	124	189	125	190
rect	124	191	125	192
rect	124	192	125	193
rect	124	194	125	195
rect	124	195	125	196
rect	124	197	125	198
rect	124	198	125	199
rect	124	200	125	201
rect	124	201	125	202
rect	124	203	125	204
rect	124	204	125	205
rect	124	206	125	207
rect	124	207	125	208
rect	124	209	125	210
rect	124	210	125	211
rect	124	212	125	213
rect	124	213	125	214
rect	124	215	125	216
rect	124	216	125	217
rect	124	218	125	219
rect	124	219	125	220
rect	124	221	125	222
rect	124	222	125	223
rect	124	224	125	225
rect	124	225	125	226
rect	124	227	125	228
rect	124	228	125	229
rect	124	230	125	231
rect	124	231	125	232
rect	124	233	125	234
rect	124	234	125	235
rect	124	236	125	237
rect	124	237	125	238
rect	124	239	125	240
rect	124	240	125	241
rect	124	242	125	243
rect	124	243	125	244
rect	124	245	125	246
rect	124	246	125	247
rect	124	248	125	249
rect	124	249	125	250
rect	124	251	125	252
rect	124	252	125	253
rect	124	254	125	255
rect	124	255	125	256
rect	124	257	125	258
rect	124	258	125	259
rect	124	260	125	261
rect	124	261	125	262
rect	124	263	125	264
rect	124	264	125	265
rect	124	266	125	267
rect	124	267	125	268
rect	124	269	125	270
rect	124	270	125	271
rect	124	272	125	273
rect	124	273	125	274
rect	124	275	125	276
rect	124	276	125	277
rect	124	278	125	279
rect	124	279	125	280
rect	124	281	125	282
rect	124	282	125	283
rect	124	284	125	285
rect	124	285	125	286
rect	124	287	125	288
rect	124	288	125	289
rect	124	290	125	291
rect	124	291	125	292
rect	124	293	125	294
rect	124	294	125	295
rect	124	296	125	297
rect	124	297	125	298
rect	124	299	125	300
rect	124	300	125	301
rect	124	302	125	303
rect	124	303	125	304
rect	124	305	125	306
rect	124	306	125	307
rect	124	308	125	309
rect	124	309	125	310
rect	124	311	125	312
rect	124	312	125	313
rect	124	314	125	315
rect	124	315	125	316
rect	124	317	125	318
rect	124	318	125	319
rect	124	320	125	321
rect	124	321	125	322
rect	124	323	125	324
rect	124	324	125	325
rect	124	326	125	327
rect	124	327	125	328
rect	124	329	125	330
rect	124	330	125	331
rect	124	332	125	333
rect	124	333	125	334
rect	124	335	125	336
rect	124	336	125	337
rect	124	338	125	339
rect	124	339	125	340
rect	124	341	125	342
rect	124	342	125	343
rect	124	344	125	345
rect	124	345	125	346
rect	124	347	125	348
rect	124	348	125	349
rect	124	350	125	351
rect	124	351	125	352
rect	124	353	125	354
rect	124	354	125	355
rect	124	356	125	357
rect	124	357	125	358
rect	124	359	125	360
rect	124	360	125	361
rect	124	362	125	363
rect	124	363	125	364
rect	124	365	125	366
rect	125	0	126	1
rect	125	2	126	3
rect	125	3	126	4
rect	125	5	126	6
rect	125	6	126	7
rect	125	8	126	9
rect	125	9	126	10
rect	125	11	126	12
rect	125	12	126	13
rect	125	14	126	15
rect	125	15	126	16
rect	125	17	126	18
rect	125	18	126	19
rect	125	20	126	21
rect	125	21	126	22
rect	125	23	126	24
rect	125	24	126	25
rect	125	26	126	27
rect	125	27	126	28
rect	125	29	126	30
rect	125	30	126	31
rect	125	32	126	33
rect	125	33	126	34
rect	125	35	126	36
rect	125	36	126	37
rect	125	38	126	39
rect	125	39	126	40
rect	125	41	126	42
rect	125	42	126	43
rect	125	44	126	45
rect	125	45	126	46
rect	125	47	126	48
rect	125	48	126	49
rect	125	50	126	51
rect	125	51	126	52
rect	125	53	126	54
rect	125	54	126	55
rect	125	56	126	57
rect	125	57	126	58
rect	125	59	126	60
rect	125	60	126	61
rect	125	62	126	63
rect	125	63	126	64
rect	125	65	126	66
rect	125	66	126	67
rect	125	68	126	69
rect	125	69	126	70
rect	125	71	126	72
rect	125	72	126	73
rect	125	74	126	75
rect	125	75	126	76
rect	125	77	126	78
rect	125	78	126	79
rect	125	80	126	81
rect	125	81	126	82
rect	125	83	126	84
rect	125	84	126	85
rect	125	86	126	87
rect	125	87	126	88
rect	125	89	126	90
rect	125	90	126	91
rect	125	92	126	93
rect	125	93	126	94
rect	125	95	126	96
rect	125	96	126	97
rect	125	98	126	99
rect	125	99	126	100
rect	125	101	126	102
rect	125	102	126	103
rect	125	104	126	105
rect	125	105	126	106
rect	125	107	126	108
rect	125	108	126	109
rect	125	110	126	111
rect	125	111	126	112
rect	125	113	126	114
rect	125	114	126	115
rect	125	116	126	117
rect	125	117	126	118
rect	125	119	126	120
rect	125	120	126	121
rect	125	122	126	123
rect	125	123	126	124
rect	125	125	126	126
rect	125	126	126	127
rect	125	128	126	129
rect	125	129	126	130
rect	125	131	126	132
rect	125	132	126	133
rect	125	134	126	135
rect	125	135	126	136
rect	125	137	126	138
rect	125	138	126	139
rect	125	140	126	141
rect	125	141	126	142
rect	125	143	126	144
rect	125	144	126	145
rect	125	146	126	147
rect	125	147	126	148
rect	125	149	126	150
rect	125	150	126	151
rect	125	152	126	153
rect	125	153	126	154
rect	125	155	126	156
rect	125	156	126	157
rect	125	158	126	159
rect	125	159	126	160
rect	125	161	126	162
rect	125	162	126	163
rect	125	164	126	165
rect	125	165	126	166
rect	125	167	126	168
rect	125	168	126	169
rect	125	170	126	171
rect	125	171	126	172
rect	125	173	126	174
rect	125	174	126	175
rect	125	176	126	177
rect	125	177	126	178
rect	125	179	126	180
rect	125	180	126	181
rect	125	182	126	183
rect	125	183	126	184
rect	125	185	126	186
rect	125	186	126	187
rect	125	188	126	189
rect	125	189	126	190
rect	125	191	126	192
rect	125	192	126	193
rect	125	194	126	195
rect	125	195	126	196
rect	125	197	126	198
rect	125	198	126	199
rect	125	200	126	201
rect	125	201	126	202
rect	125	203	126	204
rect	125	204	126	205
rect	125	206	126	207
rect	125	207	126	208
rect	125	209	126	210
rect	125	210	126	211
rect	125	212	126	213
rect	125	213	126	214
rect	125	215	126	216
rect	125	216	126	217
rect	125	218	126	219
rect	125	219	126	220
rect	125	221	126	222
rect	125	222	126	223
rect	125	224	126	225
rect	125	225	126	226
rect	125	227	126	228
rect	125	228	126	229
rect	125	230	126	231
rect	125	231	126	232
rect	125	233	126	234
rect	125	234	126	235
rect	125	236	126	237
rect	125	237	126	238
rect	125	239	126	240
rect	125	240	126	241
rect	125	242	126	243
rect	125	243	126	244
rect	125	245	126	246
rect	125	246	126	247
rect	125	248	126	249
rect	125	249	126	250
rect	125	251	126	252
rect	125	252	126	253
rect	125	254	126	255
rect	125	255	126	256
rect	125	257	126	258
rect	125	258	126	259
rect	125	260	126	261
rect	125	261	126	262
rect	125	263	126	264
rect	125	264	126	265
rect	125	266	126	267
rect	125	267	126	268
rect	125	269	126	270
rect	125	270	126	271
rect	125	272	126	273
rect	125	273	126	274
rect	125	275	126	276
rect	125	276	126	277
rect	125	278	126	279
rect	125	279	126	280
rect	125	281	126	282
rect	125	282	126	283
rect	125	284	126	285
rect	125	285	126	286
rect	125	287	126	288
rect	125	288	126	289
rect	125	290	126	291
rect	125	291	126	292
rect	125	293	126	294
rect	125	294	126	295
rect	125	296	126	297
rect	125	297	126	298
rect	125	299	126	300
rect	125	300	126	301
rect	125	302	126	303
rect	125	303	126	304
rect	125	305	126	306
rect	125	306	126	307
rect	125	308	126	309
rect	125	309	126	310
rect	125	311	126	312
rect	125	312	126	313
rect	125	314	126	315
rect	125	315	126	316
rect	125	317	126	318
rect	125	318	126	319
rect	125	320	126	321
rect	125	321	126	322
rect	125	323	126	324
rect	125	324	126	325
rect	125	326	126	327
rect	125	327	126	328
rect	125	329	126	330
rect	125	330	126	331
rect	125	332	126	333
rect	125	333	126	334
rect	125	335	126	336
rect	125	336	126	337
rect	125	338	126	339
rect	125	339	126	340
rect	125	341	126	342
rect	125	342	126	343
rect	125	344	126	345
rect	125	345	126	346
rect	125	347	126	348
rect	125	348	126	349
rect	125	350	126	351
rect	125	351	126	352
rect	125	353	126	354
rect	125	354	126	355
rect	125	356	126	357
rect	125	357	126	358
rect	125	359	126	360
rect	125	360	126	361
rect	125	362	126	363
rect	125	363	126	364
rect	125	365	126	366
rect	130	0	131	1
rect	130	2	131	3
rect	130	3	131	4
rect	130	5	131	6
rect	130	6	131	7
rect	130	8	131	9
rect	130	9	131	10
rect	130	11	131	12
rect	130	12	131	13
rect	130	14	131	15
rect	130	15	131	16
rect	130	17	131	18
rect	130	18	131	19
rect	130	20	131	21
rect	130	21	131	22
rect	130	23	131	24
rect	130	24	131	25
rect	130	26	131	27
rect	130	27	131	28
rect	130	29	131	30
rect	130	30	131	31
rect	130	32	131	33
rect	130	33	131	34
rect	130	35	131	36
rect	130	36	131	37
rect	130	38	131	39
rect	130	39	131	40
rect	130	41	131	42
rect	130	42	131	43
rect	130	44	131	45
rect	130	45	131	46
rect	130	47	131	48
rect	130	48	131	49
rect	130	50	131	51
rect	130	51	131	52
rect	130	53	131	54
rect	130	54	131	55
rect	130	56	131	57
rect	130	57	131	58
rect	130	59	131	60
rect	130	60	131	61
rect	130	62	131	63
rect	130	63	131	64
rect	130	65	131	66
rect	130	66	131	67
rect	130	68	131	69
rect	130	69	131	70
rect	130	71	131	72
rect	130	72	131	73
rect	130	74	131	75
rect	130	75	131	76
rect	130	77	131	78
rect	130	78	131	79
rect	130	80	131	81
rect	130	81	131	82
rect	130	83	131	84
rect	130	84	131	85
rect	130	86	131	87
rect	130	87	131	88
rect	130	89	131	90
rect	130	90	131	91
rect	130	92	131	93
rect	130	93	131	94
rect	130	95	131	96
rect	130	96	131	97
rect	130	98	131	99
rect	130	99	131	100
rect	130	101	131	102
rect	130	102	131	103
rect	130	104	131	105
rect	130	105	131	106
rect	130	107	131	108
rect	130	108	131	109
rect	130	110	131	111
rect	130	111	131	112
rect	130	113	131	114
rect	130	114	131	115
rect	130	116	131	117
rect	130	117	131	118
rect	130	119	131	120
rect	130	120	131	121
rect	130	122	131	123
rect	130	123	131	124
rect	130	125	131	126
rect	130	126	131	127
rect	130	128	131	129
rect	130	129	131	130
rect	130	131	131	132
rect	130	132	131	133
rect	130	134	131	135
rect	130	135	131	136
rect	130	137	131	138
rect	130	138	131	139
rect	130	140	131	141
rect	130	141	131	142
rect	130	143	131	144
rect	130	144	131	145
rect	130	146	131	147
rect	130	147	131	148
rect	130	149	131	150
rect	130	150	131	151
rect	130	152	131	153
rect	130	153	131	154
rect	130	155	131	156
rect	130	156	131	157
rect	130	158	131	159
rect	130	159	131	160
rect	130	161	131	162
rect	130	162	131	163
rect	130	164	131	165
rect	130	165	131	166
rect	130	167	131	168
rect	130	168	131	169
rect	130	170	131	171
rect	130	171	131	172
rect	130	173	131	174
rect	130	174	131	175
rect	130	176	131	177
rect	130	177	131	178
rect	130	179	131	180
rect	130	180	131	181
rect	130	182	131	183
rect	130	183	131	184
rect	130	185	131	186
rect	130	186	131	187
rect	130	188	131	189
rect	130	189	131	190
rect	130	191	131	192
rect	130	192	131	193
rect	130	194	131	195
rect	130	195	131	196
rect	130	197	131	198
rect	130	198	131	199
rect	130	200	131	201
rect	130	201	131	202
rect	130	203	131	204
rect	130	204	131	205
rect	130	206	131	207
rect	130	207	131	208
rect	130	209	131	210
rect	130	210	131	211
rect	130	212	131	213
rect	130	213	131	214
rect	130	215	131	216
rect	130	216	131	217
rect	130	218	131	219
rect	130	219	131	220
rect	130	221	131	222
rect	130	222	131	223
rect	130	224	131	225
rect	130	225	131	226
rect	130	227	131	228
rect	130	228	131	229
rect	130	230	131	231
rect	130	231	131	232
rect	130	233	131	234
rect	130	234	131	235
rect	130	236	131	237
rect	130	237	131	238
rect	130	239	131	240
rect	130	240	131	241
rect	130	242	131	243
rect	130	243	131	244
rect	130	245	131	246
rect	130	246	131	247
rect	130	248	131	249
rect	130	249	131	250
rect	130	251	131	252
rect	130	252	131	253
rect	130	254	131	255
rect	130	255	131	256
rect	130	257	131	258
rect	130	258	131	259
rect	130	260	131	261
rect	130	261	131	262
rect	130	263	131	264
rect	130	264	131	265
rect	130	266	131	267
rect	130	267	131	268
rect	130	269	131	270
rect	130	270	131	271
rect	130	272	131	273
rect	130	273	131	274
rect	130	275	131	276
rect	130	276	131	277
rect	130	278	131	279
rect	130	279	131	280
rect	130	281	131	282
rect	130	282	131	283
rect	130	284	131	285
rect	130	285	131	286
rect	130	287	131	288
rect	130	288	131	289
rect	130	290	131	291
rect	130	291	131	292
rect	130	293	131	294
rect	130	294	131	295
rect	130	296	131	297
rect	130	297	131	298
rect	130	299	131	300
rect	130	300	131	301
rect	130	302	131	303
rect	130	303	131	304
rect	130	305	131	306
rect	130	306	131	307
rect	130	308	131	309
rect	130	309	131	310
rect	130	311	131	312
rect	130	312	131	313
rect	130	314	131	315
rect	130	315	131	316
rect	130	317	131	318
rect	130	318	131	319
rect	130	320	131	321
rect	130	321	131	322
rect	130	323	131	324
rect	130	324	131	325
rect	130	326	131	327
rect	130	327	131	328
rect	130	329	131	330
rect	130	330	131	331
rect	130	332	131	333
rect	130	333	131	334
rect	130	335	131	336
rect	130	336	131	337
rect	130	337	131	338
rect	130	338	131	339
rect	130	339	131	340
rect	130	341	131	342
rect	130	342	131	343
rect	130	344	131	345
rect	130	345	131	346
rect	130	347	131	348
rect	130	348	131	349
rect	130	350	131	351
rect	130	351	131	352
rect	130	353	131	354
rect	130	354	131	355
rect	130	356	131	357
rect	130	357	131	358
rect	130	359	131	360
rect	130	360	131	361
rect	130	362	131	363
rect	130	363	131	364
rect	130	365	131	366
rect	132	0	133	1
rect	132	2	133	3
rect	132	3	133	4
rect	132	5	133	6
rect	132	6	133	7
rect	132	8	133	9
rect	132	9	133	10
rect	132	11	133	12
rect	132	12	133	13
rect	132	14	133	15
rect	132	15	133	16
rect	132	17	133	18
rect	132	18	133	19
rect	132	20	133	21
rect	132	21	133	22
rect	132	23	133	24
rect	132	24	133	25
rect	132	26	133	27
rect	132	27	133	28
rect	132	29	133	30
rect	132	30	133	31
rect	132	32	133	33
rect	132	33	133	34
rect	132	35	133	36
rect	132	36	133	37
rect	132	38	133	39
rect	132	39	133	40
rect	132	41	133	42
rect	132	42	133	43
rect	132	44	133	45
rect	132	45	133	46
rect	132	47	133	48
rect	132	48	133	49
rect	132	50	133	51
rect	132	51	133	52
rect	132	53	133	54
rect	132	54	133	55
rect	132	56	133	57
rect	132	57	133	58
rect	132	59	133	60
rect	132	60	133	61
rect	132	62	133	63
rect	132	63	133	64
rect	132	65	133	66
rect	132	66	133	67
rect	132	68	133	69
rect	132	69	133	70
rect	132	71	133	72
rect	132	72	133	73
rect	132	74	133	75
rect	132	75	133	76
rect	132	77	133	78
rect	132	78	133	79
rect	132	80	133	81
rect	132	81	133	82
rect	132	83	133	84
rect	132	84	133	85
rect	132	86	133	87
rect	132	87	133	88
rect	132	89	133	90
rect	132	90	133	91
rect	132	92	133	93
rect	132	93	133	94
rect	132	95	133	96
rect	132	96	133	97
rect	132	98	133	99
rect	132	99	133	100
rect	132	101	133	102
rect	132	102	133	103
rect	132	104	133	105
rect	132	105	133	106
rect	132	107	133	108
rect	132	108	133	109
rect	132	110	133	111
rect	132	111	133	112
rect	132	113	133	114
rect	132	114	133	115
rect	132	116	133	117
rect	132	117	133	118
rect	132	119	133	120
rect	132	120	133	121
rect	132	122	133	123
rect	132	123	133	124
rect	132	125	133	126
rect	132	126	133	127
rect	132	128	133	129
rect	132	129	133	130
rect	132	131	133	132
rect	132	132	133	133
rect	132	134	133	135
rect	132	135	133	136
rect	132	137	133	138
rect	132	138	133	139
rect	132	140	133	141
rect	132	141	133	142
rect	132	143	133	144
rect	132	144	133	145
rect	132	146	133	147
rect	132	147	133	148
rect	132	149	133	150
rect	132	150	133	151
rect	132	152	133	153
rect	132	153	133	154
rect	132	155	133	156
rect	132	156	133	157
rect	132	158	133	159
rect	132	159	133	160
rect	132	161	133	162
rect	132	162	133	163
rect	132	164	133	165
rect	132	165	133	166
rect	132	167	133	168
rect	132	168	133	169
rect	132	170	133	171
rect	132	171	133	172
rect	132	173	133	174
rect	132	174	133	175
rect	132	176	133	177
rect	132	177	133	178
rect	132	179	133	180
rect	132	180	133	181
rect	132	182	133	183
rect	132	183	133	184
rect	132	185	133	186
rect	132	186	133	187
rect	132	188	133	189
rect	132	189	133	190
rect	132	191	133	192
rect	132	192	133	193
rect	132	194	133	195
rect	132	195	133	196
rect	132	197	133	198
rect	132	198	133	199
rect	132	200	133	201
rect	132	201	133	202
rect	132	203	133	204
rect	132	204	133	205
rect	132	206	133	207
rect	132	207	133	208
rect	132	209	133	210
rect	132	210	133	211
rect	132	212	133	213
rect	132	213	133	214
rect	132	215	133	216
rect	132	216	133	217
rect	132	218	133	219
rect	132	219	133	220
rect	132	221	133	222
rect	132	222	133	223
rect	132	224	133	225
rect	132	225	133	226
rect	132	227	133	228
rect	132	228	133	229
rect	132	230	133	231
rect	132	231	133	232
rect	132	233	133	234
rect	132	234	133	235
rect	132	236	133	237
rect	132	237	133	238
rect	132	239	133	240
rect	132	240	133	241
rect	132	242	133	243
rect	132	243	133	244
rect	132	245	133	246
rect	132	246	133	247
rect	132	248	133	249
rect	132	249	133	250
rect	132	251	133	252
rect	132	252	133	253
rect	132	254	133	255
rect	132	255	133	256
rect	132	257	133	258
rect	132	258	133	259
rect	132	260	133	261
rect	132	261	133	262
rect	132	263	133	264
rect	132	264	133	265
rect	132	266	133	267
rect	132	267	133	268
rect	132	269	133	270
rect	132	270	133	271
rect	132	272	133	273
rect	132	273	133	274
rect	132	275	133	276
rect	132	276	133	277
rect	132	278	133	279
rect	132	279	133	280
rect	132	281	133	282
rect	132	282	133	283
rect	132	284	133	285
rect	132	285	133	286
rect	132	287	133	288
rect	132	288	133	289
rect	132	290	133	291
rect	132	291	133	292
rect	132	293	133	294
rect	132	294	133	295
rect	132	296	133	297
rect	132	297	133	298
rect	132	299	133	300
rect	132	300	133	301
rect	132	302	133	303
rect	132	303	133	304
rect	132	305	133	306
rect	132	306	133	307
rect	132	308	133	309
rect	132	309	133	310
rect	132	311	133	312
rect	132	312	133	313
rect	132	314	133	315
rect	132	315	133	316
rect	132	317	133	318
rect	132	318	133	319
rect	132	320	133	321
rect	132	321	133	322
rect	132	323	133	324
rect	132	324	133	325
rect	132	326	133	327
rect	132	327	133	328
rect	132	329	133	330
rect	132	330	133	331
rect	132	332	133	333
rect	132	333	133	334
rect	132	335	133	336
rect	132	336	133	337
rect	132	337	133	338
rect	132	338	133	339
rect	132	339	133	340
rect	132	341	133	342
rect	132	342	133	343
rect	132	344	133	345
rect	132	345	133	346
rect	132	347	133	348
rect	132	348	133	349
rect	132	350	133	351
rect	132	351	133	352
rect	132	353	133	354
rect	132	354	133	355
rect	132	356	133	357
rect	132	357	133	358
rect	132	359	133	360
rect	132	360	133	361
rect	132	362	133	363
rect	132	363	133	364
rect	132	365	133	366
rect	133	0	134	1
rect	133	2	134	3
rect	133	3	134	4
rect	133	5	134	6
rect	133	6	134	7
rect	133	8	134	9
rect	133	9	134	10
rect	133	11	134	12
rect	133	12	134	13
rect	133	14	134	15
rect	133	15	134	16
rect	133	17	134	18
rect	133	18	134	19
rect	133	20	134	21
rect	133	21	134	22
rect	133	23	134	24
rect	133	24	134	25
rect	133	26	134	27
rect	133	27	134	28
rect	133	29	134	30
rect	133	30	134	31
rect	133	32	134	33
rect	133	33	134	34
rect	133	35	134	36
rect	133	36	134	37
rect	133	38	134	39
rect	133	39	134	40
rect	133	41	134	42
rect	133	42	134	43
rect	133	44	134	45
rect	133	45	134	46
rect	133	47	134	48
rect	133	48	134	49
rect	133	50	134	51
rect	133	51	134	52
rect	133	53	134	54
rect	133	54	134	55
rect	133	56	134	57
rect	133	57	134	58
rect	133	59	134	60
rect	133	60	134	61
rect	133	62	134	63
rect	133	63	134	64
rect	133	65	134	66
rect	133	66	134	67
rect	133	68	134	69
rect	133	69	134	70
rect	133	71	134	72
rect	133	72	134	73
rect	133	74	134	75
rect	133	75	134	76
rect	133	77	134	78
rect	133	78	134	79
rect	133	80	134	81
rect	133	81	134	82
rect	133	83	134	84
rect	133	84	134	85
rect	133	86	134	87
rect	133	87	134	88
rect	133	89	134	90
rect	133	90	134	91
rect	133	92	134	93
rect	133	93	134	94
rect	133	95	134	96
rect	133	96	134	97
rect	133	98	134	99
rect	133	99	134	100
rect	133	101	134	102
rect	133	102	134	103
rect	133	104	134	105
rect	133	105	134	106
rect	133	107	134	108
rect	133	108	134	109
rect	133	110	134	111
rect	133	111	134	112
rect	133	113	134	114
rect	133	114	134	115
rect	133	116	134	117
rect	133	117	134	118
rect	133	119	134	120
rect	133	120	134	121
rect	133	122	134	123
rect	133	123	134	124
rect	133	125	134	126
rect	133	126	134	127
rect	133	128	134	129
rect	133	129	134	130
rect	133	131	134	132
rect	133	132	134	133
rect	133	134	134	135
rect	133	135	134	136
rect	133	137	134	138
rect	133	138	134	139
rect	133	140	134	141
rect	133	141	134	142
rect	133	143	134	144
rect	133	144	134	145
rect	133	146	134	147
rect	133	147	134	148
rect	133	149	134	150
rect	133	150	134	151
rect	133	152	134	153
rect	133	153	134	154
rect	133	155	134	156
rect	133	156	134	157
rect	133	158	134	159
rect	133	159	134	160
rect	133	161	134	162
rect	133	162	134	163
rect	133	164	134	165
rect	133	165	134	166
rect	133	167	134	168
rect	133	168	134	169
rect	133	170	134	171
rect	133	171	134	172
rect	133	173	134	174
rect	133	174	134	175
rect	133	176	134	177
rect	133	177	134	178
rect	133	179	134	180
rect	133	180	134	181
rect	133	182	134	183
rect	133	183	134	184
rect	133	185	134	186
rect	133	186	134	187
rect	133	188	134	189
rect	133	189	134	190
rect	133	191	134	192
rect	133	192	134	193
rect	133	194	134	195
rect	133	195	134	196
rect	133	197	134	198
rect	133	198	134	199
rect	133	200	134	201
rect	133	201	134	202
rect	133	203	134	204
rect	133	204	134	205
rect	133	206	134	207
rect	133	207	134	208
rect	133	209	134	210
rect	133	210	134	211
rect	133	212	134	213
rect	133	213	134	214
rect	133	215	134	216
rect	133	216	134	217
rect	133	218	134	219
rect	133	219	134	220
rect	133	221	134	222
rect	133	222	134	223
rect	133	224	134	225
rect	133	225	134	226
rect	133	227	134	228
rect	133	228	134	229
rect	133	230	134	231
rect	133	231	134	232
rect	133	233	134	234
rect	133	234	134	235
rect	133	236	134	237
rect	133	237	134	238
rect	133	239	134	240
rect	133	240	134	241
rect	133	242	134	243
rect	133	243	134	244
rect	133	245	134	246
rect	133	246	134	247
rect	133	248	134	249
rect	133	249	134	250
rect	133	251	134	252
rect	133	252	134	253
rect	133	254	134	255
rect	133	255	134	256
rect	133	257	134	258
rect	133	258	134	259
rect	133	260	134	261
rect	133	261	134	262
rect	133	263	134	264
rect	133	264	134	265
rect	133	266	134	267
rect	133	267	134	268
rect	133	269	134	270
rect	133	270	134	271
rect	133	272	134	273
rect	133	273	134	274
rect	133	275	134	276
rect	133	276	134	277
rect	133	278	134	279
rect	133	279	134	280
rect	133	281	134	282
rect	133	282	134	283
rect	133	284	134	285
rect	133	285	134	286
rect	133	287	134	288
rect	133	288	134	289
rect	133	290	134	291
rect	133	291	134	292
rect	133	293	134	294
rect	133	294	134	295
rect	133	296	134	297
rect	133	297	134	298
rect	133	299	134	300
rect	133	300	134	301
rect	133	302	134	303
rect	133	303	134	304
rect	133	305	134	306
rect	133	306	134	307
rect	133	308	134	309
rect	133	309	134	310
rect	133	311	134	312
rect	133	312	134	313
rect	133	314	134	315
rect	133	315	134	316
rect	133	317	134	318
rect	133	318	134	319
rect	133	320	134	321
rect	133	321	134	322
rect	133	323	134	324
rect	133	324	134	325
rect	133	326	134	327
rect	133	327	134	328
rect	133	329	134	330
rect	133	330	134	331
rect	133	332	134	333
rect	133	333	134	334
rect	133	335	134	336
rect	133	336	134	337
rect	133	337	134	338
rect	133	338	134	339
rect	133	339	134	340
rect	133	341	134	342
rect	133	342	134	343
rect	133	344	134	345
rect	133	345	134	346
rect	133	347	134	348
rect	133	348	134	349
rect	133	350	134	351
rect	133	351	134	352
rect	133	353	134	354
rect	133	354	134	355
rect	133	356	134	357
rect	133	357	134	358
rect	133	359	134	360
rect	133	360	134	361
rect	133	362	134	363
rect	133	363	134	364
rect	133	365	134	366
rect	134	0	135	1
rect	134	2	135	3
rect	134	3	135	4
rect	134	5	135	6
rect	134	6	135	7
rect	134	8	135	9
rect	134	9	135	10
rect	134	11	135	12
rect	134	12	135	13
rect	134	14	135	15
rect	134	15	135	16
rect	134	17	135	18
rect	134	18	135	19
rect	134	20	135	21
rect	134	21	135	22
rect	134	23	135	24
rect	134	24	135	25
rect	134	26	135	27
rect	134	27	135	28
rect	134	29	135	30
rect	134	30	135	31
rect	134	32	135	33
rect	134	33	135	34
rect	134	35	135	36
rect	134	36	135	37
rect	134	38	135	39
rect	134	39	135	40
rect	134	41	135	42
rect	134	42	135	43
rect	134	44	135	45
rect	134	45	135	46
rect	134	47	135	48
rect	134	48	135	49
rect	134	50	135	51
rect	134	51	135	52
rect	134	53	135	54
rect	134	54	135	55
rect	134	56	135	57
rect	134	57	135	58
rect	134	59	135	60
rect	134	60	135	61
rect	134	62	135	63
rect	134	63	135	64
rect	134	65	135	66
rect	134	66	135	67
rect	134	68	135	69
rect	134	69	135	70
rect	134	71	135	72
rect	134	72	135	73
rect	134	74	135	75
rect	134	75	135	76
rect	134	77	135	78
rect	134	78	135	79
rect	134	80	135	81
rect	134	81	135	82
rect	134	83	135	84
rect	134	84	135	85
rect	134	86	135	87
rect	134	87	135	88
rect	134	89	135	90
rect	134	90	135	91
rect	134	92	135	93
rect	134	93	135	94
rect	134	95	135	96
rect	134	96	135	97
rect	134	98	135	99
rect	134	99	135	100
rect	134	101	135	102
rect	134	102	135	103
rect	134	104	135	105
rect	134	105	135	106
rect	134	107	135	108
rect	134	108	135	109
rect	134	110	135	111
rect	134	111	135	112
rect	134	113	135	114
rect	134	114	135	115
rect	134	116	135	117
rect	134	117	135	118
rect	134	119	135	120
rect	134	120	135	121
rect	134	122	135	123
rect	134	123	135	124
rect	134	125	135	126
rect	134	126	135	127
rect	134	128	135	129
rect	134	129	135	130
rect	134	131	135	132
rect	134	132	135	133
rect	134	134	135	135
rect	134	135	135	136
rect	134	137	135	138
rect	134	138	135	139
rect	134	140	135	141
rect	134	141	135	142
rect	134	143	135	144
rect	134	144	135	145
rect	134	146	135	147
rect	134	147	135	148
rect	134	149	135	150
rect	134	150	135	151
rect	134	152	135	153
rect	134	153	135	154
rect	134	155	135	156
rect	134	156	135	157
rect	134	158	135	159
rect	134	159	135	160
rect	134	161	135	162
rect	134	162	135	163
rect	134	164	135	165
rect	134	165	135	166
rect	134	167	135	168
rect	134	168	135	169
rect	134	170	135	171
rect	134	171	135	172
rect	134	173	135	174
rect	134	174	135	175
rect	134	176	135	177
rect	134	177	135	178
rect	134	179	135	180
rect	134	180	135	181
rect	134	182	135	183
rect	134	183	135	184
rect	134	185	135	186
rect	134	186	135	187
rect	134	188	135	189
rect	134	189	135	190
rect	134	191	135	192
rect	134	192	135	193
rect	134	194	135	195
rect	134	195	135	196
rect	134	197	135	198
rect	134	198	135	199
rect	134	200	135	201
rect	134	201	135	202
rect	134	203	135	204
rect	134	204	135	205
rect	134	206	135	207
rect	134	207	135	208
rect	134	209	135	210
rect	134	210	135	211
rect	134	212	135	213
rect	134	213	135	214
rect	134	215	135	216
rect	134	216	135	217
rect	134	218	135	219
rect	134	219	135	220
rect	134	221	135	222
rect	134	222	135	223
rect	134	224	135	225
rect	134	225	135	226
rect	134	227	135	228
rect	134	228	135	229
rect	134	230	135	231
rect	134	231	135	232
rect	134	233	135	234
rect	134	234	135	235
rect	134	236	135	237
rect	134	237	135	238
rect	134	239	135	240
rect	134	240	135	241
rect	134	242	135	243
rect	134	243	135	244
rect	134	245	135	246
rect	134	246	135	247
rect	134	248	135	249
rect	134	249	135	250
rect	134	251	135	252
rect	134	252	135	253
rect	134	254	135	255
rect	134	255	135	256
rect	134	257	135	258
rect	134	258	135	259
rect	134	260	135	261
rect	134	261	135	262
rect	134	263	135	264
rect	134	264	135	265
rect	134	266	135	267
rect	134	267	135	268
rect	134	269	135	270
rect	134	270	135	271
rect	134	272	135	273
rect	134	273	135	274
rect	134	275	135	276
rect	134	276	135	277
rect	134	278	135	279
rect	134	279	135	280
rect	134	281	135	282
rect	134	282	135	283
rect	134	284	135	285
rect	134	285	135	286
rect	134	287	135	288
rect	134	288	135	289
rect	134	290	135	291
rect	134	291	135	292
rect	134	293	135	294
rect	134	294	135	295
rect	134	296	135	297
rect	134	297	135	298
rect	134	299	135	300
rect	134	300	135	301
rect	134	302	135	303
rect	134	303	135	304
rect	134	305	135	306
rect	134	306	135	307
rect	134	308	135	309
rect	134	309	135	310
rect	134	311	135	312
rect	134	312	135	313
rect	134	314	135	315
rect	134	315	135	316
rect	134	317	135	318
rect	134	318	135	319
rect	134	320	135	321
rect	134	321	135	322
rect	134	323	135	324
rect	134	324	135	325
rect	134	326	135	327
rect	134	327	135	328
rect	134	329	135	330
rect	134	330	135	331
rect	134	332	135	333
rect	134	333	135	334
rect	134	335	135	336
rect	134	336	135	337
rect	134	337	135	338
rect	134	338	135	339
rect	134	339	135	340
rect	134	341	135	342
rect	134	342	135	343
rect	134	344	135	345
rect	134	345	135	346
rect	134	347	135	348
rect	134	348	135	349
rect	134	350	135	351
rect	134	351	135	352
rect	134	353	135	354
rect	134	354	135	355
rect	134	356	135	357
rect	134	357	135	358
rect	134	359	135	360
rect	134	360	135	361
rect	134	362	135	363
rect	134	363	135	364
rect	134	365	135	366
rect	135	0	136	1
rect	135	2	136	3
rect	135	3	136	4
rect	135	5	136	6
rect	135	6	136	7
rect	135	8	136	9
rect	135	9	136	10
rect	135	11	136	12
rect	135	12	136	13
rect	135	14	136	15
rect	135	15	136	16
rect	135	17	136	18
rect	135	18	136	19
rect	135	20	136	21
rect	135	21	136	22
rect	135	23	136	24
rect	135	24	136	25
rect	135	26	136	27
rect	135	27	136	28
rect	135	29	136	30
rect	135	30	136	31
rect	135	32	136	33
rect	135	33	136	34
rect	135	35	136	36
rect	135	36	136	37
rect	135	38	136	39
rect	135	39	136	40
rect	135	41	136	42
rect	135	42	136	43
rect	135	44	136	45
rect	135	45	136	46
rect	135	47	136	48
rect	135	48	136	49
rect	135	50	136	51
rect	135	51	136	52
rect	135	53	136	54
rect	135	54	136	55
rect	135	56	136	57
rect	135	57	136	58
rect	135	59	136	60
rect	135	60	136	61
rect	135	62	136	63
rect	135	63	136	64
rect	135	65	136	66
rect	135	66	136	67
rect	135	68	136	69
rect	135	69	136	70
rect	135	71	136	72
rect	135	72	136	73
rect	135	74	136	75
rect	135	75	136	76
rect	135	77	136	78
rect	135	78	136	79
rect	135	80	136	81
rect	135	81	136	82
rect	135	83	136	84
rect	135	84	136	85
rect	135	86	136	87
rect	135	87	136	88
rect	135	89	136	90
rect	135	90	136	91
rect	135	92	136	93
rect	135	93	136	94
rect	135	95	136	96
rect	135	96	136	97
rect	135	98	136	99
rect	135	99	136	100
rect	135	101	136	102
rect	135	102	136	103
rect	135	104	136	105
rect	135	105	136	106
rect	135	107	136	108
rect	135	108	136	109
rect	135	110	136	111
rect	135	111	136	112
rect	135	113	136	114
rect	135	114	136	115
rect	135	116	136	117
rect	135	117	136	118
rect	135	119	136	120
rect	135	120	136	121
rect	135	122	136	123
rect	135	123	136	124
rect	135	125	136	126
rect	135	126	136	127
rect	135	128	136	129
rect	135	129	136	130
rect	135	131	136	132
rect	135	132	136	133
rect	135	134	136	135
rect	135	135	136	136
rect	135	137	136	138
rect	135	138	136	139
rect	135	140	136	141
rect	135	141	136	142
rect	135	143	136	144
rect	135	144	136	145
rect	135	146	136	147
rect	135	147	136	148
rect	135	149	136	150
rect	135	150	136	151
rect	135	152	136	153
rect	135	153	136	154
rect	135	155	136	156
rect	135	156	136	157
rect	135	158	136	159
rect	135	159	136	160
rect	135	161	136	162
rect	135	162	136	163
rect	135	164	136	165
rect	135	165	136	166
rect	135	167	136	168
rect	135	168	136	169
rect	135	170	136	171
rect	135	171	136	172
rect	135	173	136	174
rect	135	174	136	175
rect	135	176	136	177
rect	135	177	136	178
rect	135	179	136	180
rect	135	180	136	181
rect	135	182	136	183
rect	135	183	136	184
rect	135	185	136	186
rect	135	186	136	187
rect	135	188	136	189
rect	135	189	136	190
rect	135	191	136	192
rect	135	192	136	193
rect	135	194	136	195
rect	135	195	136	196
rect	135	197	136	198
rect	135	198	136	199
rect	135	200	136	201
rect	135	201	136	202
rect	135	203	136	204
rect	135	204	136	205
rect	135	206	136	207
rect	135	207	136	208
rect	135	209	136	210
rect	135	210	136	211
rect	135	212	136	213
rect	135	213	136	214
rect	135	215	136	216
rect	135	216	136	217
rect	135	218	136	219
rect	135	219	136	220
rect	135	221	136	222
rect	135	222	136	223
rect	135	224	136	225
rect	135	225	136	226
rect	135	227	136	228
rect	135	228	136	229
rect	135	230	136	231
rect	135	231	136	232
rect	135	233	136	234
rect	135	234	136	235
rect	135	236	136	237
rect	135	237	136	238
rect	135	239	136	240
rect	135	240	136	241
rect	135	242	136	243
rect	135	243	136	244
rect	135	245	136	246
rect	135	246	136	247
rect	135	248	136	249
rect	135	249	136	250
rect	135	251	136	252
rect	135	252	136	253
rect	135	254	136	255
rect	135	255	136	256
rect	135	257	136	258
rect	135	258	136	259
rect	135	260	136	261
rect	135	261	136	262
rect	135	263	136	264
rect	135	264	136	265
rect	135	266	136	267
rect	135	267	136	268
rect	135	269	136	270
rect	135	270	136	271
rect	135	272	136	273
rect	135	273	136	274
rect	135	275	136	276
rect	135	276	136	277
rect	135	278	136	279
rect	135	279	136	280
rect	135	281	136	282
rect	135	282	136	283
rect	135	284	136	285
rect	135	285	136	286
rect	135	287	136	288
rect	135	288	136	289
rect	135	290	136	291
rect	135	291	136	292
rect	135	293	136	294
rect	135	294	136	295
rect	135	296	136	297
rect	135	297	136	298
rect	135	299	136	300
rect	135	300	136	301
rect	135	302	136	303
rect	135	303	136	304
rect	135	305	136	306
rect	135	306	136	307
rect	135	308	136	309
rect	135	309	136	310
rect	135	311	136	312
rect	135	312	136	313
rect	135	314	136	315
rect	135	315	136	316
rect	135	317	136	318
rect	135	318	136	319
rect	135	320	136	321
rect	135	321	136	322
rect	135	323	136	324
rect	135	324	136	325
rect	135	326	136	327
rect	135	327	136	328
rect	135	329	136	330
rect	135	330	136	331
rect	135	332	136	333
rect	135	333	136	334
rect	135	335	136	336
rect	135	336	136	337
rect	135	337	136	338
rect	135	338	136	339
rect	135	339	136	340
rect	135	341	136	342
rect	135	342	136	343
rect	135	344	136	345
rect	135	345	136	346
rect	135	347	136	348
rect	135	348	136	349
rect	135	350	136	351
rect	135	351	136	352
rect	135	353	136	354
rect	135	354	136	355
rect	135	356	136	357
rect	135	357	136	358
rect	135	359	136	360
rect	135	360	136	361
rect	135	362	136	363
rect	135	363	136	364
rect	135	365	136	366
rect	136	0	137	1
rect	136	2	137	3
rect	136	3	137	4
rect	136	5	137	6
rect	136	6	137	7
rect	136	8	137	9
rect	136	9	137	10
rect	136	11	137	12
rect	136	12	137	13
rect	136	14	137	15
rect	136	15	137	16
rect	136	17	137	18
rect	136	18	137	19
rect	136	20	137	21
rect	136	21	137	22
rect	136	23	137	24
rect	136	24	137	25
rect	136	26	137	27
rect	136	27	137	28
rect	136	29	137	30
rect	136	30	137	31
rect	136	32	137	33
rect	136	33	137	34
rect	136	35	137	36
rect	136	36	137	37
rect	136	38	137	39
rect	136	39	137	40
rect	136	41	137	42
rect	136	42	137	43
rect	136	44	137	45
rect	136	45	137	46
rect	136	47	137	48
rect	136	48	137	49
rect	136	50	137	51
rect	136	51	137	52
rect	136	53	137	54
rect	136	54	137	55
rect	136	56	137	57
rect	136	57	137	58
rect	136	59	137	60
rect	136	60	137	61
rect	136	62	137	63
rect	136	63	137	64
rect	136	65	137	66
rect	136	66	137	67
rect	136	68	137	69
rect	136	69	137	70
rect	136	71	137	72
rect	136	72	137	73
rect	136	74	137	75
rect	136	75	137	76
rect	136	77	137	78
rect	136	78	137	79
rect	136	80	137	81
rect	136	81	137	82
rect	136	83	137	84
rect	136	84	137	85
rect	136	86	137	87
rect	136	87	137	88
rect	136	89	137	90
rect	136	90	137	91
rect	136	92	137	93
rect	136	93	137	94
rect	136	95	137	96
rect	136	96	137	97
rect	136	98	137	99
rect	136	99	137	100
rect	136	101	137	102
rect	136	102	137	103
rect	136	104	137	105
rect	136	105	137	106
rect	136	107	137	108
rect	136	108	137	109
rect	136	110	137	111
rect	136	111	137	112
rect	136	113	137	114
rect	136	114	137	115
rect	136	116	137	117
rect	136	117	137	118
rect	136	119	137	120
rect	136	120	137	121
rect	136	122	137	123
rect	136	123	137	124
rect	136	125	137	126
rect	136	126	137	127
rect	136	128	137	129
rect	136	129	137	130
rect	136	131	137	132
rect	136	132	137	133
rect	136	134	137	135
rect	136	135	137	136
rect	136	137	137	138
rect	136	138	137	139
rect	136	140	137	141
rect	136	141	137	142
rect	136	143	137	144
rect	136	144	137	145
rect	136	146	137	147
rect	136	147	137	148
rect	136	149	137	150
rect	136	150	137	151
rect	136	152	137	153
rect	136	153	137	154
rect	136	155	137	156
rect	136	156	137	157
rect	136	158	137	159
rect	136	159	137	160
rect	136	161	137	162
rect	136	162	137	163
rect	136	164	137	165
rect	136	165	137	166
rect	136	167	137	168
rect	136	168	137	169
rect	136	170	137	171
rect	136	171	137	172
rect	136	173	137	174
rect	136	174	137	175
rect	136	176	137	177
rect	136	177	137	178
rect	136	179	137	180
rect	136	180	137	181
rect	136	182	137	183
rect	136	183	137	184
rect	136	185	137	186
rect	136	186	137	187
rect	136	188	137	189
rect	136	189	137	190
rect	136	191	137	192
rect	136	192	137	193
rect	136	194	137	195
rect	136	195	137	196
rect	136	197	137	198
rect	136	198	137	199
rect	136	200	137	201
rect	136	201	137	202
rect	136	203	137	204
rect	136	204	137	205
rect	136	206	137	207
rect	136	207	137	208
rect	136	209	137	210
rect	136	210	137	211
rect	136	212	137	213
rect	136	213	137	214
rect	136	215	137	216
rect	136	216	137	217
rect	136	218	137	219
rect	136	219	137	220
rect	136	221	137	222
rect	136	222	137	223
rect	136	224	137	225
rect	136	225	137	226
rect	136	227	137	228
rect	136	228	137	229
rect	136	230	137	231
rect	136	231	137	232
rect	136	233	137	234
rect	136	234	137	235
rect	136	236	137	237
rect	136	237	137	238
rect	136	239	137	240
rect	136	240	137	241
rect	136	242	137	243
rect	136	243	137	244
rect	136	245	137	246
rect	136	246	137	247
rect	136	248	137	249
rect	136	249	137	250
rect	136	251	137	252
rect	136	252	137	253
rect	136	254	137	255
rect	136	255	137	256
rect	136	257	137	258
rect	136	258	137	259
rect	136	260	137	261
rect	136	261	137	262
rect	136	263	137	264
rect	136	264	137	265
rect	136	266	137	267
rect	136	267	137	268
rect	136	269	137	270
rect	136	270	137	271
rect	136	272	137	273
rect	136	273	137	274
rect	136	275	137	276
rect	136	276	137	277
rect	136	278	137	279
rect	136	279	137	280
rect	136	281	137	282
rect	136	282	137	283
rect	136	284	137	285
rect	136	285	137	286
rect	136	287	137	288
rect	136	288	137	289
rect	136	290	137	291
rect	136	291	137	292
rect	136	293	137	294
rect	136	294	137	295
rect	136	296	137	297
rect	136	297	137	298
rect	136	299	137	300
rect	136	300	137	301
rect	136	302	137	303
rect	136	303	137	304
rect	136	305	137	306
rect	136	306	137	307
rect	136	308	137	309
rect	136	309	137	310
rect	136	311	137	312
rect	136	312	137	313
rect	136	314	137	315
rect	136	315	137	316
rect	136	317	137	318
rect	136	318	137	319
rect	136	320	137	321
rect	136	321	137	322
rect	136	323	137	324
rect	136	324	137	325
rect	136	326	137	327
rect	136	327	137	328
rect	136	329	137	330
rect	136	330	137	331
rect	136	332	137	333
rect	136	333	137	334
rect	136	335	137	336
rect	136	336	137	337
rect	136	337	137	338
rect	136	338	137	339
rect	136	339	137	340
rect	136	341	137	342
rect	136	342	137	343
rect	136	344	137	345
rect	136	345	137	346
rect	136	347	137	348
rect	136	348	137	349
rect	136	350	137	351
rect	136	351	137	352
rect	136	353	137	354
rect	136	354	137	355
rect	136	356	137	357
rect	136	357	137	358
rect	136	359	137	360
rect	136	360	137	361
rect	136	362	137	363
rect	136	363	137	364
rect	136	365	137	366
rect	143	0	144	1
rect	143	2	144	3
rect	143	3	144	4
rect	143	5	144	6
rect	143	6	144	7
rect	143	8	144	9
rect	143	9	144	10
rect	143	11	144	12
rect	143	12	144	13
rect	143	14	144	15
rect	143	15	144	16
rect	143	17	144	18
rect	143	18	144	19
rect	143	20	144	21
rect	143	21	144	22
rect	143	23	144	24
rect	143	24	144	25
rect	143	26	144	27
rect	143	27	144	28
rect	143	29	144	30
rect	143	30	144	31
rect	143	32	144	33
rect	143	33	144	34
rect	143	35	144	36
rect	143	36	144	37
rect	143	38	144	39
rect	143	39	144	40
rect	143	41	144	42
rect	143	42	144	43
rect	143	44	144	45
rect	143	45	144	46
rect	143	47	144	48
rect	143	48	144	49
rect	143	50	144	51
rect	143	51	144	52
rect	143	53	144	54
rect	143	54	144	55
rect	143	56	144	57
rect	143	57	144	58
rect	143	59	144	60
rect	143	60	144	61
rect	143	62	144	63
rect	143	63	144	64
rect	143	65	144	66
rect	143	66	144	67
rect	143	68	144	69
rect	143	69	144	70
rect	143	71	144	72
rect	143	72	144	73
rect	143	74	144	75
rect	143	75	144	76
rect	143	77	144	78
rect	143	78	144	79
rect	143	80	144	81
rect	143	81	144	82
rect	143	83	144	84
rect	143	84	144	85
rect	143	86	144	87
rect	143	87	144	88
rect	143	89	144	90
rect	143	90	144	91
rect	143	92	144	93
rect	143	93	144	94
rect	143	95	144	96
rect	143	96	144	97
rect	143	98	144	99
rect	143	99	144	100
rect	143	101	144	102
rect	143	102	144	103
rect	143	104	144	105
rect	143	105	144	106
rect	143	107	144	108
rect	143	108	144	109
rect	143	110	144	111
rect	143	111	144	112
rect	143	113	144	114
rect	143	114	144	115
rect	143	116	144	117
rect	143	117	144	118
rect	143	119	144	120
rect	143	120	144	121
rect	143	122	144	123
rect	143	123	144	124
rect	143	125	144	126
rect	143	126	144	127
rect	143	128	144	129
rect	143	129	144	130
rect	143	131	144	132
rect	143	132	144	133
rect	143	134	144	135
rect	143	135	144	136
rect	143	137	144	138
rect	143	138	144	139
rect	143	140	144	141
rect	143	141	144	142
rect	143	143	144	144
rect	143	144	144	145
rect	143	146	144	147
rect	143	147	144	148
rect	143	149	144	150
rect	143	150	144	151
rect	143	152	144	153
rect	143	153	144	154
rect	143	155	144	156
rect	143	156	144	157
rect	143	158	144	159
rect	143	159	144	160
rect	143	161	144	162
rect	143	162	144	163
rect	143	164	144	165
rect	143	165	144	166
rect	143	167	144	168
rect	143	168	144	169
rect	143	170	144	171
rect	143	171	144	172
rect	143	173	144	174
rect	143	174	144	175
rect	143	176	144	177
rect	143	177	144	178
rect	143	179	144	180
rect	143	180	144	181
rect	143	182	144	183
rect	143	183	144	184
rect	143	185	144	186
rect	143	186	144	187
rect	143	188	144	189
rect	143	189	144	190
rect	143	191	144	192
rect	143	192	144	193
rect	143	194	144	195
rect	143	195	144	196
rect	143	197	144	198
rect	143	198	144	199
rect	143	200	144	201
rect	143	201	144	202
rect	143	203	144	204
rect	143	204	144	205
rect	143	206	144	207
rect	143	207	144	208
rect	143	209	144	210
rect	143	210	144	211
rect	143	212	144	213
rect	143	213	144	214
rect	143	215	144	216
rect	143	216	144	217
rect	143	218	144	219
rect	143	219	144	220
rect	143	221	144	222
rect	143	222	144	223
rect	143	224	144	225
rect	143	225	144	226
rect	143	227	144	228
rect	143	228	144	229
rect	143	230	144	231
rect	143	231	144	232
rect	143	233	144	234
rect	143	234	144	235
rect	143	236	144	237
rect	143	237	144	238
rect	143	239	144	240
rect	143	240	144	241
rect	143	242	144	243
rect	143	243	144	244
rect	143	245	144	246
rect	143	246	144	247
rect	143	248	144	249
rect	143	249	144	250
rect	143	251	144	252
rect	143	252	144	253
rect	143	254	144	255
rect	143	255	144	256
rect	143	257	144	258
rect	143	258	144	259
rect	143	260	144	261
rect	143	261	144	262
rect	143	263	144	264
rect	143	264	144	265
rect	143	266	144	267
rect	143	267	144	268
rect	143	269	144	270
rect	143	270	144	271
rect	143	272	144	273
rect	143	273	144	274
rect	143	275	144	276
rect	143	276	144	277
rect	143	278	144	279
rect	143	279	144	280
rect	143	281	144	282
rect	143	282	144	283
rect	143	284	144	285
rect	143	285	144	286
rect	143	287	144	288
rect	143	288	144	289
rect	143	290	144	291
rect	143	291	144	292
rect	143	293	144	294
rect	143	294	144	295
rect	143	296	144	297
rect	143	297	144	298
rect	143	299	144	300
rect	143	300	144	301
rect	143	302	144	303
rect	143	303	144	304
rect	143	304	144	305
rect	143	305	144	306
rect	143	306	144	307
rect	143	308	144	309
rect	143	309	144	310
rect	143	311	144	312
rect	143	312	144	313
rect	143	314	144	315
rect	143	315	144	316
rect	143	317	144	318
rect	143	318	144	319
rect	143	320	144	321
rect	143	321	144	322
rect	143	323	144	324
rect	143	324	144	325
rect	143	326	144	327
rect	143	327	144	328
rect	143	329	144	330
rect	143	330	144	331
rect	143	332	144	333
rect	143	333	144	334
rect	143	335	144	336
rect	143	336	144	337
rect	143	337	144	338
rect	143	338	144	339
rect	143	339	144	340
rect	143	341	144	342
rect	143	342	144	343
rect	143	344	144	345
rect	143	345	144	346
rect	143	347	144	348
rect	143	348	144	349
rect	143	350	144	351
rect	143	351	144	352
rect	143	353	144	354
rect	143	354	144	355
rect	143	356	144	357
rect	143	357	144	358
rect	143	359	144	360
rect	143	360	144	361
rect	143	362	144	363
rect	143	363	144	364
rect	143	365	144	366
rect	145	0	146	1
rect	145	2	146	3
rect	145	3	146	4
rect	145	5	146	6
rect	145	6	146	7
rect	145	8	146	9
rect	145	9	146	10
rect	145	11	146	12
rect	145	12	146	13
rect	145	14	146	15
rect	145	15	146	16
rect	145	17	146	18
rect	145	18	146	19
rect	145	20	146	21
rect	145	21	146	22
rect	145	23	146	24
rect	145	24	146	25
rect	145	26	146	27
rect	145	27	146	28
rect	145	29	146	30
rect	145	30	146	31
rect	145	32	146	33
rect	145	33	146	34
rect	145	35	146	36
rect	145	36	146	37
rect	145	38	146	39
rect	145	39	146	40
rect	145	41	146	42
rect	145	42	146	43
rect	145	44	146	45
rect	145	45	146	46
rect	145	47	146	48
rect	145	48	146	49
rect	145	50	146	51
rect	145	51	146	52
rect	145	53	146	54
rect	145	54	146	55
rect	145	56	146	57
rect	145	57	146	58
rect	145	59	146	60
rect	145	60	146	61
rect	145	62	146	63
rect	145	63	146	64
rect	145	65	146	66
rect	145	66	146	67
rect	145	68	146	69
rect	145	69	146	70
rect	145	71	146	72
rect	145	72	146	73
rect	145	74	146	75
rect	145	75	146	76
rect	145	77	146	78
rect	145	78	146	79
rect	145	80	146	81
rect	145	81	146	82
rect	145	83	146	84
rect	145	84	146	85
rect	145	86	146	87
rect	145	87	146	88
rect	145	89	146	90
rect	145	90	146	91
rect	145	92	146	93
rect	145	93	146	94
rect	145	95	146	96
rect	145	96	146	97
rect	145	98	146	99
rect	145	99	146	100
rect	145	101	146	102
rect	145	102	146	103
rect	145	104	146	105
rect	145	105	146	106
rect	145	107	146	108
rect	145	108	146	109
rect	145	110	146	111
rect	145	111	146	112
rect	145	113	146	114
rect	145	114	146	115
rect	145	116	146	117
rect	145	117	146	118
rect	145	119	146	120
rect	145	120	146	121
rect	145	122	146	123
rect	145	123	146	124
rect	145	125	146	126
rect	145	126	146	127
rect	145	128	146	129
rect	145	129	146	130
rect	145	131	146	132
rect	145	132	146	133
rect	145	134	146	135
rect	145	135	146	136
rect	145	137	146	138
rect	145	138	146	139
rect	145	140	146	141
rect	145	141	146	142
rect	145	143	146	144
rect	145	144	146	145
rect	145	146	146	147
rect	145	147	146	148
rect	145	149	146	150
rect	145	150	146	151
rect	145	152	146	153
rect	145	153	146	154
rect	145	155	146	156
rect	145	156	146	157
rect	145	158	146	159
rect	145	159	146	160
rect	145	161	146	162
rect	145	162	146	163
rect	145	164	146	165
rect	145	165	146	166
rect	145	167	146	168
rect	145	168	146	169
rect	145	170	146	171
rect	145	171	146	172
rect	145	173	146	174
rect	145	174	146	175
rect	145	176	146	177
rect	145	177	146	178
rect	145	179	146	180
rect	145	180	146	181
rect	145	182	146	183
rect	145	183	146	184
rect	145	185	146	186
rect	145	186	146	187
rect	145	188	146	189
rect	145	189	146	190
rect	145	191	146	192
rect	145	192	146	193
rect	145	194	146	195
rect	145	195	146	196
rect	145	197	146	198
rect	145	198	146	199
rect	145	200	146	201
rect	145	201	146	202
rect	145	203	146	204
rect	145	204	146	205
rect	145	206	146	207
rect	145	207	146	208
rect	145	209	146	210
rect	145	210	146	211
rect	145	212	146	213
rect	145	213	146	214
rect	145	215	146	216
rect	145	216	146	217
rect	145	218	146	219
rect	145	219	146	220
rect	145	221	146	222
rect	145	222	146	223
rect	145	224	146	225
rect	145	225	146	226
rect	145	227	146	228
rect	145	228	146	229
rect	145	230	146	231
rect	145	231	146	232
rect	145	233	146	234
rect	145	234	146	235
rect	145	236	146	237
rect	145	237	146	238
rect	145	239	146	240
rect	145	240	146	241
rect	145	242	146	243
rect	145	243	146	244
rect	145	245	146	246
rect	145	246	146	247
rect	145	248	146	249
rect	145	249	146	250
rect	145	251	146	252
rect	145	252	146	253
rect	145	254	146	255
rect	145	255	146	256
rect	145	257	146	258
rect	145	258	146	259
rect	145	260	146	261
rect	145	261	146	262
rect	145	263	146	264
rect	145	264	146	265
rect	145	266	146	267
rect	145	267	146	268
rect	145	269	146	270
rect	145	270	146	271
rect	145	272	146	273
rect	145	273	146	274
rect	145	275	146	276
rect	145	276	146	277
rect	145	278	146	279
rect	145	279	146	280
rect	145	281	146	282
rect	145	282	146	283
rect	145	284	146	285
rect	145	285	146	286
rect	145	287	146	288
rect	145	288	146	289
rect	145	290	146	291
rect	145	291	146	292
rect	145	293	146	294
rect	145	294	146	295
rect	145	296	146	297
rect	145	297	146	298
rect	145	299	146	300
rect	145	300	146	301
rect	145	302	146	303
rect	145	303	146	304
rect	145	304	146	305
rect	145	305	146	306
rect	145	306	146	307
rect	145	308	146	309
rect	145	309	146	310
rect	145	311	146	312
rect	145	312	146	313
rect	145	314	146	315
rect	145	315	146	316
rect	145	317	146	318
rect	145	318	146	319
rect	145	320	146	321
rect	145	321	146	322
rect	145	323	146	324
rect	145	324	146	325
rect	145	326	146	327
rect	145	327	146	328
rect	145	329	146	330
rect	145	330	146	331
rect	145	332	146	333
rect	145	333	146	334
rect	145	335	146	336
rect	145	336	146	337
rect	145	337	146	338
rect	145	338	146	339
rect	145	339	146	340
rect	145	341	146	342
rect	145	342	146	343
rect	145	344	146	345
rect	145	345	146	346
rect	145	347	146	348
rect	145	348	146	349
rect	145	350	146	351
rect	145	351	146	352
rect	145	353	146	354
rect	145	354	146	355
rect	145	356	146	357
rect	145	357	146	358
rect	145	359	146	360
rect	145	360	146	361
rect	145	362	146	363
rect	145	363	146	364
rect	145	365	146	366
rect	145	366	146	367
rect	145	368	146	369
rect	145	369	146	370
rect	145	370	146	371
rect	145	371	146	372
rect	145	372	146	373
rect	145	374	146	375
rect	145	375	146	376
rect	145	377	146	378
rect	145	378	146	379
rect	145	380	146	381
rect	145	381	146	382
rect	145	382	146	383
rect	145	383	146	384
rect	145	384	146	385
rect	145	386	146	387
rect	146	0	147	1
rect	146	2	147	3
rect	146	3	147	4
rect	146	5	147	6
rect	146	6	147	7
rect	146	8	147	9
rect	146	9	147	10
rect	146	11	147	12
rect	146	12	147	13
rect	146	14	147	15
rect	146	15	147	16
rect	146	17	147	18
rect	146	18	147	19
rect	146	20	147	21
rect	146	21	147	22
rect	146	23	147	24
rect	146	24	147	25
rect	146	26	147	27
rect	146	27	147	28
rect	146	29	147	30
rect	146	30	147	31
rect	146	32	147	33
rect	146	33	147	34
rect	146	35	147	36
rect	146	36	147	37
rect	146	38	147	39
rect	146	39	147	40
rect	146	41	147	42
rect	146	42	147	43
rect	146	44	147	45
rect	146	45	147	46
rect	146	47	147	48
rect	146	48	147	49
rect	146	50	147	51
rect	146	51	147	52
rect	146	53	147	54
rect	146	54	147	55
rect	146	56	147	57
rect	146	57	147	58
rect	146	59	147	60
rect	146	60	147	61
rect	146	62	147	63
rect	146	63	147	64
rect	146	65	147	66
rect	146	66	147	67
rect	146	68	147	69
rect	146	69	147	70
rect	146	71	147	72
rect	146	72	147	73
rect	146	74	147	75
rect	146	75	147	76
rect	146	77	147	78
rect	146	78	147	79
rect	146	80	147	81
rect	146	81	147	82
rect	146	83	147	84
rect	146	84	147	85
rect	146	86	147	87
rect	146	87	147	88
rect	146	89	147	90
rect	146	90	147	91
rect	146	92	147	93
rect	146	93	147	94
rect	146	95	147	96
rect	146	96	147	97
rect	146	98	147	99
rect	146	99	147	100
rect	146	101	147	102
rect	146	102	147	103
rect	146	104	147	105
rect	146	105	147	106
rect	146	107	147	108
rect	146	108	147	109
rect	146	110	147	111
rect	146	111	147	112
rect	146	113	147	114
rect	146	114	147	115
rect	146	116	147	117
rect	146	117	147	118
rect	146	119	147	120
rect	146	120	147	121
rect	146	122	147	123
rect	146	123	147	124
rect	146	125	147	126
rect	146	126	147	127
rect	146	128	147	129
rect	146	129	147	130
rect	146	131	147	132
rect	146	132	147	133
rect	146	134	147	135
rect	146	135	147	136
rect	146	137	147	138
rect	146	138	147	139
rect	146	140	147	141
rect	146	141	147	142
rect	146	143	147	144
rect	146	144	147	145
rect	146	146	147	147
rect	146	147	147	148
rect	146	149	147	150
rect	146	150	147	151
rect	146	152	147	153
rect	146	153	147	154
rect	146	155	147	156
rect	146	156	147	157
rect	146	158	147	159
rect	146	159	147	160
rect	146	161	147	162
rect	146	162	147	163
rect	146	164	147	165
rect	146	165	147	166
rect	146	167	147	168
rect	146	168	147	169
rect	146	170	147	171
rect	146	171	147	172
rect	146	173	147	174
rect	146	174	147	175
rect	146	176	147	177
rect	146	177	147	178
rect	146	179	147	180
rect	146	180	147	181
rect	146	182	147	183
rect	146	183	147	184
rect	146	185	147	186
rect	146	186	147	187
rect	146	188	147	189
rect	146	189	147	190
rect	146	191	147	192
rect	146	192	147	193
rect	146	194	147	195
rect	146	195	147	196
rect	146	197	147	198
rect	146	198	147	199
rect	146	200	147	201
rect	146	201	147	202
rect	146	203	147	204
rect	146	204	147	205
rect	146	206	147	207
rect	146	207	147	208
rect	146	209	147	210
rect	146	210	147	211
rect	146	212	147	213
rect	146	213	147	214
rect	146	215	147	216
rect	146	216	147	217
rect	146	218	147	219
rect	146	219	147	220
rect	146	221	147	222
rect	146	222	147	223
rect	146	224	147	225
rect	146	225	147	226
rect	146	227	147	228
rect	146	228	147	229
rect	146	230	147	231
rect	146	231	147	232
rect	146	233	147	234
rect	146	234	147	235
rect	146	236	147	237
rect	146	237	147	238
rect	146	239	147	240
rect	146	240	147	241
rect	146	242	147	243
rect	146	243	147	244
rect	146	245	147	246
rect	146	246	147	247
rect	146	248	147	249
rect	146	249	147	250
rect	146	251	147	252
rect	146	252	147	253
rect	146	254	147	255
rect	146	255	147	256
rect	146	257	147	258
rect	146	258	147	259
rect	146	260	147	261
rect	146	261	147	262
rect	146	263	147	264
rect	146	264	147	265
rect	146	266	147	267
rect	146	267	147	268
rect	146	269	147	270
rect	146	270	147	271
rect	146	272	147	273
rect	146	273	147	274
rect	146	275	147	276
rect	146	276	147	277
rect	146	278	147	279
rect	146	279	147	280
rect	146	281	147	282
rect	146	282	147	283
rect	146	284	147	285
rect	146	285	147	286
rect	146	287	147	288
rect	146	288	147	289
rect	146	290	147	291
rect	146	291	147	292
rect	146	293	147	294
rect	146	294	147	295
rect	146	296	147	297
rect	146	297	147	298
rect	146	299	147	300
rect	146	300	147	301
rect	146	302	147	303
rect	146	303	147	304
rect	146	304	147	305
rect	146	305	147	306
rect	146	306	147	307
rect	146	308	147	309
rect	146	309	147	310
rect	146	311	147	312
rect	146	312	147	313
rect	146	314	147	315
rect	146	315	147	316
rect	146	317	147	318
rect	146	318	147	319
rect	146	320	147	321
rect	146	321	147	322
rect	146	323	147	324
rect	146	324	147	325
rect	146	326	147	327
rect	146	327	147	328
rect	146	329	147	330
rect	146	330	147	331
rect	146	332	147	333
rect	146	333	147	334
rect	146	335	147	336
rect	146	336	147	337
rect	146	337	147	338
rect	146	338	147	339
rect	146	339	147	340
rect	146	341	147	342
rect	146	342	147	343
rect	146	344	147	345
rect	146	345	147	346
rect	146	347	147	348
rect	146	348	147	349
rect	146	350	147	351
rect	146	351	147	352
rect	146	353	147	354
rect	146	354	147	355
rect	146	356	147	357
rect	146	357	147	358
rect	146	359	147	360
rect	146	360	147	361
rect	146	362	147	363
rect	146	363	147	364
rect	146	365	147	366
rect	146	366	147	367
rect	146	368	147	369
rect	146	369	147	370
rect	146	370	147	371
rect	146	371	147	372
rect	146	372	147	373
rect	146	374	147	375
rect	146	375	147	376
rect	146	377	147	378
rect	146	378	147	379
rect	146	380	147	381
rect	146	381	147	382
rect	146	382	147	383
rect	146	383	147	384
rect	146	384	147	385
rect	146	386	147	387
rect	147	0	148	1
rect	147	2	148	3
rect	147	3	148	4
rect	147	5	148	6
rect	147	6	148	7
rect	147	8	148	9
rect	147	9	148	10
rect	147	11	148	12
rect	147	12	148	13
rect	147	14	148	15
rect	147	15	148	16
rect	147	17	148	18
rect	147	18	148	19
rect	147	20	148	21
rect	147	21	148	22
rect	147	23	148	24
rect	147	24	148	25
rect	147	26	148	27
rect	147	27	148	28
rect	147	29	148	30
rect	147	30	148	31
rect	147	32	148	33
rect	147	33	148	34
rect	147	35	148	36
rect	147	36	148	37
rect	147	38	148	39
rect	147	39	148	40
rect	147	41	148	42
rect	147	42	148	43
rect	147	44	148	45
rect	147	45	148	46
rect	147	47	148	48
rect	147	48	148	49
rect	147	50	148	51
rect	147	51	148	52
rect	147	53	148	54
rect	147	54	148	55
rect	147	56	148	57
rect	147	57	148	58
rect	147	59	148	60
rect	147	60	148	61
rect	147	62	148	63
rect	147	63	148	64
rect	147	65	148	66
rect	147	66	148	67
rect	147	68	148	69
rect	147	69	148	70
rect	147	71	148	72
rect	147	72	148	73
rect	147	74	148	75
rect	147	75	148	76
rect	147	77	148	78
rect	147	78	148	79
rect	147	80	148	81
rect	147	81	148	82
rect	147	83	148	84
rect	147	84	148	85
rect	147	86	148	87
rect	147	87	148	88
rect	147	89	148	90
rect	147	90	148	91
rect	147	92	148	93
rect	147	93	148	94
rect	147	95	148	96
rect	147	96	148	97
rect	147	98	148	99
rect	147	99	148	100
rect	147	101	148	102
rect	147	102	148	103
rect	147	104	148	105
rect	147	105	148	106
rect	147	107	148	108
rect	147	108	148	109
rect	147	110	148	111
rect	147	111	148	112
rect	147	113	148	114
rect	147	114	148	115
rect	147	116	148	117
rect	147	117	148	118
rect	147	119	148	120
rect	147	120	148	121
rect	147	122	148	123
rect	147	123	148	124
rect	147	125	148	126
rect	147	126	148	127
rect	147	128	148	129
rect	147	129	148	130
rect	147	131	148	132
rect	147	132	148	133
rect	147	134	148	135
rect	147	135	148	136
rect	147	137	148	138
rect	147	138	148	139
rect	147	140	148	141
rect	147	141	148	142
rect	147	143	148	144
rect	147	144	148	145
rect	147	146	148	147
rect	147	147	148	148
rect	147	149	148	150
rect	147	150	148	151
rect	147	152	148	153
rect	147	153	148	154
rect	147	155	148	156
rect	147	156	148	157
rect	147	158	148	159
rect	147	159	148	160
rect	147	161	148	162
rect	147	162	148	163
rect	147	164	148	165
rect	147	165	148	166
rect	147	167	148	168
rect	147	168	148	169
rect	147	170	148	171
rect	147	171	148	172
rect	147	173	148	174
rect	147	174	148	175
rect	147	176	148	177
rect	147	177	148	178
rect	147	179	148	180
rect	147	180	148	181
rect	147	182	148	183
rect	147	183	148	184
rect	147	185	148	186
rect	147	186	148	187
rect	147	188	148	189
rect	147	189	148	190
rect	147	191	148	192
rect	147	192	148	193
rect	147	194	148	195
rect	147	195	148	196
rect	147	197	148	198
rect	147	198	148	199
rect	147	200	148	201
rect	147	201	148	202
rect	147	203	148	204
rect	147	204	148	205
rect	147	206	148	207
rect	147	207	148	208
rect	147	209	148	210
rect	147	210	148	211
rect	147	212	148	213
rect	147	213	148	214
rect	147	215	148	216
rect	147	216	148	217
rect	147	218	148	219
rect	147	219	148	220
rect	147	221	148	222
rect	147	222	148	223
rect	147	224	148	225
rect	147	225	148	226
rect	147	227	148	228
rect	147	228	148	229
rect	147	230	148	231
rect	147	231	148	232
rect	147	233	148	234
rect	147	234	148	235
rect	147	236	148	237
rect	147	237	148	238
rect	147	239	148	240
rect	147	240	148	241
rect	147	242	148	243
rect	147	243	148	244
rect	147	245	148	246
rect	147	246	148	247
rect	147	248	148	249
rect	147	249	148	250
rect	147	251	148	252
rect	147	252	148	253
rect	147	254	148	255
rect	147	255	148	256
rect	147	257	148	258
rect	147	258	148	259
rect	147	260	148	261
rect	147	261	148	262
rect	147	263	148	264
rect	147	264	148	265
rect	147	266	148	267
rect	147	267	148	268
rect	147	269	148	270
rect	147	270	148	271
rect	147	272	148	273
rect	147	273	148	274
rect	147	275	148	276
rect	147	276	148	277
rect	147	278	148	279
rect	147	279	148	280
rect	147	281	148	282
rect	147	282	148	283
rect	147	284	148	285
rect	147	285	148	286
rect	147	287	148	288
rect	147	288	148	289
rect	147	290	148	291
rect	147	291	148	292
rect	147	293	148	294
rect	147	294	148	295
rect	147	296	148	297
rect	147	297	148	298
rect	147	299	148	300
rect	147	300	148	301
rect	147	302	148	303
rect	147	303	148	304
rect	147	304	148	305
rect	147	305	148	306
rect	147	306	148	307
rect	147	308	148	309
rect	147	309	148	310
rect	147	311	148	312
rect	147	312	148	313
rect	147	314	148	315
rect	147	315	148	316
rect	147	317	148	318
rect	147	318	148	319
rect	147	320	148	321
rect	147	321	148	322
rect	147	323	148	324
rect	147	324	148	325
rect	147	326	148	327
rect	147	327	148	328
rect	147	329	148	330
rect	147	330	148	331
rect	147	332	148	333
rect	147	333	148	334
rect	147	335	148	336
rect	147	336	148	337
rect	147	337	148	338
rect	147	338	148	339
rect	147	339	148	340
rect	147	341	148	342
rect	147	342	148	343
rect	147	344	148	345
rect	147	345	148	346
rect	147	347	148	348
rect	147	348	148	349
rect	147	350	148	351
rect	147	351	148	352
rect	147	353	148	354
rect	147	354	148	355
rect	147	356	148	357
rect	147	357	148	358
rect	147	359	148	360
rect	147	360	148	361
rect	147	362	148	363
rect	147	363	148	364
rect	147	365	148	366
rect	147	366	148	367
rect	147	368	148	369
rect	147	369	148	370
rect	147	370	148	371
rect	147	371	148	372
rect	147	372	148	373
rect	147	374	148	375
rect	147	375	148	376
rect	147	377	148	378
rect	147	378	148	379
rect	147	380	148	381
rect	147	381	148	382
rect	147	382	148	383
rect	147	383	148	384
rect	147	384	148	385
rect	147	386	148	387
rect	148	0	149	1
rect	148	2	149	3
rect	148	3	149	4
rect	148	5	149	6
rect	148	6	149	7
rect	148	8	149	9
rect	148	9	149	10
rect	148	11	149	12
rect	148	12	149	13
rect	148	14	149	15
rect	148	15	149	16
rect	148	17	149	18
rect	148	18	149	19
rect	148	20	149	21
rect	148	21	149	22
rect	148	23	149	24
rect	148	24	149	25
rect	148	26	149	27
rect	148	27	149	28
rect	148	29	149	30
rect	148	30	149	31
rect	148	32	149	33
rect	148	33	149	34
rect	148	35	149	36
rect	148	36	149	37
rect	148	38	149	39
rect	148	39	149	40
rect	148	41	149	42
rect	148	42	149	43
rect	148	44	149	45
rect	148	45	149	46
rect	148	47	149	48
rect	148	48	149	49
rect	148	50	149	51
rect	148	51	149	52
rect	148	53	149	54
rect	148	54	149	55
rect	148	56	149	57
rect	148	57	149	58
rect	148	59	149	60
rect	148	60	149	61
rect	148	62	149	63
rect	148	63	149	64
rect	148	65	149	66
rect	148	66	149	67
rect	148	68	149	69
rect	148	69	149	70
rect	148	71	149	72
rect	148	72	149	73
rect	148	74	149	75
rect	148	75	149	76
rect	148	77	149	78
rect	148	78	149	79
rect	148	80	149	81
rect	148	81	149	82
rect	148	83	149	84
rect	148	84	149	85
rect	148	86	149	87
rect	148	87	149	88
rect	148	89	149	90
rect	148	90	149	91
rect	148	92	149	93
rect	148	93	149	94
rect	148	95	149	96
rect	148	96	149	97
rect	148	98	149	99
rect	148	99	149	100
rect	148	101	149	102
rect	148	102	149	103
rect	148	104	149	105
rect	148	105	149	106
rect	148	107	149	108
rect	148	108	149	109
rect	148	110	149	111
rect	148	111	149	112
rect	148	113	149	114
rect	148	114	149	115
rect	148	116	149	117
rect	148	117	149	118
rect	148	119	149	120
rect	148	120	149	121
rect	148	122	149	123
rect	148	123	149	124
rect	148	125	149	126
rect	148	126	149	127
rect	148	128	149	129
rect	148	129	149	130
rect	148	131	149	132
rect	148	132	149	133
rect	148	134	149	135
rect	148	135	149	136
rect	148	137	149	138
rect	148	138	149	139
rect	148	140	149	141
rect	148	141	149	142
rect	148	143	149	144
rect	148	144	149	145
rect	148	146	149	147
rect	148	147	149	148
rect	148	149	149	150
rect	148	150	149	151
rect	148	152	149	153
rect	148	153	149	154
rect	148	155	149	156
rect	148	156	149	157
rect	148	158	149	159
rect	148	159	149	160
rect	148	161	149	162
rect	148	162	149	163
rect	148	164	149	165
rect	148	165	149	166
rect	148	167	149	168
rect	148	168	149	169
rect	148	170	149	171
rect	148	171	149	172
rect	148	173	149	174
rect	148	174	149	175
rect	148	176	149	177
rect	148	177	149	178
rect	148	179	149	180
rect	148	180	149	181
rect	148	182	149	183
rect	148	183	149	184
rect	148	185	149	186
rect	148	186	149	187
rect	148	188	149	189
rect	148	189	149	190
rect	148	191	149	192
rect	148	192	149	193
rect	148	194	149	195
rect	148	195	149	196
rect	148	197	149	198
rect	148	198	149	199
rect	148	200	149	201
rect	148	201	149	202
rect	148	203	149	204
rect	148	204	149	205
rect	148	206	149	207
rect	148	207	149	208
rect	148	209	149	210
rect	148	210	149	211
rect	148	212	149	213
rect	148	213	149	214
rect	148	215	149	216
rect	148	216	149	217
rect	148	218	149	219
rect	148	219	149	220
rect	148	221	149	222
rect	148	222	149	223
rect	148	224	149	225
rect	148	225	149	226
rect	148	227	149	228
rect	148	228	149	229
rect	148	230	149	231
rect	148	231	149	232
rect	148	233	149	234
rect	148	234	149	235
rect	148	236	149	237
rect	148	237	149	238
rect	148	239	149	240
rect	148	240	149	241
rect	148	242	149	243
rect	148	243	149	244
rect	148	245	149	246
rect	148	246	149	247
rect	148	248	149	249
rect	148	249	149	250
rect	148	251	149	252
rect	148	252	149	253
rect	148	254	149	255
rect	148	255	149	256
rect	148	257	149	258
rect	148	258	149	259
rect	148	260	149	261
rect	148	261	149	262
rect	148	263	149	264
rect	148	264	149	265
rect	148	266	149	267
rect	148	267	149	268
rect	148	269	149	270
rect	148	270	149	271
rect	148	272	149	273
rect	148	273	149	274
rect	148	275	149	276
rect	148	276	149	277
rect	148	278	149	279
rect	148	279	149	280
rect	148	281	149	282
rect	148	282	149	283
rect	148	284	149	285
rect	148	285	149	286
rect	148	287	149	288
rect	148	288	149	289
rect	148	290	149	291
rect	148	291	149	292
rect	148	293	149	294
rect	148	294	149	295
rect	148	296	149	297
rect	148	297	149	298
rect	148	299	149	300
rect	148	300	149	301
rect	148	302	149	303
rect	148	303	149	304
rect	148	304	149	305
rect	148	305	149	306
rect	148	306	149	307
rect	148	308	149	309
rect	148	309	149	310
rect	148	311	149	312
rect	148	312	149	313
rect	148	314	149	315
rect	148	315	149	316
rect	148	317	149	318
rect	148	318	149	319
rect	148	320	149	321
rect	148	321	149	322
rect	148	323	149	324
rect	148	324	149	325
rect	148	326	149	327
rect	148	327	149	328
rect	148	329	149	330
rect	148	330	149	331
rect	148	332	149	333
rect	148	333	149	334
rect	148	335	149	336
rect	148	336	149	337
rect	148	337	149	338
rect	148	338	149	339
rect	148	339	149	340
rect	148	341	149	342
rect	148	342	149	343
rect	148	344	149	345
rect	148	345	149	346
rect	148	347	149	348
rect	148	348	149	349
rect	148	350	149	351
rect	148	351	149	352
rect	148	353	149	354
rect	148	354	149	355
rect	148	356	149	357
rect	148	357	149	358
rect	148	359	149	360
rect	148	360	149	361
rect	148	362	149	363
rect	148	363	149	364
rect	148	365	149	366
rect	148	366	149	367
rect	148	368	149	369
rect	148	369	149	370
rect	148	370	149	371
rect	148	371	149	372
rect	148	372	149	373
rect	148	374	149	375
rect	148	375	149	376
rect	148	377	149	378
rect	148	378	149	379
rect	148	380	149	381
rect	148	381	149	382
rect	148	382	149	383
rect	148	383	149	384
rect	148	384	149	385
rect	148	386	149	387
rect	149	0	150	1
rect	149	2	150	3
rect	149	3	150	4
rect	149	5	150	6
rect	149	6	150	7
rect	149	8	150	9
rect	149	9	150	10
rect	149	11	150	12
rect	149	12	150	13
rect	149	14	150	15
rect	149	15	150	16
rect	149	17	150	18
rect	149	18	150	19
rect	149	20	150	21
rect	149	21	150	22
rect	149	23	150	24
rect	149	24	150	25
rect	149	26	150	27
rect	149	27	150	28
rect	149	29	150	30
rect	149	30	150	31
rect	149	32	150	33
rect	149	33	150	34
rect	149	35	150	36
rect	149	36	150	37
rect	149	38	150	39
rect	149	39	150	40
rect	149	41	150	42
rect	149	42	150	43
rect	149	44	150	45
rect	149	45	150	46
rect	149	47	150	48
rect	149	48	150	49
rect	149	50	150	51
rect	149	51	150	52
rect	149	53	150	54
rect	149	54	150	55
rect	149	56	150	57
rect	149	57	150	58
rect	149	59	150	60
rect	149	60	150	61
rect	149	62	150	63
rect	149	63	150	64
rect	149	65	150	66
rect	149	66	150	67
rect	149	68	150	69
rect	149	69	150	70
rect	149	71	150	72
rect	149	72	150	73
rect	149	74	150	75
rect	149	75	150	76
rect	149	77	150	78
rect	149	78	150	79
rect	149	80	150	81
rect	149	81	150	82
rect	149	83	150	84
rect	149	84	150	85
rect	149	86	150	87
rect	149	87	150	88
rect	149	89	150	90
rect	149	90	150	91
rect	149	92	150	93
rect	149	93	150	94
rect	149	95	150	96
rect	149	96	150	97
rect	149	98	150	99
rect	149	99	150	100
rect	149	101	150	102
rect	149	102	150	103
rect	149	104	150	105
rect	149	105	150	106
rect	149	107	150	108
rect	149	108	150	109
rect	149	110	150	111
rect	149	111	150	112
rect	149	113	150	114
rect	149	114	150	115
rect	149	116	150	117
rect	149	117	150	118
rect	149	119	150	120
rect	149	120	150	121
rect	149	122	150	123
rect	149	123	150	124
rect	149	125	150	126
rect	149	126	150	127
rect	149	128	150	129
rect	149	129	150	130
rect	149	131	150	132
rect	149	132	150	133
rect	149	134	150	135
rect	149	135	150	136
rect	149	137	150	138
rect	149	138	150	139
rect	149	140	150	141
rect	149	141	150	142
rect	149	143	150	144
rect	149	144	150	145
rect	149	146	150	147
rect	149	147	150	148
rect	149	149	150	150
rect	149	150	150	151
rect	149	152	150	153
rect	149	153	150	154
rect	149	155	150	156
rect	149	156	150	157
rect	149	158	150	159
rect	149	159	150	160
rect	149	161	150	162
rect	149	162	150	163
rect	149	164	150	165
rect	149	165	150	166
rect	149	167	150	168
rect	149	168	150	169
rect	149	170	150	171
rect	149	171	150	172
rect	149	173	150	174
rect	149	174	150	175
rect	149	176	150	177
rect	149	177	150	178
rect	149	179	150	180
rect	149	180	150	181
rect	149	182	150	183
rect	149	183	150	184
rect	149	185	150	186
rect	149	186	150	187
rect	149	188	150	189
rect	149	189	150	190
rect	149	191	150	192
rect	149	192	150	193
rect	149	194	150	195
rect	149	195	150	196
rect	149	197	150	198
rect	149	198	150	199
rect	149	200	150	201
rect	149	201	150	202
rect	149	203	150	204
rect	149	204	150	205
rect	149	206	150	207
rect	149	207	150	208
rect	149	209	150	210
rect	149	210	150	211
rect	149	212	150	213
rect	149	213	150	214
rect	149	215	150	216
rect	149	216	150	217
rect	149	218	150	219
rect	149	219	150	220
rect	149	221	150	222
rect	149	222	150	223
rect	149	224	150	225
rect	149	225	150	226
rect	149	227	150	228
rect	149	228	150	229
rect	149	230	150	231
rect	149	231	150	232
rect	149	233	150	234
rect	149	234	150	235
rect	149	236	150	237
rect	149	237	150	238
rect	149	239	150	240
rect	149	240	150	241
rect	149	242	150	243
rect	149	243	150	244
rect	149	245	150	246
rect	149	246	150	247
rect	149	248	150	249
rect	149	249	150	250
rect	149	251	150	252
rect	149	252	150	253
rect	149	254	150	255
rect	149	255	150	256
rect	149	257	150	258
rect	149	258	150	259
rect	149	260	150	261
rect	149	261	150	262
rect	149	263	150	264
rect	149	264	150	265
rect	149	266	150	267
rect	149	267	150	268
rect	149	269	150	270
rect	149	270	150	271
rect	149	272	150	273
rect	149	273	150	274
rect	149	275	150	276
rect	149	276	150	277
rect	149	278	150	279
rect	149	279	150	280
rect	149	281	150	282
rect	149	282	150	283
rect	149	284	150	285
rect	149	285	150	286
rect	149	287	150	288
rect	149	288	150	289
rect	149	290	150	291
rect	149	291	150	292
rect	149	293	150	294
rect	149	294	150	295
rect	149	296	150	297
rect	149	297	150	298
rect	149	299	150	300
rect	149	300	150	301
rect	149	302	150	303
rect	149	303	150	304
rect	149	304	150	305
rect	149	305	150	306
rect	149	306	150	307
rect	149	308	150	309
rect	149	309	150	310
rect	149	311	150	312
rect	149	312	150	313
rect	149	314	150	315
rect	149	315	150	316
rect	149	317	150	318
rect	149	318	150	319
rect	149	320	150	321
rect	149	321	150	322
rect	149	323	150	324
rect	149	324	150	325
rect	149	326	150	327
rect	149	327	150	328
rect	149	329	150	330
rect	149	330	150	331
rect	149	332	150	333
rect	149	333	150	334
rect	149	335	150	336
rect	149	336	150	337
rect	149	337	150	338
rect	149	338	150	339
rect	149	339	150	340
rect	149	341	150	342
rect	149	342	150	343
rect	149	344	150	345
rect	149	345	150	346
rect	149	347	150	348
rect	149	348	150	349
rect	149	350	150	351
rect	149	351	150	352
rect	149	353	150	354
rect	149	354	150	355
rect	149	356	150	357
rect	149	357	150	358
rect	149	359	150	360
rect	149	360	150	361
rect	149	362	150	363
rect	149	363	150	364
rect	149	365	150	366
rect	149	366	150	367
rect	149	368	150	369
rect	149	369	150	370
rect	149	370	150	371
rect	149	371	150	372
rect	149	372	150	373
rect	149	374	150	375
rect	149	375	150	376
rect	149	377	150	378
rect	149	378	150	379
rect	149	380	150	381
rect	149	381	150	382
rect	149	382	150	383
rect	149	383	150	384
rect	149	384	150	385
rect	149	386	150	387
rect	160	0	161	1
rect	160	2	161	3
rect	160	3	161	4
rect	160	5	161	6
rect	160	6	161	7
rect	160	8	161	9
rect	160	9	161	10
rect	160	11	161	12
rect	160	12	161	13
rect	160	14	161	15
rect	160	15	161	16
rect	160	17	161	18
rect	160	18	161	19
rect	160	20	161	21
rect	160	21	161	22
rect	160	23	161	24
rect	160	24	161	25
rect	160	26	161	27
rect	160	27	161	28
rect	160	29	161	30
rect	160	30	161	31
rect	160	32	161	33
rect	160	33	161	34
rect	160	35	161	36
rect	160	36	161	37
rect	160	38	161	39
rect	160	39	161	40
rect	160	41	161	42
rect	160	42	161	43
rect	160	44	161	45
rect	160	45	161	46
rect	160	47	161	48
rect	160	48	161	49
rect	160	50	161	51
rect	160	51	161	52
rect	160	53	161	54
rect	160	54	161	55
rect	160	56	161	57
rect	160	57	161	58
rect	160	59	161	60
rect	160	60	161	61
rect	160	62	161	63
rect	160	63	161	64
rect	160	65	161	66
rect	160	66	161	67
rect	160	68	161	69
rect	160	69	161	70
rect	160	71	161	72
rect	160	72	161	73
rect	160	74	161	75
rect	160	75	161	76
rect	160	77	161	78
rect	160	78	161	79
rect	160	80	161	81
rect	160	81	161	82
rect	160	83	161	84
rect	160	84	161	85
rect	160	86	161	87
rect	160	87	161	88
rect	160	89	161	90
rect	160	90	161	91
rect	160	92	161	93
rect	160	93	161	94
rect	160	95	161	96
rect	160	96	161	97
rect	160	98	161	99
rect	160	99	161	100
rect	160	101	161	102
rect	160	102	161	103
rect	160	104	161	105
rect	160	105	161	106
rect	160	107	161	108
rect	160	108	161	109
rect	160	110	161	111
rect	160	111	161	112
rect	160	113	161	114
rect	160	114	161	115
rect	160	116	161	117
rect	160	117	161	118
rect	160	119	161	120
rect	160	120	161	121
rect	160	122	161	123
rect	160	123	161	124
rect	160	125	161	126
rect	160	126	161	127
rect	160	128	161	129
rect	160	129	161	130
rect	160	131	161	132
rect	160	132	161	133
rect	160	134	161	135
rect	160	135	161	136
rect	160	137	161	138
rect	160	138	161	139
rect	160	140	161	141
rect	160	141	161	142
rect	160	143	161	144
rect	160	144	161	145
rect	160	146	161	147
rect	160	147	161	148
rect	160	149	161	150
rect	160	150	161	151
rect	160	152	161	153
rect	160	153	161	154
rect	160	155	161	156
rect	160	156	161	157
rect	160	158	161	159
rect	160	159	161	160
rect	160	161	161	162
rect	160	162	161	163
rect	160	164	161	165
rect	160	165	161	166
rect	160	167	161	168
rect	160	168	161	169
rect	160	170	161	171
rect	160	171	161	172
rect	160	173	161	174
rect	160	174	161	175
rect	160	176	161	177
rect	160	177	161	178
rect	160	179	161	180
rect	160	180	161	181
rect	160	182	161	183
rect	160	183	161	184
rect	160	185	161	186
rect	160	186	161	187
rect	160	188	161	189
rect	160	189	161	190
rect	160	191	161	192
rect	160	192	161	193
rect	160	194	161	195
rect	160	195	161	196
rect	160	197	161	198
rect	160	198	161	199
rect	160	200	161	201
rect	160	201	161	202
rect	160	203	161	204
rect	160	204	161	205
rect	160	206	161	207
rect	160	207	161	208
rect	160	209	161	210
rect	160	210	161	211
rect	160	212	161	213
rect	160	213	161	214
rect	160	215	161	216
rect	160	216	161	217
rect	160	218	161	219
rect	160	219	161	220
rect	160	221	161	222
rect	160	222	161	223
rect	160	224	161	225
rect	160	225	161	226
rect	160	227	161	228
rect	160	228	161	229
rect	160	230	161	231
rect	160	231	161	232
rect	160	233	161	234
rect	160	234	161	235
rect	160	236	161	237
rect	160	237	161	238
rect	160	239	161	240
rect	160	240	161	241
rect	160	242	161	243
rect	160	243	161	244
rect	160	245	161	246
rect	160	246	161	247
rect	160	248	161	249
rect	160	249	161	250
rect	160	251	161	252
rect	160	252	161	253
rect	160	254	161	255
rect	160	255	161	256
rect	160	257	161	258
rect	160	258	161	259
rect	160	260	161	261
rect	160	261	161	262
rect	160	263	161	264
rect	160	264	161	265
rect	160	266	161	267
rect	160	267	161	268
rect	160	269	161	270
rect	160	270	161	271
rect	160	272	161	273
rect	160	273	161	274
rect	160	275	161	276
rect	160	276	161	277
rect	160	278	161	279
rect	160	279	161	280
rect	160	281	161	282
rect	160	282	161	283
rect	160	284	161	285
rect	160	285	161	286
rect	160	287	161	288
rect	160	288	161	289
rect	160	290	161	291
rect	160	291	161	292
rect	160	293	161	294
rect	160	294	161	295
rect	160	296	161	297
rect	160	297	161	298
rect	160	299	161	300
rect	160	300	161	301
rect	160	302	161	303
rect	160	303	161	304
rect	160	304	161	305
rect	160	305	161	306
rect	160	306	161	307
rect	160	308	161	309
rect	160	309	161	310
rect	160	311	161	312
rect	160	312	161	313
rect	160	314	161	315
rect	160	315	161	316
rect	160	317	161	318
rect	160	318	161	319
rect	160	320	161	321
rect	160	321	161	322
rect	160	323	161	324
rect	160	324	161	325
rect	160	326	161	327
rect	160	327	161	328
rect	160	328	161	329
rect	160	329	161	330
rect	160	330	161	331
rect	160	332	161	333
rect	160	333	161	334
rect	160	335	161	336
rect	160	336	161	337
rect	160	337	161	338
rect	160	338	161	339
rect	160	339	161	340
rect	160	340	161	341
rect	160	341	161	342
rect	160	342	161	343
rect	160	343	161	344
rect	160	344	161	345
rect	160	345	161	346
rect	160	347	161	348
rect	160	348	161	349
rect	160	350	161	351
rect	160	351	161	352
rect	160	353	161	354
rect	160	354	161	355
rect	160	356	161	357
rect	160	357	161	358
rect	160	359	161	360
rect	160	360	161	361
rect	160	362	161	363
rect	160	363	161	364
rect	160	365	161	366
rect	160	366	161	367
rect	160	368	161	369
rect	160	369	161	370
rect	160	370	161	371
rect	160	371	161	372
rect	160	372	161	373
rect	160	373	161	374
rect	160	374	161	375
rect	160	375	161	376
rect	160	376	161	377
rect	160	377	161	378
rect	160	378	161	379
rect	160	379	161	380
rect	160	380	161	381
rect	160	381	161	382
rect	160	382	161	383
rect	160	383	161	384
rect	160	384	161	385
rect	160	385	161	386
rect	160	386	161	387
rect	162	0	163	1
rect	162	2	163	3
rect	162	3	163	4
rect	162	5	163	6
rect	162	6	163	7
rect	162	8	163	9
rect	162	9	163	10
rect	162	11	163	12
rect	162	12	163	13
rect	162	14	163	15
rect	162	15	163	16
rect	162	17	163	18
rect	162	18	163	19
rect	162	20	163	21
rect	162	21	163	22
rect	162	23	163	24
rect	162	24	163	25
rect	162	26	163	27
rect	162	27	163	28
rect	162	29	163	30
rect	162	30	163	31
rect	162	32	163	33
rect	162	33	163	34
rect	162	35	163	36
rect	162	36	163	37
rect	162	38	163	39
rect	162	39	163	40
rect	162	41	163	42
rect	162	42	163	43
rect	162	44	163	45
rect	162	45	163	46
rect	162	47	163	48
rect	162	48	163	49
rect	162	50	163	51
rect	162	51	163	52
rect	162	53	163	54
rect	162	54	163	55
rect	162	56	163	57
rect	162	57	163	58
rect	162	59	163	60
rect	162	60	163	61
rect	162	62	163	63
rect	162	63	163	64
rect	162	65	163	66
rect	162	66	163	67
rect	162	68	163	69
rect	162	69	163	70
rect	162	71	163	72
rect	162	72	163	73
rect	162	74	163	75
rect	162	75	163	76
rect	162	77	163	78
rect	162	78	163	79
rect	162	80	163	81
rect	162	81	163	82
rect	162	83	163	84
rect	162	84	163	85
rect	162	86	163	87
rect	162	87	163	88
rect	162	89	163	90
rect	162	90	163	91
rect	162	92	163	93
rect	162	93	163	94
rect	162	95	163	96
rect	162	96	163	97
rect	162	98	163	99
rect	162	99	163	100
rect	162	101	163	102
rect	162	102	163	103
rect	162	104	163	105
rect	162	105	163	106
rect	162	107	163	108
rect	162	108	163	109
rect	162	110	163	111
rect	162	111	163	112
rect	162	113	163	114
rect	162	114	163	115
rect	162	116	163	117
rect	162	117	163	118
rect	162	119	163	120
rect	162	120	163	121
rect	162	122	163	123
rect	162	123	163	124
rect	162	125	163	126
rect	162	126	163	127
rect	162	128	163	129
rect	162	129	163	130
rect	162	131	163	132
rect	162	132	163	133
rect	162	134	163	135
rect	162	135	163	136
rect	162	137	163	138
rect	162	138	163	139
rect	162	140	163	141
rect	162	141	163	142
rect	162	143	163	144
rect	162	144	163	145
rect	162	146	163	147
rect	162	147	163	148
rect	162	149	163	150
rect	162	150	163	151
rect	162	152	163	153
rect	162	153	163	154
rect	162	155	163	156
rect	162	156	163	157
rect	162	158	163	159
rect	162	159	163	160
rect	162	161	163	162
rect	162	162	163	163
rect	162	164	163	165
rect	162	165	163	166
rect	162	167	163	168
rect	162	168	163	169
rect	162	170	163	171
rect	162	171	163	172
rect	162	173	163	174
rect	162	174	163	175
rect	162	176	163	177
rect	162	177	163	178
rect	162	179	163	180
rect	162	180	163	181
rect	162	182	163	183
rect	162	183	163	184
rect	162	185	163	186
rect	162	186	163	187
rect	162	188	163	189
rect	162	189	163	190
rect	162	191	163	192
rect	162	192	163	193
rect	162	194	163	195
rect	162	195	163	196
rect	162	197	163	198
rect	162	198	163	199
rect	162	200	163	201
rect	162	201	163	202
rect	162	203	163	204
rect	162	204	163	205
rect	162	206	163	207
rect	162	207	163	208
rect	162	209	163	210
rect	162	210	163	211
rect	162	212	163	213
rect	162	213	163	214
rect	162	215	163	216
rect	162	216	163	217
rect	162	218	163	219
rect	162	219	163	220
rect	162	221	163	222
rect	162	222	163	223
rect	162	224	163	225
rect	162	225	163	226
rect	162	227	163	228
rect	162	228	163	229
rect	162	230	163	231
rect	162	231	163	232
rect	162	233	163	234
rect	162	234	163	235
rect	162	236	163	237
rect	162	237	163	238
rect	162	239	163	240
rect	162	240	163	241
rect	162	242	163	243
rect	162	243	163	244
rect	162	245	163	246
rect	162	246	163	247
rect	162	248	163	249
rect	162	249	163	250
rect	162	251	163	252
rect	162	252	163	253
rect	162	254	163	255
rect	162	255	163	256
rect	162	257	163	258
rect	162	258	163	259
rect	162	260	163	261
rect	162	261	163	262
rect	162	263	163	264
rect	162	264	163	265
rect	162	266	163	267
rect	162	267	163	268
rect	162	269	163	270
rect	162	270	163	271
rect	162	272	163	273
rect	162	273	163	274
rect	162	275	163	276
rect	162	276	163	277
rect	162	278	163	279
rect	162	279	163	280
rect	162	281	163	282
rect	162	282	163	283
rect	162	284	163	285
rect	162	285	163	286
rect	162	287	163	288
rect	162	288	163	289
rect	162	290	163	291
rect	162	291	163	292
rect	162	293	163	294
rect	162	294	163	295
rect	162	296	163	297
rect	162	297	163	298
rect	162	299	163	300
rect	162	300	163	301
rect	162	302	163	303
rect	162	303	163	304
rect	162	304	163	305
rect	162	305	163	306
rect	162	306	163	307
rect	162	308	163	309
rect	162	309	163	310
rect	162	311	163	312
rect	162	312	163	313
rect	162	314	163	315
rect	162	315	163	316
rect	162	317	163	318
rect	162	318	163	319
rect	162	320	163	321
rect	162	321	163	322
rect	162	323	163	324
rect	162	324	163	325
rect	162	326	163	327
rect	162	327	163	328
rect	162	328	163	329
rect	162	329	163	330
rect	162	330	163	331
rect	162	332	163	333
rect	162	333	163	334
rect	162	335	163	336
rect	162	336	163	337
rect	162	337	163	338
rect	162	338	163	339
rect	162	339	163	340
rect	162	340	163	341
rect	162	341	163	342
rect	162	342	163	343
rect	162	343	163	344
rect	162	344	163	345
rect	162	345	163	346
rect	162	347	163	348
rect	162	348	163	349
rect	162	350	163	351
rect	162	351	163	352
rect	162	353	163	354
rect	162	354	163	355
rect	162	356	163	357
rect	162	357	163	358
rect	162	359	163	360
rect	162	360	163	361
rect	162	362	163	363
rect	162	363	163	364
rect	162	365	163	366
rect	162	366	163	367
rect	162	368	163	369
rect	163	0	164	1
rect	163	2	164	3
rect	163	3	164	4
rect	163	5	164	6
rect	163	6	164	7
rect	163	8	164	9
rect	163	9	164	10
rect	163	11	164	12
rect	163	12	164	13
rect	163	14	164	15
rect	163	15	164	16
rect	163	17	164	18
rect	163	18	164	19
rect	163	20	164	21
rect	163	21	164	22
rect	163	23	164	24
rect	163	24	164	25
rect	163	26	164	27
rect	163	27	164	28
rect	163	29	164	30
rect	163	30	164	31
rect	163	32	164	33
rect	163	33	164	34
rect	163	35	164	36
rect	163	36	164	37
rect	163	38	164	39
rect	163	39	164	40
rect	163	41	164	42
rect	163	42	164	43
rect	163	44	164	45
rect	163	45	164	46
rect	163	47	164	48
rect	163	48	164	49
rect	163	50	164	51
rect	163	51	164	52
rect	163	53	164	54
rect	163	54	164	55
rect	163	56	164	57
rect	163	57	164	58
rect	163	59	164	60
rect	163	60	164	61
rect	163	62	164	63
rect	163	63	164	64
rect	163	65	164	66
rect	163	66	164	67
rect	163	68	164	69
rect	163	69	164	70
rect	163	71	164	72
rect	163	72	164	73
rect	163	74	164	75
rect	163	75	164	76
rect	163	77	164	78
rect	163	78	164	79
rect	163	80	164	81
rect	163	81	164	82
rect	163	83	164	84
rect	163	84	164	85
rect	163	86	164	87
rect	163	87	164	88
rect	163	89	164	90
rect	163	90	164	91
rect	163	92	164	93
rect	163	93	164	94
rect	163	95	164	96
rect	163	96	164	97
rect	163	98	164	99
rect	163	99	164	100
rect	163	101	164	102
rect	163	102	164	103
rect	163	104	164	105
rect	163	105	164	106
rect	163	107	164	108
rect	163	108	164	109
rect	163	110	164	111
rect	163	111	164	112
rect	163	113	164	114
rect	163	114	164	115
rect	163	116	164	117
rect	163	117	164	118
rect	163	119	164	120
rect	163	120	164	121
rect	163	122	164	123
rect	163	123	164	124
rect	163	125	164	126
rect	163	126	164	127
rect	163	128	164	129
rect	163	129	164	130
rect	163	131	164	132
rect	163	132	164	133
rect	163	134	164	135
rect	163	135	164	136
rect	163	137	164	138
rect	163	138	164	139
rect	163	140	164	141
rect	163	141	164	142
rect	163	143	164	144
rect	163	144	164	145
rect	163	146	164	147
rect	163	147	164	148
rect	163	149	164	150
rect	163	150	164	151
rect	163	152	164	153
rect	163	153	164	154
rect	163	155	164	156
rect	163	156	164	157
rect	163	158	164	159
rect	163	159	164	160
rect	163	161	164	162
rect	163	162	164	163
rect	163	164	164	165
rect	163	165	164	166
rect	163	167	164	168
rect	163	168	164	169
rect	163	170	164	171
rect	163	171	164	172
rect	163	173	164	174
rect	163	174	164	175
rect	163	176	164	177
rect	163	177	164	178
rect	163	179	164	180
rect	163	180	164	181
rect	163	182	164	183
rect	163	183	164	184
rect	163	185	164	186
rect	163	186	164	187
rect	163	188	164	189
rect	163	189	164	190
rect	163	191	164	192
rect	163	192	164	193
rect	163	194	164	195
rect	163	195	164	196
rect	163	197	164	198
rect	163	198	164	199
rect	163	200	164	201
rect	163	201	164	202
rect	163	203	164	204
rect	163	204	164	205
rect	163	206	164	207
rect	163	207	164	208
rect	163	209	164	210
rect	163	210	164	211
rect	163	212	164	213
rect	163	213	164	214
rect	163	215	164	216
rect	163	216	164	217
rect	163	218	164	219
rect	163	219	164	220
rect	163	221	164	222
rect	163	222	164	223
rect	163	224	164	225
rect	163	225	164	226
rect	163	227	164	228
rect	163	228	164	229
rect	163	230	164	231
rect	163	231	164	232
rect	163	233	164	234
rect	163	234	164	235
rect	163	236	164	237
rect	163	237	164	238
rect	163	239	164	240
rect	163	240	164	241
rect	163	242	164	243
rect	163	243	164	244
rect	163	245	164	246
rect	163	246	164	247
rect	163	248	164	249
rect	163	249	164	250
rect	163	251	164	252
rect	163	252	164	253
rect	163	254	164	255
rect	163	255	164	256
rect	163	257	164	258
rect	163	258	164	259
rect	163	260	164	261
rect	163	261	164	262
rect	163	263	164	264
rect	163	264	164	265
rect	163	266	164	267
rect	163	267	164	268
rect	163	269	164	270
rect	163	270	164	271
rect	163	272	164	273
rect	163	273	164	274
rect	163	275	164	276
rect	163	276	164	277
rect	163	278	164	279
rect	163	279	164	280
rect	163	281	164	282
rect	163	282	164	283
rect	163	284	164	285
rect	163	285	164	286
rect	163	287	164	288
rect	163	288	164	289
rect	163	290	164	291
rect	163	291	164	292
rect	163	293	164	294
rect	163	294	164	295
rect	163	296	164	297
rect	163	297	164	298
rect	163	299	164	300
rect	163	300	164	301
rect	163	302	164	303
rect	163	303	164	304
rect	163	304	164	305
rect	163	305	164	306
rect	163	306	164	307
rect	163	308	164	309
rect	163	309	164	310
rect	163	311	164	312
rect	163	312	164	313
rect	163	314	164	315
rect	163	315	164	316
rect	163	317	164	318
rect	163	318	164	319
rect	163	320	164	321
rect	163	321	164	322
rect	163	323	164	324
rect	163	324	164	325
rect	163	326	164	327
rect	163	327	164	328
rect	163	328	164	329
rect	163	329	164	330
rect	163	330	164	331
rect	163	332	164	333
rect	163	333	164	334
rect	163	335	164	336
rect	163	336	164	337
rect	163	337	164	338
rect	163	338	164	339
rect	163	339	164	340
rect	163	340	164	341
rect	163	341	164	342
rect	163	342	164	343
rect	163	343	164	344
rect	163	344	164	345
rect	163	345	164	346
rect	163	347	164	348
rect	163	348	164	349
rect	163	350	164	351
rect	163	351	164	352
rect	163	353	164	354
rect	163	354	164	355
rect	163	356	164	357
rect	163	357	164	358
rect	163	359	164	360
rect	163	360	164	361
rect	163	362	164	363
rect	163	363	164	364
rect	163	365	164	366
rect	163	366	164	367
rect	163	368	164	369
rect	164	0	165	1
rect	164	2	165	3
rect	164	3	165	4
rect	164	5	165	6
rect	164	6	165	7
rect	164	8	165	9
rect	164	9	165	10
rect	164	11	165	12
rect	164	12	165	13
rect	164	14	165	15
rect	164	15	165	16
rect	164	17	165	18
rect	164	18	165	19
rect	164	20	165	21
rect	164	21	165	22
rect	164	23	165	24
rect	164	24	165	25
rect	164	26	165	27
rect	164	27	165	28
rect	164	29	165	30
rect	164	30	165	31
rect	164	32	165	33
rect	164	33	165	34
rect	164	35	165	36
rect	164	36	165	37
rect	164	38	165	39
rect	164	39	165	40
rect	164	41	165	42
rect	164	42	165	43
rect	164	44	165	45
rect	164	45	165	46
rect	164	47	165	48
rect	164	48	165	49
rect	164	50	165	51
rect	164	51	165	52
rect	164	53	165	54
rect	164	54	165	55
rect	164	56	165	57
rect	164	57	165	58
rect	164	59	165	60
rect	164	60	165	61
rect	164	62	165	63
rect	164	63	165	64
rect	164	65	165	66
rect	164	66	165	67
rect	164	68	165	69
rect	164	69	165	70
rect	164	71	165	72
rect	164	72	165	73
rect	164	74	165	75
rect	164	75	165	76
rect	164	77	165	78
rect	164	78	165	79
rect	164	80	165	81
rect	164	81	165	82
rect	164	83	165	84
rect	164	84	165	85
rect	164	86	165	87
rect	164	87	165	88
rect	164	89	165	90
rect	164	90	165	91
rect	164	92	165	93
rect	164	93	165	94
rect	164	95	165	96
rect	164	96	165	97
rect	164	98	165	99
rect	164	99	165	100
rect	164	101	165	102
rect	164	102	165	103
rect	164	104	165	105
rect	164	105	165	106
rect	164	107	165	108
rect	164	108	165	109
rect	164	110	165	111
rect	164	111	165	112
rect	164	113	165	114
rect	164	114	165	115
rect	164	116	165	117
rect	164	117	165	118
rect	164	119	165	120
rect	164	120	165	121
rect	164	122	165	123
rect	164	123	165	124
rect	164	125	165	126
rect	164	126	165	127
rect	164	128	165	129
rect	164	129	165	130
rect	164	131	165	132
rect	164	132	165	133
rect	164	134	165	135
rect	164	135	165	136
rect	164	137	165	138
rect	164	138	165	139
rect	164	140	165	141
rect	164	141	165	142
rect	164	143	165	144
rect	164	144	165	145
rect	164	146	165	147
rect	164	147	165	148
rect	164	149	165	150
rect	164	150	165	151
rect	164	152	165	153
rect	164	153	165	154
rect	164	155	165	156
rect	164	156	165	157
rect	164	158	165	159
rect	164	159	165	160
rect	164	161	165	162
rect	164	162	165	163
rect	164	164	165	165
rect	164	165	165	166
rect	164	167	165	168
rect	164	168	165	169
rect	164	170	165	171
rect	164	171	165	172
rect	164	173	165	174
rect	164	174	165	175
rect	164	176	165	177
rect	164	177	165	178
rect	164	179	165	180
rect	164	180	165	181
rect	164	182	165	183
rect	164	183	165	184
rect	164	185	165	186
rect	164	186	165	187
rect	164	188	165	189
rect	164	189	165	190
rect	164	191	165	192
rect	164	192	165	193
rect	164	194	165	195
rect	164	195	165	196
rect	164	197	165	198
rect	164	198	165	199
rect	164	200	165	201
rect	164	201	165	202
rect	164	203	165	204
rect	164	204	165	205
rect	164	206	165	207
rect	164	207	165	208
rect	164	209	165	210
rect	164	210	165	211
rect	164	212	165	213
rect	164	213	165	214
rect	164	215	165	216
rect	164	216	165	217
rect	164	218	165	219
rect	164	219	165	220
rect	164	221	165	222
rect	164	222	165	223
rect	164	224	165	225
rect	164	225	165	226
rect	164	227	165	228
rect	164	228	165	229
rect	164	230	165	231
rect	164	231	165	232
rect	164	233	165	234
rect	164	234	165	235
rect	164	236	165	237
rect	164	237	165	238
rect	164	239	165	240
rect	164	240	165	241
rect	164	242	165	243
rect	164	243	165	244
rect	164	245	165	246
rect	164	246	165	247
rect	164	248	165	249
rect	164	249	165	250
rect	164	251	165	252
rect	164	252	165	253
rect	164	254	165	255
rect	164	255	165	256
rect	164	257	165	258
rect	164	258	165	259
rect	164	260	165	261
rect	164	261	165	262
rect	164	263	165	264
rect	164	264	165	265
rect	164	266	165	267
rect	164	267	165	268
rect	164	269	165	270
rect	164	270	165	271
rect	164	272	165	273
rect	164	273	165	274
rect	164	275	165	276
rect	164	276	165	277
rect	164	278	165	279
rect	164	279	165	280
rect	164	281	165	282
rect	164	282	165	283
rect	164	284	165	285
rect	164	285	165	286
rect	164	287	165	288
rect	164	288	165	289
rect	164	290	165	291
rect	164	291	165	292
rect	164	293	165	294
rect	164	294	165	295
rect	164	296	165	297
rect	164	297	165	298
rect	164	299	165	300
rect	164	300	165	301
rect	164	302	165	303
rect	164	303	165	304
rect	164	304	165	305
rect	164	305	165	306
rect	164	306	165	307
rect	164	308	165	309
rect	164	309	165	310
rect	164	311	165	312
rect	164	312	165	313
rect	164	314	165	315
rect	164	315	165	316
rect	164	317	165	318
rect	164	318	165	319
rect	164	320	165	321
rect	164	321	165	322
rect	164	323	165	324
rect	164	324	165	325
rect	164	326	165	327
rect	164	327	165	328
rect	164	328	165	329
rect	164	329	165	330
rect	164	330	165	331
rect	164	332	165	333
rect	164	333	165	334
rect	164	335	165	336
rect	164	336	165	337
rect	164	337	165	338
rect	164	338	165	339
rect	164	339	165	340
rect	164	340	165	341
rect	164	341	165	342
rect	164	342	165	343
rect	164	343	165	344
rect	164	344	165	345
rect	164	345	165	346
rect	164	347	165	348
rect	164	348	165	349
rect	164	350	165	351
rect	164	351	165	352
rect	164	353	165	354
rect	164	354	165	355
rect	164	356	165	357
rect	164	357	165	358
rect	164	359	165	360
rect	164	360	165	361
rect	164	362	165	363
rect	164	363	165	364
rect	164	365	165	366
rect	164	366	165	367
rect	164	368	165	369
rect	165	0	166	1
rect	165	2	166	3
rect	165	3	166	4
rect	165	5	166	6
rect	165	6	166	7
rect	165	8	166	9
rect	165	9	166	10
rect	165	11	166	12
rect	165	12	166	13
rect	165	14	166	15
rect	165	15	166	16
rect	165	17	166	18
rect	165	18	166	19
rect	165	20	166	21
rect	165	21	166	22
rect	165	23	166	24
rect	165	24	166	25
rect	165	26	166	27
rect	165	27	166	28
rect	165	29	166	30
rect	165	30	166	31
rect	165	32	166	33
rect	165	33	166	34
rect	165	35	166	36
rect	165	36	166	37
rect	165	38	166	39
rect	165	39	166	40
rect	165	41	166	42
rect	165	42	166	43
rect	165	44	166	45
rect	165	45	166	46
rect	165	47	166	48
rect	165	48	166	49
rect	165	50	166	51
rect	165	51	166	52
rect	165	53	166	54
rect	165	54	166	55
rect	165	56	166	57
rect	165	57	166	58
rect	165	59	166	60
rect	165	60	166	61
rect	165	62	166	63
rect	165	63	166	64
rect	165	65	166	66
rect	165	66	166	67
rect	165	68	166	69
rect	165	69	166	70
rect	165	71	166	72
rect	165	72	166	73
rect	165	74	166	75
rect	165	75	166	76
rect	165	77	166	78
rect	165	78	166	79
rect	165	80	166	81
rect	165	81	166	82
rect	165	83	166	84
rect	165	84	166	85
rect	165	86	166	87
rect	165	87	166	88
rect	165	89	166	90
rect	165	90	166	91
rect	165	92	166	93
rect	165	93	166	94
rect	165	95	166	96
rect	165	96	166	97
rect	165	98	166	99
rect	165	99	166	100
rect	165	101	166	102
rect	165	102	166	103
rect	165	104	166	105
rect	165	105	166	106
rect	165	107	166	108
rect	165	108	166	109
rect	165	110	166	111
rect	165	111	166	112
rect	165	113	166	114
rect	165	114	166	115
rect	165	116	166	117
rect	165	117	166	118
rect	165	119	166	120
rect	165	120	166	121
rect	165	122	166	123
rect	165	123	166	124
rect	165	125	166	126
rect	165	126	166	127
rect	165	128	166	129
rect	165	129	166	130
rect	165	131	166	132
rect	165	132	166	133
rect	165	134	166	135
rect	165	135	166	136
rect	165	137	166	138
rect	165	138	166	139
rect	165	140	166	141
rect	165	141	166	142
rect	165	143	166	144
rect	165	144	166	145
rect	165	146	166	147
rect	165	147	166	148
rect	165	149	166	150
rect	165	150	166	151
rect	165	152	166	153
rect	165	153	166	154
rect	165	155	166	156
rect	165	156	166	157
rect	165	158	166	159
rect	165	159	166	160
rect	165	161	166	162
rect	165	162	166	163
rect	165	164	166	165
rect	165	165	166	166
rect	165	167	166	168
rect	165	168	166	169
rect	165	170	166	171
rect	165	171	166	172
rect	165	173	166	174
rect	165	174	166	175
rect	165	176	166	177
rect	165	177	166	178
rect	165	179	166	180
rect	165	180	166	181
rect	165	182	166	183
rect	165	183	166	184
rect	165	185	166	186
rect	165	186	166	187
rect	165	188	166	189
rect	165	189	166	190
rect	165	191	166	192
rect	165	192	166	193
rect	165	194	166	195
rect	165	195	166	196
rect	165	197	166	198
rect	165	198	166	199
rect	165	200	166	201
rect	165	201	166	202
rect	165	203	166	204
rect	165	204	166	205
rect	165	206	166	207
rect	165	207	166	208
rect	165	209	166	210
rect	165	210	166	211
rect	165	212	166	213
rect	165	213	166	214
rect	165	215	166	216
rect	165	216	166	217
rect	165	218	166	219
rect	165	219	166	220
rect	165	221	166	222
rect	165	222	166	223
rect	165	224	166	225
rect	165	225	166	226
rect	165	227	166	228
rect	165	228	166	229
rect	165	230	166	231
rect	165	231	166	232
rect	165	233	166	234
rect	165	234	166	235
rect	165	236	166	237
rect	165	237	166	238
rect	165	239	166	240
rect	165	240	166	241
rect	165	242	166	243
rect	165	243	166	244
rect	165	245	166	246
rect	165	246	166	247
rect	165	248	166	249
rect	165	249	166	250
rect	165	251	166	252
rect	165	252	166	253
rect	165	254	166	255
rect	165	255	166	256
rect	165	257	166	258
rect	165	258	166	259
rect	165	260	166	261
rect	165	261	166	262
rect	165	263	166	264
rect	165	264	166	265
rect	165	266	166	267
rect	165	267	166	268
rect	165	269	166	270
rect	165	270	166	271
rect	165	272	166	273
rect	165	273	166	274
rect	165	275	166	276
rect	165	276	166	277
rect	165	278	166	279
rect	165	279	166	280
rect	165	281	166	282
rect	165	282	166	283
rect	165	284	166	285
rect	165	285	166	286
rect	165	287	166	288
rect	165	288	166	289
rect	165	290	166	291
rect	165	291	166	292
rect	165	293	166	294
rect	165	294	166	295
rect	165	296	166	297
rect	165	297	166	298
rect	165	299	166	300
rect	165	300	166	301
rect	165	302	166	303
rect	165	303	166	304
rect	165	304	166	305
rect	165	305	166	306
rect	165	306	166	307
rect	165	308	166	309
rect	165	309	166	310
rect	165	311	166	312
rect	165	312	166	313
rect	165	314	166	315
rect	165	315	166	316
rect	165	317	166	318
rect	165	318	166	319
rect	165	320	166	321
rect	165	321	166	322
rect	165	323	166	324
rect	165	324	166	325
rect	165	326	166	327
rect	165	327	166	328
rect	165	328	166	329
rect	165	329	166	330
rect	165	330	166	331
rect	165	332	166	333
rect	165	333	166	334
rect	165	335	166	336
rect	165	336	166	337
rect	165	337	166	338
rect	165	338	166	339
rect	165	339	166	340
rect	165	340	166	341
rect	165	341	166	342
rect	165	342	166	343
rect	165	343	166	344
rect	165	344	166	345
rect	165	345	166	346
rect	165	347	166	348
rect	165	348	166	349
rect	165	350	166	351
rect	165	351	166	352
rect	165	353	166	354
rect	165	354	166	355
rect	165	356	166	357
rect	165	357	166	358
rect	165	359	166	360
rect	165	360	166	361
rect	165	362	166	363
rect	165	363	166	364
rect	165	365	166	366
rect	165	366	166	367
rect	165	368	166	369
rect	166	0	167	1
rect	166	2	167	3
rect	166	3	167	4
rect	166	5	167	6
rect	166	6	167	7
rect	166	8	167	9
rect	166	9	167	10
rect	166	11	167	12
rect	166	12	167	13
rect	166	14	167	15
rect	166	15	167	16
rect	166	17	167	18
rect	166	18	167	19
rect	166	20	167	21
rect	166	21	167	22
rect	166	23	167	24
rect	166	24	167	25
rect	166	26	167	27
rect	166	27	167	28
rect	166	29	167	30
rect	166	30	167	31
rect	166	32	167	33
rect	166	33	167	34
rect	166	35	167	36
rect	166	36	167	37
rect	166	38	167	39
rect	166	39	167	40
rect	166	41	167	42
rect	166	42	167	43
rect	166	44	167	45
rect	166	45	167	46
rect	166	47	167	48
rect	166	48	167	49
rect	166	50	167	51
rect	166	51	167	52
rect	166	53	167	54
rect	166	54	167	55
rect	166	56	167	57
rect	166	57	167	58
rect	166	59	167	60
rect	166	60	167	61
rect	166	62	167	63
rect	166	63	167	64
rect	166	65	167	66
rect	166	66	167	67
rect	166	68	167	69
rect	166	69	167	70
rect	166	71	167	72
rect	166	72	167	73
rect	166	74	167	75
rect	166	75	167	76
rect	166	77	167	78
rect	166	78	167	79
rect	166	80	167	81
rect	166	81	167	82
rect	166	83	167	84
rect	166	84	167	85
rect	166	86	167	87
rect	166	87	167	88
rect	166	89	167	90
rect	166	90	167	91
rect	166	92	167	93
rect	166	93	167	94
rect	166	95	167	96
rect	166	96	167	97
rect	166	98	167	99
rect	166	99	167	100
rect	166	101	167	102
rect	166	102	167	103
rect	166	104	167	105
rect	166	105	167	106
rect	166	107	167	108
rect	166	108	167	109
rect	166	110	167	111
rect	166	111	167	112
rect	166	113	167	114
rect	166	114	167	115
rect	166	116	167	117
rect	166	117	167	118
rect	166	119	167	120
rect	166	120	167	121
rect	166	122	167	123
rect	166	123	167	124
rect	166	125	167	126
rect	166	126	167	127
rect	166	128	167	129
rect	166	129	167	130
rect	166	131	167	132
rect	166	132	167	133
rect	166	134	167	135
rect	166	135	167	136
rect	166	137	167	138
rect	166	138	167	139
rect	166	140	167	141
rect	166	141	167	142
rect	166	143	167	144
rect	166	144	167	145
rect	166	146	167	147
rect	166	147	167	148
rect	166	149	167	150
rect	166	150	167	151
rect	166	152	167	153
rect	166	153	167	154
rect	166	155	167	156
rect	166	156	167	157
rect	166	158	167	159
rect	166	159	167	160
rect	166	161	167	162
rect	166	162	167	163
rect	166	164	167	165
rect	166	165	167	166
rect	166	167	167	168
rect	166	168	167	169
rect	166	170	167	171
rect	166	171	167	172
rect	166	173	167	174
rect	166	174	167	175
rect	166	176	167	177
rect	166	177	167	178
rect	166	179	167	180
rect	166	180	167	181
rect	166	182	167	183
rect	166	183	167	184
rect	166	185	167	186
rect	166	186	167	187
rect	166	188	167	189
rect	166	189	167	190
rect	166	191	167	192
rect	166	192	167	193
rect	166	194	167	195
rect	166	195	167	196
rect	166	197	167	198
rect	166	198	167	199
rect	166	200	167	201
rect	166	201	167	202
rect	166	203	167	204
rect	166	204	167	205
rect	166	206	167	207
rect	166	207	167	208
rect	166	209	167	210
rect	166	210	167	211
rect	166	212	167	213
rect	166	213	167	214
rect	166	215	167	216
rect	166	216	167	217
rect	166	218	167	219
rect	166	219	167	220
rect	166	221	167	222
rect	166	222	167	223
rect	166	224	167	225
rect	166	225	167	226
rect	166	227	167	228
rect	166	228	167	229
rect	166	230	167	231
rect	166	231	167	232
rect	166	233	167	234
rect	166	234	167	235
rect	166	236	167	237
rect	166	237	167	238
rect	166	239	167	240
rect	166	240	167	241
rect	166	242	167	243
rect	166	243	167	244
rect	166	245	167	246
rect	166	246	167	247
rect	166	248	167	249
rect	166	249	167	250
rect	166	251	167	252
rect	166	252	167	253
rect	166	254	167	255
rect	166	255	167	256
rect	166	257	167	258
rect	166	258	167	259
rect	166	260	167	261
rect	166	261	167	262
rect	166	263	167	264
rect	166	264	167	265
rect	166	266	167	267
rect	166	267	167	268
rect	166	269	167	270
rect	166	270	167	271
rect	166	272	167	273
rect	166	273	167	274
rect	166	275	167	276
rect	166	276	167	277
rect	166	278	167	279
rect	166	279	167	280
rect	166	281	167	282
rect	166	282	167	283
rect	166	284	167	285
rect	166	285	167	286
rect	166	287	167	288
rect	166	288	167	289
rect	166	290	167	291
rect	166	291	167	292
rect	166	293	167	294
rect	166	294	167	295
rect	166	296	167	297
rect	166	297	167	298
rect	166	299	167	300
rect	166	300	167	301
rect	166	302	167	303
rect	166	303	167	304
rect	166	304	167	305
rect	166	305	167	306
rect	166	306	167	307
rect	166	308	167	309
rect	166	309	167	310
rect	166	311	167	312
rect	166	312	167	313
rect	166	314	167	315
rect	166	315	167	316
rect	166	317	167	318
rect	166	318	167	319
rect	166	320	167	321
rect	166	321	167	322
rect	166	323	167	324
rect	166	324	167	325
rect	166	326	167	327
rect	166	327	167	328
rect	166	328	167	329
rect	166	329	167	330
rect	166	330	167	331
rect	166	332	167	333
rect	166	333	167	334
rect	166	335	167	336
rect	166	336	167	337
rect	166	337	167	338
rect	166	338	167	339
rect	166	339	167	340
rect	166	340	167	341
rect	166	341	167	342
rect	166	342	167	343
rect	166	343	167	344
rect	166	344	167	345
rect	166	345	167	346
rect	166	347	167	348
rect	166	348	167	349
rect	166	350	167	351
rect	166	351	167	352
rect	166	353	167	354
rect	166	354	167	355
rect	166	356	167	357
rect	166	357	167	358
rect	166	359	167	360
rect	166	360	167	361
rect	166	362	167	363
rect	166	363	167	364
rect	166	365	167	366
rect	166	366	167	367
rect	166	368	167	369
rect	173	0	174	1
rect	173	2	174	3
rect	173	3	174	4
rect	173	5	174	6
rect	173	6	174	7
rect	173	8	174	9
rect	173	9	174	10
rect	173	11	174	12
rect	173	12	174	13
rect	173	14	174	15
rect	173	15	174	16
rect	173	17	174	18
rect	173	18	174	19
rect	173	20	174	21
rect	173	21	174	22
rect	173	23	174	24
rect	173	24	174	25
rect	173	26	174	27
rect	173	27	174	28
rect	173	29	174	30
rect	173	30	174	31
rect	173	32	174	33
rect	173	33	174	34
rect	173	35	174	36
rect	173	36	174	37
rect	173	38	174	39
rect	173	39	174	40
rect	173	41	174	42
rect	173	42	174	43
rect	173	44	174	45
rect	173	45	174	46
rect	173	47	174	48
rect	173	48	174	49
rect	173	50	174	51
rect	173	51	174	52
rect	173	53	174	54
rect	173	54	174	55
rect	173	56	174	57
rect	173	57	174	58
rect	173	59	174	60
rect	173	60	174	61
rect	173	62	174	63
rect	173	63	174	64
rect	173	65	174	66
rect	173	66	174	67
rect	173	68	174	69
rect	173	69	174	70
rect	173	71	174	72
rect	173	72	174	73
rect	173	74	174	75
rect	173	75	174	76
rect	173	77	174	78
rect	173	78	174	79
rect	173	80	174	81
rect	173	81	174	82
rect	173	83	174	84
rect	173	84	174	85
rect	173	86	174	87
rect	173	87	174	88
rect	173	89	174	90
rect	173	90	174	91
rect	173	92	174	93
rect	173	93	174	94
rect	173	95	174	96
rect	173	96	174	97
rect	173	98	174	99
rect	173	99	174	100
rect	173	101	174	102
rect	173	102	174	103
rect	173	104	174	105
rect	173	105	174	106
rect	173	107	174	108
rect	173	108	174	109
rect	173	110	174	111
rect	173	111	174	112
rect	173	113	174	114
rect	173	114	174	115
rect	173	116	174	117
rect	173	117	174	118
rect	173	119	174	120
rect	173	120	174	121
rect	173	122	174	123
rect	173	123	174	124
rect	173	125	174	126
rect	173	126	174	127
rect	173	128	174	129
rect	173	129	174	130
rect	173	131	174	132
rect	173	132	174	133
rect	173	134	174	135
rect	173	135	174	136
rect	173	137	174	138
rect	173	138	174	139
rect	173	140	174	141
rect	173	141	174	142
rect	173	143	174	144
rect	173	144	174	145
rect	173	146	174	147
rect	173	147	174	148
rect	173	149	174	150
rect	173	150	174	151
rect	173	152	174	153
rect	173	153	174	154
rect	173	155	174	156
rect	173	156	174	157
rect	173	158	174	159
rect	173	159	174	160
rect	173	161	174	162
rect	173	162	174	163
rect	173	164	174	165
rect	173	165	174	166
rect	173	167	174	168
rect	173	168	174	169
rect	173	170	174	171
rect	173	171	174	172
rect	173	173	174	174
rect	173	174	174	175
rect	173	176	174	177
rect	173	177	174	178
rect	173	179	174	180
rect	173	180	174	181
rect	173	182	174	183
rect	173	183	174	184
rect	173	185	174	186
rect	173	186	174	187
rect	173	188	174	189
rect	173	189	174	190
rect	173	191	174	192
rect	173	192	174	193
rect	173	194	174	195
rect	173	195	174	196
rect	173	197	174	198
rect	173	198	174	199
rect	173	200	174	201
rect	173	201	174	202
rect	173	203	174	204
rect	173	204	174	205
rect	173	206	174	207
rect	173	207	174	208
rect	173	209	174	210
rect	173	210	174	211
rect	173	212	174	213
rect	173	213	174	214
rect	173	215	174	216
rect	173	216	174	217
rect	173	218	174	219
rect	173	219	174	220
rect	173	221	174	222
rect	173	222	174	223
rect	173	224	174	225
rect	173	225	174	226
rect	173	227	174	228
rect	173	228	174	229
rect	173	230	174	231
rect	173	231	174	232
rect	173	233	174	234
rect	173	234	174	235
rect	173	236	174	237
rect	173	237	174	238
rect	173	239	174	240
rect	173	240	174	241
rect	173	242	174	243
rect	173	243	174	244
rect	173	245	174	246
rect	173	246	174	247
rect	173	248	174	249
rect	173	249	174	250
rect	173	251	174	252
rect	173	252	174	253
rect	173	254	174	255
rect	173	255	174	256
rect	173	257	174	258
rect	173	258	174	259
rect	173	260	174	261
rect	173	261	174	262
rect	173	263	174	264
rect	173	264	174	265
rect	173	266	174	267
rect	173	267	174	268
rect	173	269	174	270
rect	173	270	174	271
rect	173	272	174	273
rect	173	273	174	274
rect	173	275	174	276
rect	173	276	174	277
rect	173	278	174	279
rect	173	279	174	280
rect	173	281	174	282
rect	173	282	174	283
rect	173	284	174	285
rect	173	285	174	286
rect	173	287	174	288
rect	173	288	174	289
rect	173	290	174	291
rect	173	291	174	292
rect	173	293	174	294
rect	173	294	174	295
rect	173	296	174	297
rect	173	297	174	298
rect	173	299	174	300
rect	173	300	174	301
rect	173	302	174	303
rect	173	303	174	304
rect	173	304	174	305
rect	173	305	174	306
rect	173	306	174	307
rect	173	308	174	309
rect	173	309	174	310
rect	173	311	174	312
rect	173	312	174	313
rect	173	314	174	315
rect	173	315	174	316
rect	173	317	174	318
rect	173	318	174	319
rect	173	319	174	320
rect	173	320	174	321
rect	173	321	174	322
rect	173	323	174	324
rect	173	324	174	325
rect	173	326	174	327
rect	173	327	174	328
rect	173	328	174	329
rect	173	329	174	330
rect	173	330	174	331
rect	173	332	174	333
rect	173	333	174	334
rect	173	335	174	336
rect	173	336	174	337
rect	173	337	174	338
rect	173	338	174	339
rect	173	339	174	340
rect	173	340	174	341
rect	173	341	174	342
rect	173	342	174	343
rect	173	343	174	344
rect	173	344	174	345
rect	173	345	174	346
rect	173	347	174	348
rect	173	348	174	349
rect	173	350	174	351
rect	173	351	174	352
rect	173	352	174	353
rect	173	353	174	354
rect	173	354	174	355
rect	173	356	174	357
rect	173	357	174	358
rect	173	358	174	359
rect	173	359	174	360
rect	173	360	174	361
rect	173	362	174	363
rect	173	363	174	364
rect	173	365	174	366
rect	173	366	174	367
rect	173	368	174	369
rect	175	0	176	1
rect	175	2	176	3
rect	175	3	176	4
rect	175	5	176	6
rect	175	6	176	7
rect	175	8	176	9
rect	175	9	176	10
rect	175	11	176	12
rect	175	12	176	13
rect	175	14	176	15
rect	175	15	176	16
rect	175	17	176	18
rect	175	18	176	19
rect	175	20	176	21
rect	175	21	176	22
rect	175	23	176	24
rect	175	24	176	25
rect	175	26	176	27
rect	175	27	176	28
rect	175	29	176	30
rect	175	30	176	31
rect	175	32	176	33
rect	175	33	176	34
rect	175	35	176	36
rect	175	36	176	37
rect	175	38	176	39
rect	175	39	176	40
rect	175	41	176	42
rect	175	42	176	43
rect	175	44	176	45
rect	175	45	176	46
rect	175	47	176	48
rect	175	48	176	49
rect	175	50	176	51
rect	175	51	176	52
rect	175	53	176	54
rect	175	54	176	55
rect	175	56	176	57
rect	175	57	176	58
rect	175	59	176	60
rect	175	60	176	61
rect	175	62	176	63
rect	175	63	176	64
rect	175	65	176	66
rect	175	66	176	67
rect	175	68	176	69
rect	175	69	176	70
rect	175	71	176	72
rect	175	72	176	73
rect	175	74	176	75
rect	175	75	176	76
rect	175	77	176	78
rect	175	78	176	79
rect	175	80	176	81
rect	175	81	176	82
rect	175	83	176	84
rect	175	84	176	85
rect	175	86	176	87
rect	175	87	176	88
rect	175	89	176	90
rect	175	90	176	91
rect	175	92	176	93
rect	175	93	176	94
rect	175	95	176	96
rect	175	96	176	97
rect	175	98	176	99
rect	175	99	176	100
rect	175	101	176	102
rect	175	102	176	103
rect	175	104	176	105
rect	175	105	176	106
rect	175	107	176	108
rect	175	108	176	109
rect	175	110	176	111
rect	175	111	176	112
rect	175	113	176	114
rect	175	114	176	115
rect	175	116	176	117
rect	175	117	176	118
rect	175	119	176	120
rect	175	120	176	121
rect	175	122	176	123
rect	175	123	176	124
rect	175	125	176	126
rect	175	126	176	127
rect	175	128	176	129
rect	175	129	176	130
rect	175	131	176	132
rect	175	132	176	133
rect	175	134	176	135
rect	175	135	176	136
rect	175	137	176	138
rect	175	138	176	139
rect	175	140	176	141
rect	175	141	176	142
rect	175	143	176	144
rect	175	144	176	145
rect	175	146	176	147
rect	175	147	176	148
rect	175	149	176	150
rect	175	150	176	151
rect	175	152	176	153
rect	175	153	176	154
rect	175	155	176	156
rect	175	156	176	157
rect	175	158	176	159
rect	175	159	176	160
rect	175	161	176	162
rect	175	162	176	163
rect	175	164	176	165
rect	175	165	176	166
rect	175	167	176	168
rect	175	168	176	169
rect	175	170	176	171
rect	175	171	176	172
rect	175	173	176	174
rect	175	174	176	175
rect	175	176	176	177
rect	175	177	176	178
rect	175	179	176	180
rect	175	180	176	181
rect	175	182	176	183
rect	175	183	176	184
rect	175	185	176	186
rect	175	186	176	187
rect	175	188	176	189
rect	175	189	176	190
rect	175	191	176	192
rect	175	192	176	193
rect	175	194	176	195
rect	175	195	176	196
rect	175	197	176	198
rect	175	198	176	199
rect	175	200	176	201
rect	175	201	176	202
rect	175	203	176	204
rect	175	204	176	205
rect	175	206	176	207
rect	175	207	176	208
rect	175	209	176	210
rect	175	210	176	211
rect	175	212	176	213
rect	175	213	176	214
rect	175	215	176	216
rect	175	216	176	217
rect	175	218	176	219
rect	175	219	176	220
rect	175	221	176	222
rect	175	222	176	223
rect	175	224	176	225
rect	175	225	176	226
rect	175	227	176	228
rect	175	228	176	229
rect	175	230	176	231
rect	175	231	176	232
rect	175	233	176	234
rect	175	234	176	235
rect	175	236	176	237
rect	175	237	176	238
rect	175	239	176	240
rect	175	240	176	241
rect	175	242	176	243
rect	175	243	176	244
rect	175	245	176	246
rect	175	246	176	247
rect	175	248	176	249
rect	175	249	176	250
rect	175	251	176	252
rect	175	252	176	253
rect	175	254	176	255
rect	175	255	176	256
rect	175	257	176	258
rect	175	258	176	259
rect	175	260	176	261
rect	175	261	176	262
rect	175	263	176	264
rect	175	264	176	265
rect	175	266	176	267
rect	175	267	176	268
rect	175	269	176	270
rect	175	270	176	271
rect	175	272	176	273
rect	175	273	176	274
rect	175	275	176	276
rect	175	276	176	277
rect	175	278	176	279
rect	175	279	176	280
rect	175	281	176	282
rect	175	282	176	283
rect	175	284	176	285
rect	175	285	176	286
rect	175	287	176	288
rect	175	288	176	289
rect	175	290	176	291
rect	175	291	176	292
rect	175	293	176	294
rect	175	294	176	295
rect	175	296	176	297
rect	175	297	176	298
rect	175	299	176	300
rect	175	300	176	301
rect	175	302	176	303
rect	175	303	176	304
rect	175	304	176	305
rect	175	305	176	306
rect	175	306	176	307
rect	175	308	176	309
rect	175	309	176	310
rect	175	311	176	312
rect	175	312	176	313
rect	175	314	176	315
rect	175	315	176	316
rect	175	317	176	318
rect	175	318	176	319
rect	175	319	176	320
rect	175	320	176	321
rect	175	321	176	322
rect	175	323	176	324
rect	175	324	176	325
rect	175	326	176	327
rect	175	327	176	328
rect	175	328	176	329
rect	175	329	176	330
rect	175	330	176	331
rect	175	332	176	333
rect	175	333	176	334
rect	175	335	176	336
rect	175	336	176	337
rect	175	337	176	338
rect	175	338	176	339
rect	175	339	176	340
rect	175	340	176	341
rect	175	341	176	342
rect	175	342	176	343
rect	175	343	176	344
rect	175	344	176	345
rect	175	345	176	346
rect	175	347	176	348
rect	175	348	176	349
rect	175	350	176	351
rect	175	351	176	352
rect	175	352	176	353
rect	175	353	176	354
rect	175	354	176	355
rect	175	356	176	357
rect	175	357	176	358
rect	175	358	176	359
rect	175	359	176	360
rect	175	360	176	361
rect	175	362	176	363
rect	175	363	176	364
rect	175	365	176	366
rect	175	366	176	367
rect	175	368	176	369
rect	176	0	177	1
rect	176	2	177	3
rect	176	3	177	4
rect	176	5	177	6
rect	176	6	177	7
rect	176	8	177	9
rect	176	9	177	10
rect	176	11	177	12
rect	176	12	177	13
rect	176	14	177	15
rect	176	15	177	16
rect	176	17	177	18
rect	176	18	177	19
rect	176	20	177	21
rect	176	21	177	22
rect	176	23	177	24
rect	176	24	177	25
rect	176	26	177	27
rect	176	27	177	28
rect	176	29	177	30
rect	176	30	177	31
rect	176	32	177	33
rect	176	33	177	34
rect	176	35	177	36
rect	176	36	177	37
rect	176	38	177	39
rect	176	39	177	40
rect	176	41	177	42
rect	176	42	177	43
rect	176	44	177	45
rect	176	45	177	46
rect	176	47	177	48
rect	176	48	177	49
rect	176	50	177	51
rect	176	51	177	52
rect	176	53	177	54
rect	176	54	177	55
rect	176	56	177	57
rect	176	57	177	58
rect	176	59	177	60
rect	176	60	177	61
rect	176	62	177	63
rect	176	63	177	64
rect	176	65	177	66
rect	176	66	177	67
rect	176	68	177	69
rect	176	69	177	70
rect	176	71	177	72
rect	176	72	177	73
rect	176	74	177	75
rect	176	75	177	76
rect	176	77	177	78
rect	176	78	177	79
rect	176	80	177	81
rect	176	81	177	82
rect	176	83	177	84
rect	176	84	177	85
rect	176	86	177	87
rect	176	87	177	88
rect	176	89	177	90
rect	176	90	177	91
rect	176	92	177	93
rect	176	93	177	94
rect	176	95	177	96
rect	176	96	177	97
rect	176	98	177	99
rect	176	99	177	100
rect	176	101	177	102
rect	176	102	177	103
rect	176	104	177	105
rect	176	105	177	106
rect	176	107	177	108
rect	176	108	177	109
rect	176	110	177	111
rect	176	111	177	112
rect	176	113	177	114
rect	176	114	177	115
rect	176	116	177	117
rect	176	117	177	118
rect	176	119	177	120
rect	176	120	177	121
rect	176	122	177	123
rect	176	123	177	124
rect	176	125	177	126
rect	176	126	177	127
rect	176	128	177	129
rect	176	129	177	130
rect	176	131	177	132
rect	176	132	177	133
rect	176	134	177	135
rect	176	135	177	136
rect	176	137	177	138
rect	176	138	177	139
rect	176	140	177	141
rect	176	141	177	142
rect	176	143	177	144
rect	176	144	177	145
rect	176	146	177	147
rect	176	147	177	148
rect	176	149	177	150
rect	176	150	177	151
rect	176	152	177	153
rect	176	153	177	154
rect	176	155	177	156
rect	176	156	177	157
rect	176	158	177	159
rect	176	159	177	160
rect	176	161	177	162
rect	176	162	177	163
rect	176	164	177	165
rect	176	165	177	166
rect	176	167	177	168
rect	176	168	177	169
rect	176	170	177	171
rect	176	171	177	172
rect	176	173	177	174
rect	176	174	177	175
rect	176	176	177	177
rect	176	177	177	178
rect	176	179	177	180
rect	176	180	177	181
rect	176	182	177	183
rect	176	183	177	184
rect	176	185	177	186
rect	176	186	177	187
rect	176	188	177	189
rect	176	189	177	190
rect	176	191	177	192
rect	176	192	177	193
rect	176	194	177	195
rect	176	195	177	196
rect	176	197	177	198
rect	176	198	177	199
rect	176	200	177	201
rect	176	201	177	202
rect	176	203	177	204
rect	176	204	177	205
rect	176	206	177	207
rect	176	207	177	208
rect	176	209	177	210
rect	176	210	177	211
rect	176	212	177	213
rect	176	213	177	214
rect	176	215	177	216
rect	176	216	177	217
rect	176	218	177	219
rect	176	219	177	220
rect	176	221	177	222
rect	176	222	177	223
rect	176	224	177	225
rect	176	225	177	226
rect	176	227	177	228
rect	176	228	177	229
rect	176	230	177	231
rect	176	231	177	232
rect	176	233	177	234
rect	176	234	177	235
rect	176	236	177	237
rect	176	237	177	238
rect	176	239	177	240
rect	176	240	177	241
rect	176	242	177	243
rect	176	243	177	244
rect	176	245	177	246
rect	176	246	177	247
rect	176	248	177	249
rect	176	249	177	250
rect	176	251	177	252
rect	176	252	177	253
rect	176	254	177	255
rect	176	255	177	256
rect	176	257	177	258
rect	176	258	177	259
rect	176	260	177	261
rect	176	261	177	262
rect	176	263	177	264
rect	176	264	177	265
rect	176	266	177	267
rect	176	267	177	268
rect	176	269	177	270
rect	176	270	177	271
rect	176	272	177	273
rect	176	273	177	274
rect	176	275	177	276
rect	176	276	177	277
rect	176	278	177	279
rect	176	279	177	280
rect	176	281	177	282
rect	176	282	177	283
rect	176	284	177	285
rect	176	285	177	286
rect	176	287	177	288
rect	176	288	177	289
rect	176	290	177	291
rect	176	291	177	292
rect	176	293	177	294
rect	176	294	177	295
rect	176	296	177	297
rect	176	297	177	298
rect	176	299	177	300
rect	176	300	177	301
rect	176	302	177	303
rect	176	303	177	304
rect	176	304	177	305
rect	176	305	177	306
rect	176	306	177	307
rect	176	308	177	309
rect	176	309	177	310
rect	176	311	177	312
rect	176	312	177	313
rect	176	314	177	315
rect	176	315	177	316
rect	176	317	177	318
rect	176	318	177	319
rect	176	319	177	320
rect	176	320	177	321
rect	176	321	177	322
rect	176	323	177	324
rect	176	324	177	325
rect	176	326	177	327
rect	176	327	177	328
rect	176	328	177	329
rect	176	329	177	330
rect	176	330	177	331
rect	176	332	177	333
rect	176	333	177	334
rect	176	335	177	336
rect	176	336	177	337
rect	176	337	177	338
rect	176	338	177	339
rect	176	339	177	340
rect	176	340	177	341
rect	176	341	177	342
rect	176	342	177	343
rect	176	343	177	344
rect	176	344	177	345
rect	176	345	177	346
rect	176	347	177	348
rect	176	348	177	349
rect	176	350	177	351
rect	176	351	177	352
rect	176	352	177	353
rect	176	353	177	354
rect	176	354	177	355
rect	176	356	177	357
rect	176	357	177	358
rect	176	358	177	359
rect	176	359	177	360
rect	176	360	177	361
rect	176	362	177	363
rect	176	363	177	364
rect	176	365	177	366
rect	176	366	177	367
rect	176	368	177	369
rect	177	0	178	1
rect	177	2	178	3
rect	177	3	178	4
rect	177	5	178	6
rect	177	6	178	7
rect	177	8	178	9
rect	177	9	178	10
rect	177	11	178	12
rect	177	12	178	13
rect	177	14	178	15
rect	177	15	178	16
rect	177	17	178	18
rect	177	18	178	19
rect	177	20	178	21
rect	177	21	178	22
rect	177	23	178	24
rect	177	24	178	25
rect	177	26	178	27
rect	177	27	178	28
rect	177	29	178	30
rect	177	30	178	31
rect	177	32	178	33
rect	177	33	178	34
rect	177	35	178	36
rect	177	36	178	37
rect	177	38	178	39
rect	177	39	178	40
rect	177	41	178	42
rect	177	42	178	43
rect	177	44	178	45
rect	177	45	178	46
rect	177	47	178	48
rect	177	48	178	49
rect	177	50	178	51
rect	177	51	178	52
rect	177	53	178	54
rect	177	54	178	55
rect	177	56	178	57
rect	177	57	178	58
rect	177	59	178	60
rect	177	60	178	61
rect	177	62	178	63
rect	177	63	178	64
rect	177	65	178	66
rect	177	66	178	67
rect	177	68	178	69
rect	177	69	178	70
rect	177	71	178	72
rect	177	72	178	73
rect	177	74	178	75
rect	177	75	178	76
rect	177	77	178	78
rect	177	78	178	79
rect	177	80	178	81
rect	177	81	178	82
rect	177	83	178	84
rect	177	84	178	85
rect	177	86	178	87
rect	177	87	178	88
rect	177	89	178	90
rect	177	90	178	91
rect	177	92	178	93
rect	177	93	178	94
rect	177	95	178	96
rect	177	96	178	97
rect	177	98	178	99
rect	177	99	178	100
rect	177	101	178	102
rect	177	102	178	103
rect	177	104	178	105
rect	177	105	178	106
rect	177	107	178	108
rect	177	108	178	109
rect	177	110	178	111
rect	177	111	178	112
rect	177	113	178	114
rect	177	114	178	115
rect	177	116	178	117
rect	177	117	178	118
rect	177	119	178	120
rect	177	120	178	121
rect	177	122	178	123
rect	177	123	178	124
rect	177	125	178	126
rect	177	126	178	127
rect	177	128	178	129
rect	177	129	178	130
rect	177	131	178	132
rect	177	132	178	133
rect	177	134	178	135
rect	177	135	178	136
rect	177	137	178	138
rect	177	138	178	139
rect	177	140	178	141
rect	177	141	178	142
rect	177	143	178	144
rect	177	144	178	145
rect	177	146	178	147
rect	177	147	178	148
rect	177	149	178	150
rect	177	150	178	151
rect	177	152	178	153
rect	177	153	178	154
rect	177	155	178	156
rect	177	156	178	157
rect	177	158	178	159
rect	177	159	178	160
rect	177	161	178	162
rect	177	162	178	163
rect	177	164	178	165
rect	177	165	178	166
rect	177	167	178	168
rect	177	168	178	169
rect	177	170	178	171
rect	177	171	178	172
rect	177	173	178	174
rect	177	174	178	175
rect	177	176	178	177
rect	177	177	178	178
rect	177	179	178	180
rect	177	180	178	181
rect	177	182	178	183
rect	177	183	178	184
rect	177	185	178	186
rect	177	186	178	187
rect	177	188	178	189
rect	177	189	178	190
rect	177	191	178	192
rect	177	192	178	193
rect	177	194	178	195
rect	177	195	178	196
rect	177	197	178	198
rect	177	198	178	199
rect	177	200	178	201
rect	177	201	178	202
rect	177	203	178	204
rect	177	204	178	205
rect	177	206	178	207
rect	177	207	178	208
rect	177	209	178	210
rect	177	210	178	211
rect	177	212	178	213
rect	177	213	178	214
rect	177	215	178	216
rect	177	216	178	217
rect	177	218	178	219
rect	177	219	178	220
rect	177	221	178	222
rect	177	222	178	223
rect	177	224	178	225
rect	177	225	178	226
rect	177	227	178	228
rect	177	228	178	229
rect	177	230	178	231
rect	177	231	178	232
rect	177	233	178	234
rect	177	234	178	235
rect	177	236	178	237
rect	177	237	178	238
rect	177	239	178	240
rect	177	240	178	241
rect	177	242	178	243
rect	177	243	178	244
rect	177	245	178	246
rect	177	246	178	247
rect	177	248	178	249
rect	177	249	178	250
rect	177	251	178	252
rect	177	252	178	253
rect	177	254	178	255
rect	177	255	178	256
rect	177	257	178	258
rect	177	258	178	259
rect	177	260	178	261
rect	177	261	178	262
rect	177	263	178	264
rect	177	264	178	265
rect	177	266	178	267
rect	177	267	178	268
rect	177	269	178	270
rect	177	270	178	271
rect	177	272	178	273
rect	177	273	178	274
rect	177	275	178	276
rect	177	276	178	277
rect	177	278	178	279
rect	177	279	178	280
rect	177	281	178	282
rect	177	282	178	283
rect	177	284	178	285
rect	177	285	178	286
rect	177	287	178	288
rect	177	288	178	289
rect	177	290	178	291
rect	177	291	178	292
rect	177	293	178	294
rect	177	294	178	295
rect	177	296	178	297
rect	177	297	178	298
rect	177	299	178	300
rect	177	300	178	301
rect	177	302	178	303
rect	177	303	178	304
rect	177	304	178	305
rect	177	305	178	306
rect	177	306	178	307
rect	177	308	178	309
rect	177	309	178	310
rect	177	311	178	312
rect	177	312	178	313
rect	177	314	178	315
rect	177	315	178	316
rect	177	317	178	318
rect	177	318	178	319
rect	177	319	178	320
rect	177	320	178	321
rect	177	321	178	322
rect	177	323	178	324
rect	177	324	178	325
rect	177	326	178	327
rect	177	327	178	328
rect	177	328	178	329
rect	177	329	178	330
rect	177	330	178	331
rect	177	332	178	333
rect	177	333	178	334
rect	177	335	178	336
rect	177	336	178	337
rect	177	337	178	338
rect	177	338	178	339
rect	177	339	178	340
rect	177	340	178	341
rect	177	341	178	342
rect	177	342	178	343
rect	177	343	178	344
rect	177	344	178	345
rect	177	345	178	346
rect	177	347	178	348
rect	177	348	178	349
rect	177	350	178	351
rect	177	351	178	352
rect	177	352	178	353
rect	177	353	178	354
rect	177	354	178	355
rect	177	356	178	357
rect	177	357	178	358
rect	177	358	178	359
rect	177	359	178	360
rect	177	360	178	361
rect	177	362	178	363
rect	177	363	178	364
rect	177	365	178	366
rect	177	366	178	367
rect	177	368	178	369
rect	178	0	179	1
rect	178	2	179	3
rect	178	3	179	4
rect	178	5	179	6
rect	178	6	179	7
rect	178	8	179	9
rect	178	9	179	10
rect	178	11	179	12
rect	178	12	179	13
rect	178	14	179	15
rect	178	15	179	16
rect	178	17	179	18
rect	178	18	179	19
rect	178	20	179	21
rect	178	21	179	22
rect	178	23	179	24
rect	178	24	179	25
rect	178	26	179	27
rect	178	27	179	28
rect	178	29	179	30
rect	178	30	179	31
rect	178	32	179	33
rect	178	33	179	34
rect	178	35	179	36
rect	178	36	179	37
rect	178	38	179	39
rect	178	39	179	40
rect	178	41	179	42
rect	178	42	179	43
rect	178	44	179	45
rect	178	45	179	46
rect	178	47	179	48
rect	178	48	179	49
rect	178	50	179	51
rect	178	51	179	52
rect	178	53	179	54
rect	178	54	179	55
rect	178	56	179	57
rect	178	57	179	58
rect	178	59	179	60
rect	178	60	179	61
rect	178	62	179	63
rect	178	63	179	64
rect	178	65	179	66
rect	178	66	179	67
rect	178	68	179	69
rect	178	69	179	70
rect	178	71	179	72
rect	178	72	179	73
rect	178	74	179	75
rect	178	75	179	76
rect	178	77	179	78
rect	178	78	179	79
rect	178	80	179	81
rect	178	81	179	82
rect	178	83	179	84
rect	178	84	179	85
rect	178	86	179	87
rect	178	87	179	88
rect	178	89	179	90
rect	178	90	179	91
rect	178	92	179	93
rect	178	93	179	94
rect	178	95	179	96
rect	178	96	179	97
rect	178	98	179	99
rect	178	99	179	100
rect	178	101	179	102
rect	178	102	179	103
rect	178	104	179	105
rect	178	105	179	106
rect	178	107	179	108
rect	178	108	179	109
rect	178	110	179	111
rect	178	111	179	112
rect	178	113	179	114
rect	178	114	179	115
rect	178	116	179	117
rect	178	117	179	118
rect	178	119	179	120
rect	178	120	179	121
rect	178	122	179	123
rect	178	123	179	124
rect	178	125	179	126
rect	178	126	179	127
rect	178	128	179	129
rect	178	129	179	130
rect	178	131	179	132
rect	178	132	179	133
rect	178	134	179	135
rect	178	135	179	136
rect	178	137	179	138
rect	178	138	179	139
rect	178	140	179	141
rect	178	141	179	142
rect	178	143	179	144
rect	178	144	179	145
rect	178	146	179	147
rect	178	147	179	148
rect	178	149	179	150
rect	178	150	179	151
rect	178	152	179	153
rect	178	153	179	154
rect	178	155	179	156
rect	178	156	179	157
rect	178	158	179	159
rect	178	159	179	160
rect	178	161	179	162
rect	178	162	179	163
rect	178	164	179	165
rect	178	165	179	166
rect	178	167	179	168
rect	178	168	179	169
rect	178	170	179	171
rect	178	171	179	172
rect	178	173	179	174
rect	178	174	179	175
rect	178	176	179	177
rect	178	177	179	178
rect	178	179	179	180
rect	178	180	179	181
rect	178	182	179	183
rect	178	183	179	184
rect	178	185	179	186
rect	178	186	179	187
rect	178	188	179	189
rect	178	189	179	190
rect	178	191	179	192
rect	178	192	179	193
rect	178	194	179	195
rect	178	195	179	196
rect	178	197	179	198
rect	178	198	179	199
rect	178	200	179	201
rect	178	201	179	202
rect	178	203	179	204
rect	178	204	179	205
rect	178	206	179	207
rect	178	207	179	208
rect	178	209	179	210
rect	178	210	179	211
rect	178	212	179	213
rect	178	213	179	214
rect	178	215	179	216
rect	178	216	179	217
rect	178	218	179	219
rect	178	219	179	220
rect	178	221	179	222
rect	178	222	179	223
rect	178	224	179	225
rect	178	225	179	226
rect	178	227	179	228
rect	178	228	179	229
rect	178	230	179	231
rect	178	231	179	232
rect	178	233	179	234
rect	178	234	179	235
rect	178	236	179	237
rect	178	237	179	238
rect	178	239	179	240
rect	178	240	179	241
rect	178	242	179	243
rect	178	243	179	244
rect	178	245	179	246
rect	178	246	179	247
rect	178	248	179	249
rect	178	249	179	250
rect	178	251	179	252
rect	178	252	179	253
rect	178	254	179	255
rect	178	255	179	256
rect	178	257	179	258
rect	178	258	179	259
rect	178	260	179	261
rect	178	261	179	262
rect	178	263	179	264
rect	178	264	179	265
rect	178	266	179	267
rect	178	267	179	268
rect	178	269	179	270
rect	178	270	179	271
rect	178	272	179	273
rect	178	273	179	274
rect	178	275	179	276
rect	178	276	179	277
rect	178	278	179	279
rect	178	279	179	280
rect	178	281	179	282
rect	178	282	179	283
rect	178	284	179	285
rect	178	285	179	286
rect	178	287	179	288
rect	178	288	179	289
rect	178	290	179	291
rect	178	291	179	292
rect	178	293	179	294
rect	178	294	179	295
rect	178	296	179	297
rect	178	297	179	298
rect	178	299	179	300
rect	178	300	179	301
rect	178	302	179	303
rect	178	303	179	304
rect	178	304	179	305
rect	178	305	179	306
rect	178	306	179	307
rect	178	308	179	309
rect	178	309	179	310
rect	178	311	179	312
rect	178	312	179	313
rect	178	314	179	315
rect	178	315	179	316
rect	178	317	179	318
rect	178	318	179	319
rect	178	319	179	320
rect	178	320	179	321
rect	178	321	179	322
rect	178	323	179	324
rect	178	324	179	325
rect	178	326	179	327
rect	178	327	179	328
rect	178	328	179	329
rect	178	329	179	330
rect	178	330	179	331
rect	178	332	179	333
rect	178	333	179	334
rect	178	335	179	336
rect	178	336	179	337
rect	178	337	179	338
rect	178	338	179	339
rect	178	339	179	340
rect	178	340	179	341
rect	178	341	179	342
rect	178	342	179	343
rect	178	343	179	344
rect	178	344	179	345
rect	178	345	179	346
rect	178	347	179	348
rect	178	348	179	349
rect	178	350	179	351
rect	178	351	179	352
rect	178	352	179	353
rect	178	353	179	354
rect	178	354	179	355
rect	178	356	179	357
rect	178	357	179	358
rect	178	358	179	359
rect	178	359	179	360
rect	178	360	179	361
rect	178	362	179	363
rect	178	363	179	364
rect	178	365	179	366
rect	178	366	179	367
rect	178	368	179	369
rect	179	0	180	1
rect	179	2	180	3
rect	179	3	180	4
rect	179	5	180	6
rect	179	6	180	7
rect	179	8	180	9
rect	179	9	180	10
rect	179	11	180	12
rect	179	12	180	13
rect	179	14	180	15
rect	179	15	180	16
rect	179	17	180	18
rect	179	18	180	19
rect	179	20	180	21
rect	179	21	180	22
rect	179	23	180	24
rect	179	24	180	25
rect	179	26	180	27
rect	179	27	180	28
rect	179	29	180	30
rect	179	30	180	31
rect	179	32	180	33
rect	179	33	180	34
rect	179	35	180	36
rect	179	36	180	37
rect	179	38	180	39
rect	179	39	180	40
rect	179	41	180	42
rect	179	42	180	43
rect	179	44	180	45
rect	179	45	180	46
rect	179	47	180	48
rect	179	48	180	49
rect	179	50	180	51
rect	179	51	180	52
rect	179	53	180	54
rect	179	54	180	55
rect	179	56	180	57
rect	179	57	180	58
rect	179	59	180	60
rect	179	60	180	61
rect	179	62	180	63
rect	179	63	180	64
rect	179	65	180	66
rect	179	66	180	67
rect	179	68	180	69
rect	179	69	180	70
rect	179	71	180	72
rect	179	72	180	73
rect	179	74	180	75
rect	179	75	180	76
rect	179	77	180	78
rect	179	78	180	79
rect	179	80	180	81
rect	179	81	180	82
rect	179	83	180	84
rect	179	84	180	85
rect	179	86	180	87
rect	179	87	180	88
rect	179	89	180	90
rect	179	90	180	91
rect	179	92	180	93
rect	179	93	180	94
rect	179	95	180	96
rect	179	96	180	97
rect	179	98	180	99
rect	179	99	180	100
rect	179	101	180	102
rect	179	102	180	103
rect	179	104	180	105
rect	179	105	180	106
rect	179	107	180	108
rect	179	108	180	109
rect	179	110	180	111
rect	179	111	180	112
rect	179	113	180	114
rect	179	114	180	115
rect	179	116	180	117
rect	179	117	180	118
rect	179	119	180	120
rect	179	120	180	121
rect	179	122	180	123
rect	179	123	180	124
rect	179	125	180	126
rect	179	126	180	127
rect	179	128	180	129
rect	179	129	180	130
rect	179	131	180	132
rect	179	132	180	133
rect	179	134	180	135
rect	179	135	180	136
rect	179	137	180	138
rect	179	138	180	139
rect	179	140	180	141
rect	179	141	180	142
rect	179	143	180	144
rect	179	144	180	145
rect	179	146	180	147
rect	179	147	180	148
rect	179	149	180	150
rect	179	150	180	151
rect	179	152	180	153
rect	179	153	180	154
rect	179	155	180	156
rect	179	156	180	157
rect	179	158	180	159
rect	179	159	180	160
rect	179	161	180	162
rect	179	162	180	163
rect	179	164	180	165
rect	179	165	180	166
rect	179	167	180	168
rect	179	168	180	169
rect	179	170	180	171
rect	179	171	180	172
rect	179	173	180	174
rect	179	174	180	175
rect	179	176	180	177
rect	179	177	180	178
rect	179	179	180	180
rect	179	180	180	181
rect	179	182	180	183
rect	179	183	180	184
rect	179	185	180	186
rect	179	186	180	187
rect	179	188	180	189
rect	179	189	180	190
rect	179	191	180	192
rect	179	192	180	193
rect	179	194	180	195
rect	179	195	180	196
rect	179	197	180	198
rect	179	198	180	199
rect	179	200	180	201
rect	179	201	180	202
rect	179	203	180	204
rect	179	204	180	205
rect	179	206	180	207
rect	179	207	180	208
rect	179	209	180	210
rect	179	210	180	211
rect	179	212	180	213
rect	179	213	180	214
rect	179	215	180	216
rect	179	216	180	217
rect	179	218	180	219
rect	179	219	180	220
rect	179	221	180	222
rect	179	222	180	223
rect	179	224	180	225
rect	179	225	180	226
rect	179	227	180	228
rect	179	228	180	229
rect	179	230	180	231
rect	179	231	180	232
rect	179	233	180	234
rect	179	234	180	235
rect	179	236	180	237
rect	179	237	180	238
rect	179	239	180	240
rect	179	240	180	241
rect	179	242	180	243
rect	179	243	180	244
rect	179	245	180	246
rect	179	246	180	247
rect	179	248	180	249
rect	179	249	180	250
rect	179	251	180	252
rect	179	252	180	253
rect	179	254	180	255
rect	179	255	180	256
rect	179	257	180	258
rect	179	258	180	259
rect	179	260	180	261
rect	179	261	180	262
rect	179	263	180	264
rect	179	264	180	265
rect	179	266	180	267
rect	179	267	180	268
rect	179	269	180	270
rect	179	270	180	271
rect	179	272	180	273
rect	179	273	180	274
rect	179	275	180	276
rect	179	276	180	277
rect	179	278	180	279
rect	179	279	180	280
rect	179	281	180	282
rect	179	282	180	283
rect	179	284	180	285
rect	179	285	180	286
rect	179	287	180	288
rect	179	288	180	289
rect	179	290	180	291
rect	179	291	180	292
rect	179	293	180	294
rect	179	294	180	295
rect	179	296	180	297
rect	179	297	180	298
rect	179	299	180	300
rect	179	300	180	301
rect	179	302	180	303
rect	179	303	180	304
rect	179	304	180	305
rect	179	305	180	306
rect	179	306	180	307
rect	179	308	180	309
rect	179	309	180	310
rect	179	311	180	312
rect	179	312	180	313
rect	179	314	180	315
rect	179	315	180	316
rect	179	317	180	318
rect	179	318	180	319
rect	179	319	180	320
rect	179	320	180	321
rect	179	321	180	322
rect	179	323	180	324
rect	179	324	180	325
rect	179	326	180	327
rect	179	327	180	328
rect	179	328	180	329
rect	179	329	180	330
rect	179	330	180	331
rect	179	332	180	333
rect	179	333	180	334
rect	179	335	180	336
rect	179	336	180	337
rect	179	337	180	338
rect	179	338	180	339
rect	179	339	180	340
rect	179	340	180	341
rect	179	341	180	342
rect	179	342	180	343
rect	179	343	180	344
rect	179	344	180	345
rect	179	345	180	346
rect	179	347	180	348
rect	179	348	180	349
rect	179	350	180	351
rect	179	351	180	352
rect	179	352	180	353
rect	179	353	180	354
rect	179	354	180	355
rect	179	356	180	357
rect	179	357	180	358
rect	179	358	180	359
rect	179	359	180	360
rect	179	360	180	361
rect	179	362	180	363
rect	179	363	180	364
rect	179	365	180	366
rect	179	366	180	367
rect	179	368	180	369
rect	192	0	193	1
rect	192	1	193	2
rect	192	2	193	3
rect	192	3	193	4
rect	192	5	193	6
rect	192	6	193	7
rect	192	8	193	9
rect	192	9	193	10
rect	192	11	193	12
rect	192	12	193	13
rect	192	14	193	15
rect	192	15	193	16
rect	192	17	193	18
rect	192	18	193	19
rect	192	20	193	21
rect	192	21	193	22
rect	192	23	193	24
rect	192	24	193	25
rect	192	26	193	27
rect	192	27	193	28
rect	192	29	193	30
rect	192	30	193	31
rect	192	32	193	33
rect	192	33	193	34
rect	192	35	193	36
rect	192	36	193	37
rect	192	38	193	39
rect	192	39	193	40
rect	192	41	193	42
rect	192	42	193	43
rect	192	44	193	45
rect	192	45	193	46
rect	192	47	193	48
rect	192	48	193	49
rect	192	50	193	51
rect	192	51	193	52
rect	192	53	193	54
rect	192	54	193	55
rect	192	56	193	57
rect	192	57	193	58
rect	192	59	193	60
rect	192	60	193	61
rect	192	62	193	63
rect	192	63	193	64
rect	192	65	193	66
rect	192	66	193	67
rect	192	68	193	69
rect	192	69	193	70
rect	192	71	193	72
rect	192	72	193	73
rect	192	74	193	75
rect	192	75	193	76
rect	192	77	193	78
rect	192	78	193	79
rect	192	80	193	81
rect	192	81	193	82
rect	192	83	193	84
rect	192	84	193	85
rect	192	86	193	87
rect	192	87	193	88
rect	192	89	193	90
rect	192	90	193	91
rect	192	92	193	93
rect	192	93	193	94
rect	192	95	193	96
rect	192	96	193	97
rect	192	98	193	99
rect	192	99	193	100
rect	192	101	193	102
rect	192	102	193	103
rect	192	104	193	105
rect	192	105	193	106
rect	192	107	193	108
rect	192	108	193	109
rect	192	110	193	111
rect	192	111	193	112
rect	192	113	193	114
rect	192	114	193	115
rect	192	116	193	117
rect	192	117	193	118
rect	192	119	193	120
rect	192	120	193	121
rect	192	122	193	123
rect	192	123	193	124
rect	192	125	193	126
rect	192	126	193	127
rect	192	128	193	129
rect	192	129	193	130
rect	192	131	193	132
rect	192	132	193	133
rect	192	134	193	135
rect	192	135	193	136
rect	192	137	193	138
rect	192	138	193	139
rect	192	140	193	141
rect	192	141	193	142
rect	192	143	193	144
rect	192	144	193	145
rect	192	146	193	147
rect	192	147	193	148
rect	192	149	193	150
rect	192	150	193	151
rect	192	152	193	153
rect	192	153	193	154
rect	192	155	193	156
rect	192	156	193	157
rect	192	158	193	159
rect	192	159	193	160
rect	192	161	193	162
rect	192	162	193	163
rect	192	164	193	165
rect	192	165	193	166
rect	192	167	193	168
rect	192	168	193	169
rect	192	170	193	171
rect	192	171	193	172
rect	192	173	193	174
rect	192	174	193	175
rect	192	176	193	177
rect	192	177	193	178
rect	192	179	193	180
rect	192	180	193	181
rect	192	182	193	183
rect	192	183	193	184
rect	192	185	193	186
rect	192	186	193	187
rect	192	188	193	189
rect	192	189	193	190
rect	192	191	193	192
rect	192	192	193	193
rect	192	194	193	195
rect	192	195	193	196
rect	192	197	193	198
rect	192	198	193	199
rect	192	200	193	201
rect	192	201	193	202
rect	192	203	193	204
rect	192	204	193	205
rect	192	206	193	207
rect	192	207	193	208
rect	192	209	193	210
rect	192	210	193	211
rect	192	212	193	213
rect	192	213	193	214
rect	192	215	193	216
rect	192	216	193	217
rect	192	218	193	219
rect	192	219	193	220
rect	192	221	193	222
rect	192	222	193	223
rect	192	224	193	225
rect	192	225	193	226
rect	192	227	193	228
rect	192	228	193	229
rect	192	230	193	231
rect	192	231	193	232
rect	192	233	193	234
rect	192	234	193	235
rect	192	236	193	237
rect	192	237	193	238
rect	192	239	193	240
rect	192	240	193	241
rect	192	242	193	243
rect	192	243	193	244
rect	192	245	193	246
rect	192	246	193	247
rect	192	248	193	249
rect	192	249	193	250
rect	192	251	193	252
rect	192	252	193	253
rect	192	254	193	255
rect	192	255	193	256
rect	192	257	193	258
rect	192	258	193	259
rect	192	260	193	261
rect	192	261	193	262
rect	192	262	193	263
rect	192	263	193	264
rect	192	264	193	265
rect	192	266	193	267
rect	192	267	193	268
rect	192	269	193	270
rect	192	270	193	271
rect	192	272	193	273
rect	192	273	193	274
rect	192	275	193	276
rect	192	276	193	277
rect	192	278	193	279
rect	192	279	193	280
rect	192	281	193	282
rect	192	282	193	283
rect	192	284	193	285
rect	192	285	193	286
rect	192	287	193	288
rect	192	288	193	289
rect	192	290	193	291
rect	192	291	193	292
rect	192	293	193	294
rect	192	294	193	295
rect	192	296	193	297
rect	192	297	193	298
rect	192	299	193	300
rect	192	300	193	301
rect	192	302	193	303
rect	192	303	193	304
rect	192	304	193	305
rect	192	305	193	306
rect	192	306	193	307
rect	192	308	193	309
rect	192	309	193	310
rect	192	311	193	312
rect	192	312	193	313
rect	192	314	193	315
rect	192	315	193	316
rect	192	317	193	318
rect	192	318	193	319
rect	192	319	193	320
rect	192	320	193	321
rect	192	321	193	322
rect	192	322	193	323
rect	192	323	193	324
rect	192	324	193	325
rect	192	325	193	326
rect	192	326	193	327
rect	192	327	193	328
rect	192	328	193	329
rect	192	329	193	330
rect	192	330	193	331
rect	192	332	193	333
rect	192	333	193	334
rect	192	335	193	336
rect	192	336	193	337
rect	192	337	193	338
rect	192	338	193	339
rect	192	339	193	340
rect	192	340	193	341
rect	192	341	193	342
rect	192	342	193	343
rect	192	343	193	344
rect	192	344	193	345
rect	192	345	193	346
rect	192	347	193	348
rect	192	348	193	349
rect	192	349	193	350
rect	192	350	193	351
rect	192	351	193	352
rect	192	352	193	353
rect	192	353	193	354
rect	192	354	193	355
rect	192	355	193	356
rect	192	356	193	357
rect	192	357	193	358
rect	192	358	193	359
rect	192	359	193	360
rect	192	360	193	361
rect	192	361	193	362
rect	192	362	193	363
rect	192	363	193	364
rect	192	364	193	365
rect	192	365	193	366
rect	192	366	193	367
rect	192	367	193	368
rect	192	368	193	369
rect	194	0	195	1
rect	194	1	195	2
rect	194	2	195	3
rect	194	3	195	4
rect	194	5	195	6
rect	194	6	195	7
rect	194	8	195	9
rect	194	9	195	10
rect	194	11	195	12
rect	194	12	195	13
rect	194	14	195	15
rect	194	15	195	16
rect	194	17	195	18
rect	194	18	195	19
rect	194	20	195	21
rect	194	21	195	22
rect	194	23	195	24
rect	194	24	195	25
rect	194	26	195	27
rect	194	27	195	28
rect	194	29	195	30
rect	194	30	195	31
rect	194	32	195	33
rect	194	33	195	34
rect	194	35	195	36
rect	194	36	195	37
rect	194	38	195	39
rect	194	39	195	40
rect	194	41	195	42
rect	194	42	195	43
rect	194	44	195	45
rect	194	45	195	46
rect	194	47	195	48
rect	194	48	195	49
rect	194	50	195	51
rect	194	51	195	52
rect	194	53	195	54
rect	194	54	195	55
rect	194	56	195	57
rect	194	57	195	58
rect	194	59	195	60
rect	194	60	195	61
rect	194	62	195	63
rect	194	63	195	64
rect	194	65	195	66
rect	194	66	195	67
rect	194	68	195	69
rect	194	69	195	70
rect	194	71	195	72
rect	194	72	195	73
rect	194	74	195	75
rect	194	75	195	76
rect	194	77	195	78
rect	194	78	195	79
rect	194	80	195	81
rect	194	81	195	82
rect	194	83	195	84
rect	194	84	195	85
rect	194	86	195	87
rect	194	87	195	88
rect	194	89	195	90
rect	194	90	195	91
rect	194	92	195	93
rect	194	93	195	94
rect	194	95	195	96
rect	194	96	195	97
rect	194	98	195	99
rect	194	99	195	100
rect	194	101	195	102
rect	194	102	195	103
rect	194	104	195	105
rect	194	105	195	106
rect	194	107	195	108
rect	194	108	195	109
rect	194	110	195	111
rect	194	111	195	112
rect	194	113	195	114
rect	194	114	195	115
rect	194	116	195	117
rect	194	117	195	118
rect	194	119	195	120
rect	194	120	195	121
rect	194	122	195	123
rect	194	123	195	124
rect	194	125	195	126
rect	194	126	195	127
rect	194	128	195	129
rect	194	129	195	130
rect	194	131	195	132
rect	194	132	195	133
rect	194	134	195	135
rect	194	135	195	136
rect	194	137	195	138
rect	194	138	195	139
rect	194	140	195	141
rect	194	141	195	142
rect	194	143	195	144
rect	194	144	195	145
rect	194	146	195	147
rect	194	147	195	148
rect	194	149	195	150
rect	194	150	195	151
rect	194	152	195	153
rect	194	153	195	154
rect	194	155	195	156
rect	194	156	195	157
rect	194	158	195	159
rect	194	159	195	160
rect	194	161	195	162
rect	194	162	195	163
rect	194	164	195	165
rect	194	165	195	166
rect	194	167	195	168
rect	194	168	195	169
rect	194	170	195	171
rect	194	171	195	172
rect	194	173	195	174
rect	194	174	195	175
rect	194	176	195	177
rect	194	177	195	178
rect	194	179	195	180
rect	194	180	195	181
rect	194	182	195	183
rect	194	183	195	184
rect	194	185	195	186
rect	194	186	195	187
rect	194	188	195	189
rect	194	189	195	190
rect	194	191	195	192
rect	194	192	195	193
rect	194	194	195	195
rect	194	195	195	196
rect	194	197	195	198
rect	194	198	195	199
rect	194	200	195	201
rect	194	201	195	202
rect	194	203	195	204
rect	194	204	195	205
rect	194	206	195	207
rect	194	207	195	208
rect	194	209	195	210
rect	194	210	195	211
rect	194	212	195	213
rect	194	213	195	214
rect	194	215	195	216
rect	194	216	195	217
rect	194	218	195	219
rect	194	219	195	220
rect	194	221	195	222
rect	194	222	195	223
rect	194	224	195	225
rect	194	225	195	226
rect	194	227	195	228
rect	194	228	195	229
rect	194	230	195	231
rect	194	231	195	232
rect	194	233	195	234
rect	194	234	195	235
rect	194	236	195	237
rect	194	237	195	238
rect	194	239	195	240
rect	194	240	195	241
rect	194	242	195	243
rect	194	243	195	244
rect	194	245	195	246
rect	194	246	195	247
rect	194	248	195	249
rect	194	249	195	250
rect	194	251	195	252
rect	194	252	195	253
rect	194	254	195	255
rect	194	255	195	256
rect	194	257	195	258
rect	194	258	195	259
rect	194	260	195	261
rect	194	261	195	262
rect	194	262	195	263
rect	194	263	195	264
rect	194	264	195	265
rect	194	266	195	267
rect	194	267	195	268
rect	194	269	195	270
rect	194	270	195	271
rect	194	272	195	273
rect	194	273	195	274
rect	194	275	195	276
rect	194	276	195	277
rect	194	278	195	279
rect	194	279	195	280
rect	194	281	195	282
rect	194	282	195	283
rect	194	284	195	285
rect	194	285	195	286
rect	194	287	195	288
rect	194	288	195	289
rect	194	290	195	291
rect	194	291	195	292
rect	194	293	195	294
rect	194	294	195	295
rect	194	296	195	297
rect	194	297	195	298
rect	194	299	195	300
rect	194	300	195	301
rect	194	302	195	303
rect	194	303	195	304
rect	194	304	195	305
rect	194	305	195	306
rect	194	306	195	307
rect	194	308	195	309
rect	194	309	195	310
rect	194	311	195	312
rect	194	312	195	313
rect	194	314	195	315
rect	194	315	195	316
rect	194	317	195	318
rect	194	318	195	319
rect	194	319	195	320
rect	194	320	195	321
rect	194	321	195	322
rect	194	322	195	323
rect	194	323	195	324
rect	194	324	195	325
rect	194	325	195	326
rect	194	326	195	327
rect	194	327	195	328
rect	194	328	195	329
rect	194	329	195	330
rect	194	330	195	331
rect	194	332	195	333
rect	194	333	195	334
rect	194	335	195	336
rect	194	336	195	337
rect	194	337	195	338
rect	194	338	195	339
rect	194	339	195	340
rect	194	340	195	341
rect	194	341	195	342
rect	194	342	195	343
rect	194	343	195	344
rect	194	344	195	345
rect	194	345	195	346
rect	194	347	195	348
rect	195	0	196	1
rect	195	1	196	2
rect	195	2	196	3
rect	195	3	196	4
rect	195	5	196	6
rect	195	6	196	7
rect	195	8	196	9
rect	195	9	196	10
rect	195	11	196	12
rect	195	12	196	13
rect	195	14	196	15
rect	195	15	196	16
rect	195	17	196	18
rect	195	18	196	19
rect	195	20	196	21
rect	195	21	196	22
rect	195	23	196	24
rect	195	24	196	25
rect	195	26	196	27
rect	195	27	196	28
rect	195	29	196	30
rect	195	30	196	31
rect	195	32	196	33
rect	195	33	196	34
rect	195	35	196	36
rect	195	36	196	37
rect	195	38	196	39
rect	195	39	196	40
rect	195	41	196	42
rect	195	42	196	43
rect	195	44	196	45
rect	195	45	196	46
rect	195	47	196	48
rect	195	48	196	49
rect	195	50	196	51
rect	195	51	196	52
rect	195	53	196	54
rect	195	54	196	55
rect	195	56	196	57
rect	195	57	196	58
rect	195	59	196	60
rect	195	60	196	61
rect	195	62	196	63
rect	195	63	196	64
rect	195	65	196	66
rect	195	66	196	67
rect	195	68	196	69
rect	195	69	196	70
rect	195	71	196	72
rect	195	72	196	73
rect	195	74	196	75
rect	195	75	196	76
rect	195	77	196	78
rect	195	78	196	79
rect	195	80	196	81
rect	195	81	196	82
rect	195	83	196	84
rect	195	84	196	85
rect	195	86	196	87
rect	195	87	196	88
rect	195	89	196	90
rect	195	90	196	91
rect	195	92	196	93
rect	195	93	196	94
rect	195	95	196	96
rect	195	96	196	97
rect	195	98	196	99
rect	195	99	196	100
rect	195	101	196	102
rect	195	102	196	103
rect	195	104	196	105
rect	195	105	196	106
rect	195	107	196	108
rect	195	108	196	109
rect	195	110	196	111
rect	195	111	196	112
rect	195	113	196	114
rect	195	114	196	115
rect	195	116	196	117
rect	195	117	196	118
rect	195	119	196	120
rect	195	120	196	121
rect	195	122	196	123
rect	195	123	196	124
rect	195	125	196	126
rect	195	126	196	127
rect	195	128	196	129
rect	195	129	196	130
rect	195	131	196	132
rect	195	132	196	133
rect	195	134	196	135
rect	195	135	196	136
rect	195	137	196	138
rect	195	138	196	139
rect	195	140	196	141
rect	195	141	196	142
rect	195	143	196	144
rect	195	144	196	145
rect	195	146	196	147
rect	195	147	196	148
rect	195	149	196	150
rect	195	150	196	151
rect	195	152	196	153
rect	195	153	196	154
rect	195	155	196	156
rect	195	156	196	157
rect	195	158	196	159
rect	195	159	196	160
rect	195	161	196	162
rect	195	162	196	163
rect	195	164	196	165
rect	195	165	196	166
rect	195	167	196	168
rect	195	168	196	169
rect	195	170	196	171
rect	195	171	196	172
rect	195	173	196	174
rect	195	174	196	175
rect	195	176	196	177
rect	195	177	196	178
rect	195	179	196	180
rect	195	180	196	181
rect	195	182	196	183
rect	195	183	196	184
rect	195	185	196	186
rect	195	186	196	187
rect	195	188	196	189
rect	195	189	196	190
rect	195	191	196	192
rect	195	192	196	193
rect	195	194	196	195
rect	195	195	196	196
rect	195	197	196	198
rect	195	198	196	199
rect	195	200	196	201
rect	195	201	196	202
rect	195	203	196	204
rect	195	204	196	205
rect	195	206	196	207
rect	195	207	196	208
rect	195	209	196	210
rect	195	210	196	211
rect	195	212	196	213
rect	195	213	196	214
rect	195	215	196	216
rect	195	216	196	217
rect	195	218	196	219
rect	195	219	196	220
rect	195	221	196	222
rect	195	222	196	223
rect	195	224	196	225
rect	195	225	196	226
rect	195	227	196	228
rect	195	228	196	229
rect	195	230	196	231
rect	195	231	196	232
rect	195	233	196	234
rect	195	234	196	235
rect	195	236	196	237
rect	195	237	196	238
rect	195	239	196	240
rect	195	240	196	241
rect	195	242	196	243
rect	195	243	196	244
rect	195	245	196	246
rect	195	246	196	247
rect	195	248	196	249
rect	195	249	196	250
rect	195	251	196	252
rect	195	252	196	253
rect	195	254	196	255
rect	195	255	196	256
rect	195	257	196	258
rect	195	258	196	259
rect	195	260	196	261
rect	195	261	196	262
rect	195	262	196	263
rect	195	263	196	264
rect	195	264	196	265
rect	195	266	196	267
rect	195	267	196	268
rect	195	269	196	270
rect	195	270	196	271
rect	195	272	196	273
rect	195	273	196	274
rect	195	275	196	276
rect	195	276	196	277
rect	195	278	196	279
rect	195	279	196	280
rect	195	281	196	282
rect	195	282	196	283
rect	195	284	196	285
rect	195	285	196	286
rect	195	287	196	288
rect	195	288	196	289
rect	195	290	196	291
rect	195	291	196	292
rect	195	293	196	294
rect	195	294	196	295
rect	195	296	196	297
rect	195	297	196	298
rect	195	299	196	300
rect	195	300	196	301
rect	195	302	196	303
rect	195	303	196	304
rect	195	304	196	305
rect	195	305	196	306
rect	195	306	196	307
rect	195	308	196	309
rect	195	309	196	310
rect	195	311	196	312
rect	195	312	196	313
rect	195	314	196	315
rect	195	315	196	316
rect	195	317	196	318
rect	195	318	196	319
rect	195	319	196	320
rect	195	320	196	321
rect	195	321	196	322
rect	195	322	196	323
rect	195	323	196	324
rect	195	324	196	325
rect	195	325	196	326
rect	195	326	196	327
rect	195	327	196	328
rect	195	328	196	329
rect	195	329	196	330
rect	195	330	196	331
rect	195	332	196	333
rect	195	333	196	334
rect	195	335	196	336
rect	195	336	196	337
rect	195	337	196	338
rect	195	338	196	339
rect	195	339	196	340
rect	195	340	196	341
rect	195	341	196	342
rect	195	342	196	343
rect	195	343	196	344
rect	195	344	196	345
rect	195	345	196	346
rect	195	347	196	348
rect	196	0	197	1
rect	196	1	197	2
rect	196	2	197	3
rect	196	3	197	4
rect	196	5	197	6
rect	196	6	197	7
rect	196	8	197	9
rect	196	9	197	10
rect	196	11	197	12
rect	196	12	197	13
rect	196	14	197	15
rect	196	15	197	16
rect	196	17	197	18
rect	196	18	197	19
rect	196	20	197	21
rect	196	21	197	22
rect	196	23	197	24
rect	196	24	197	25
rect	196	26	197	27
rect	196	27	197	28
rect	196	29	197	30
rect	196	30	197	31
rect	196	32	197	33
rect	196	33	197	34
rect	196	35	197	36
rect	196	36	197	37
rect	196	38	197	39
rect	196	39	197	40
rect	196	41	197	42
rect	196	42	197	43
rect	196	44	197	45
rect	196	45	197	46
rect	196	47	197	48
rect	196	48	197	49
rect	196	50	197	51
rect	196	51	197	52
rect	196	53	197	54
rect	196	54	197	55
rect	196	56	197	57
rect	196	57	197	58
rect	196	59	197	60
rect	196	60	197	61
rect	196	62	197	63
rect	196	63	197	64
rect	196	65	197	66
rect	196	66	197	67
rect	196	68	197	69
rect	196	69	197	70
rect	196	71	197	72
rect	196	72	197	73
rect	196	74	197	75
rect	196	75	197	76
rect	196	77	197	78
rect	196	78	197	79
rect	196	80	197	81
rect	196	81	197	82
rect	196	83	197	84
rect	196	84	197	85
rect	196	86	197	87
rect	196	87	197	88
rect	196	89	197	90
rect	196	90	197	91
rect	196	92	197	93
rect	196	93	197	94
rect	196	95	197	96
rect	196	96	197	97
rect	196	98	197	99
rect	196	99	197	100
rect	196	101	197	102
rect	196	102	197	103
rect	196	104	197	105
rect	196	105	197	106
rect	196	107	197	108
rect	196	108	197	109
rect	196	110	197	111
rect	196	111	197	112
rect	196	113	197	114
rect	196	114	197	115
rect	196	116	197	117
rect	196	117	197	118
rect	196	119	197	120
rect	196	120	197	121
rect	196	122	197	123
rect	196	123	197	124
rect	196	125	197	126
rect	196	126	197	127
rect	196	128	197	129
rect	196	129	197	130
rect	196	131	197	132
rect	196	132	197	133
rect	196	134	197	135
rect	196	135	197	136
rect	196	137	197	138
rect	196	138	197	139
rect	196	140	197	141
rect	196	141	197	142
rect	196	143	197	144
rect	196	144	197	145
rect	196	146	197	147
rect	196	147	197	148
rect	196	149	197	150
rect	196	150	197	151
rect	196	152	197	153
rect	196	153	197	154
rect	196	155	197	156
rect	196	156	197	157
rect	196	158	197	159
rect	196	159	197	160
rect	196	161	197	162
rect	196	162	197	163
rect	196	164	197	165
rect	196	165	197	166
rect	196	167	197	168
rect	196	168	197	169
rect	196	170	197	171
rect	196	171	197	172
rect	196	173	197	174
rect	196	174	197	175
rect	196	176	197	177
rect	196	177	197	178
rect	196	179	197	180
rect	196	180	197	181
rect	196	182	197	183
rect	196	183	197	184
rect	196	185	197	186
rect	196	186	197	187
rect	196	188	197	189
rect	196	189	197	190
rect	196	191	197	192
rect	196	192	197	193
rect	196	194	197	195
rect	196	195	197	196
rect	196	197	197	198
rect	196	198	197	199
rect	196	200	197	201
rect	196	201	197	202
rect	196	203	197	204
rect	196	204	197	205
rect	196	206	197	207
rect	196	207	197	208
rect	196	209	197	210
rect	196	210	197	211
rect	196	212	197	213
rect	196	213	197	214
rect	196	215	197	216
rect	196	216	197	217
rect	196	218	197	219
rect	196	219	197	220
rect	196	221	197	222
rect	196	222	197	223
rect	196	224	197	225
rect	196	225	197	226
rect	196	227	197	228
rect	196	228	197	229
rect	196	230	197	231
rect	196	231	197	232
rect	196	233	197	234
rect	196	234	197	235
rect	196	236	197	237
rect	196	237	197	238
rect	196	239	197	240
rect	196	240	197	241
rect	196	242	197	243
rect	196	243	197	244
rect	196	245	197	246
rect	196	246	197	247
rect	196	248	197	249
rect	196	249	197	250
rect	196	251	197	252
rect	196	252	197	253
rect	196	254	197	255
rect	196	255	197	256
rect	196	257	197	258
rect	196	258	197	259
rect	196	260	197	261
rect	196	261	197	262
rect	196	262	197	263
rect	196	263	197	264
rect	196	264	197	265
rect	196	266	197	267
rect	196	267	197	268
rect	196	269	197	270
rect	196	270	197	271
rect	196	272	197	273
rect	196	273	197	274
rect	196	275	197	276
rect	196	276	197	277
rect	196	278	197	279
rect	196	279	197	280
rect	196	281	197	282
rect	196	282	197	283
rect	196	284	197	285
rect	196	285	197	286
rect	196	287	197	288
rect	196	288	197	289
rect	196	290	197	291
rect	196	291	197	292
rect	196	293	197	294
rect	196	294	197	295
rect	196	296	197	297
rect	196	297	197	298
rect	196	299	197	300
rect	196	300	197	301
rect	196	302	197	303
rect	196	303	197	304
rect	196	304	197	305
rect	196	305	197	306
rect	196	306	197	307
rect	196	308	197	309
rect	196	309	197	310
rect	196	311	197	312
rect	196	312	197	313
rect	196	314	197	315
rect	196	315	197	316
rect	196	317	197	318
rect	196	318	197	319
rect	196	319	197	320
rect	196	320	197	321
rect	196	321	197	322
rect	196	322	197	323
rect	196	323	197	324
rect	196	324	197	325
rect	196	325	197	326
rect	196	326	197	327
rect	196	327	197	328
rect	196	328	197	329
rect	196	329	197	330
rect	196	330	197	331
rect	196	332	197	333
rect	196	333	197	334
rect	196	335	197	336
rect	196	336	197	337
rect	196	337	197	338
rect	196	338	197	339
rect	196	339	197	340
rect	196	340	197	341
rect	196	341	197	342
rect	196	342	197	343
rect	196	343	197	344
rect	196	344	197	345
rect	196	345	197	346
rect	196	347	197	348
rect	197	0	198	1
rect	197	1	198	2
rect	197	2	198	3
rect	197	3	198	4
rect	197	5	198	6
rect	197	6	198	7
rect	197	8	198	9
rect	197	9	198	10
rect	197	11	198	12
rect	197	12	198	13
rect	197	14	198	15
rect	197	15	198	16
rect	197	17	198	18
rect	197	18	198	19
rect	197	20	198	21
rect	197	21	198	22
rect	197	23	198	24
rect	197	24	198	25
rect	197	26	198	27
rect	197	27	198	28
rect	197	29	198	30
rect	197	30	198	31
rect	197	32	198	33
rect	197	33	198	34
rect	197	35	198	36
rect	197	36	198	37
rect	197	38	198	39
rect	197	39	198	40
rect	197	41	198	42
rect	197	42	198	43
rect	197	44	198	45
rect	197	45	198	46
rect	197	47	198	48
rect	197	48	198	49
rect	197	50	198	51
rect	197	51	198	52
rect	197	53	198	54
rect	197	54	198	55
rect	197	56	198	57
rect	197	57	198	58
rect	197	59	198	60
rect	197	60	198	61
rect	197	62	198	63
rect	197	63	198	64
rect	197	65	198	66
rect	197	66	198	67
rect	197	68	198	69
rect	197	69	198	70
rect	197	71	198	72
rect	197	72	198	73
rect	197	74	198	75
rect	197	75	198	76
rect	197	77	198	78
rect	197	78	198	79
rect	197	80	198	81
rect	197	81	198	82
rect	197	83	198	84
rect	197	84	198	85
rect	197	86	198	87
rect	197	87	198	88
rect	197	89	198	90
rect	197	90	198	91
rect	197	92	198	93
rect	197	93	198	94
rect	197	95	198	96
rect	197	96	198	97
rect	197	98	198	99
rect	197	99	198	100
rect	197	101	198	102
rect	197	102	198	103
rect	197	104	198	105
rect	197	105	198	106
rect	197	107	198	108
rect	197	108	198	109
rect	197	110	198	111
rect	197	111	198	112
rect	197	113	198	114
rect	197	114	198	115
rect	197	116	198	117
rect	197	117	198	118
rect	197	119	198	120
rect	197	120	198	121
rect	197	122	198	123
rect	197	123	198	124
rect	197	125	198	126
rect	197	126	198	127
rect	197	128	198	129
rect	197	129	198	130
rect	197	131	198	132
rect	197	132	198	133
rect	197	134	198	135
rect	197	135	198	136
rect	197	137	198	138
rect	197	138	198	139
rect	197	140	198	141
rect	197	141	198	142
rect	197	143	198	144
rect	197	144	198	145
rect	197	146	198	147
rect	197	147	198	148
rect	197	149	198	150
rect	197	150	198	151
rect	197	152	198	153
rect	197	153	198	154
rect	197	155	198	156
rect	197	156	198	157
rect	197	158	198	159
rect	197	159	198	160
rect	197	161	198	162
rect	197	162	198	163
rect	197	164	198	165
rect	197	165	198	166
rect	197	167	198	168
rect	197	168	198	169
rect	197	170	198	171
rect	197	171	198	172
rect	197	173	198	174
rect	197	174	198	175
rect	197	176	198	177
rect	197	177	198	178
rect	197	179	198	180
rect	197	180	198	181
rect	197	182	198	183
rect	197	183	198	184
rect	197	185	198	186
rect	197	186	198	187
rect	197	188	198	189
rect	197	189	198	190
rect	197	191	198	192
rect	197	192	198	193
rect	197	194	198	195
rect	197	195	198	196
rect	197	197	198	198
rect	197	198	198	199
rect	197	200	198	201
rect	197	201	198	202
rect	197	203	198	204
rect	197	204	198	205
rect	197	206	198	207
rect	197	207	198	208
rect	197	209	198	210
rect	197	210	198	211
rect	197	212	198	213
rect	197	213	198	214
rect	197	215	198	216
rect	197	216	198	217
rect	197	218	198	219
rect	197	219	198	220
rect	197	221	198	222
rect	197	222	198	223
rect	197	224	198	225
rect	197	225	198	226
rect	197	227	198	228
rect	197	228	198	229
rect	197	230	198	231
rect	197	231	198	232
rect	197	233	198	234
rect	197	234	198	235
rect	197	236	198	237
rect	197	237	198	238
rect	197	239	198	240
rect	197	240	198	241
rect	197	242	198	243
rect	197	243	198	244
rect	197	245	198	246
rect	197	246	198	247
rect	197	248	198	249
rect	197	249	198	250
rect	197	251	198	252
rect	197	252	198	253
rect	197	254	198	255
rect	197	255	198	256
rect	197	257	198	258
rect	197	258	198	259
rect	197	260	198	261
rect	197	261	198	262
rect	197	262	198	263
rect	197	263	198	264
rect	197	264	198	265
rect	197	266	198	267
rect	197	267	198	268
rect	197	269	198	270
rect	197	270	198	271
rect	197	272	198	273
rect	197	273	198	274
rect	197	275	198	276
rect	197	276	198	277
rect	197	278	198	279
rect	197	279	198	280
rect	197	281	198	282
rect	197	282	198	283
rect	197	284	198	285
rect	197	285	198	286
rect	197	287	198	288
rect	197	288	198	289
rect	197	290	198	291
rect	197	291	198	292
rect	197	293	198	294
rect	197	294	198	295
rect	197	296	198	297
rect	197	297	198	298
rect	197	299	198	300
rect	197	300	198	301
rect	197	302	198	303
rect	197	303	198	304
rect	197	304	198	305
rect	197	305	198	306
rect	197	306	198	307
rect	197	308	198	309
rect	197	309	198	310
rect	197	311	198	312
rect	197	312	198	313
rect	197	314	198	315
rect	197	315	198	316
rect	197	317	198	318
rect	197	318	198	319
rect	197	319	198	320
rect	197	320	198	321
rect	197	321	198	322
rect	197	322	198	323
rect	197	323	198	324
rect	197	324	198	325
rect	197	325	198	326
rect	197	326	198	327
rect	197	327	198	328
rect	197	328	198	329
rect	197	329	198	330
rect	197	330	198	331
rect	197	332	198	333
rect	197	333	198	334
rect	197	335	198	336
rect	197	336	198	337
rect	197	337	198	338
rect	197	338	198	339
rect	197	339	198	340
rect	197	340	198	341
rect	197	341	198	342
rect	197	342	198	343
rect	197	343	198	344
rect	197	344	198	345
rect	197	345	198	346
rect	197	347	198	348
rect	198	0	199	1
rect	198	1	199	2
rect	198	2	199	3
rect	198	3	199	4
rect	198	5	199	6
rect	198	6	199	7
rect	198	8	199	9
rect	198	9	199	10
rect	198	11	199	12
rect	198	12	199	13
rect	198	14	199	15
rect	198	15	199	16
rect	198	17	199	18
rect	198	18	199	19
rect	198	20	199	21
rect	198	21	199	22
rect	198	23	199	24
rect	198	24	199	25
rect	198	26	199	27
rect	198	27	199	28
rect	198	29	199	30
rect	198	30	199	31
rect	198	32	199	33
rect	198	33	199	34
rect	198	35	199	36
rect	198	36	199	37
rect	198	38	199	39
rect	198	39	199	40
rect	198	41	199	42
rect	198	42	199	43
rect	198	44	199	45
rect	198	45	199	46
rect	198	47	199	48
rect	198	48	199	49
rect	198	50	199	51
rect	198	51	199	52
rect	198	53	199	54
rect	198	54	199	55
rect	198	56	199	57
rect	198	57	199	58
rect	198	59	199	60
rect	198	60	199	61
rect	198	62	199	63
rect	198	63	199	64
rect	198	65	199	66
rect	198	66	199	67
rect	198	68	199	69
rect	198	69	199	70
rect	198	71	199	72
rect	198	72	199	73
rect	198	74	199	75
rect	198	75	199	76
rect	198	77	199	78
rect	198	78	199	79
rect	198	80	199	81
rect	198	81	199	82
rect	198	83	199	84
rect	198	84	199	85
rect	198	86	199	87
rect	198	87	199	88
rect	198	89	199	90
rect	198	90	199	91
rect	198	92	199	93
rect	198	93	199	94
rect	198	95	199	96
rect	198	96	199	97
rect	198	98	199	99
rect	198	99	199	100
rect	198	101	199	102
rect	198	102	199	103
rect	198	104	199	105
rect	198	105	199	106
rect	198	107	199	108
rect	198	108	199	109
rect	198	110	199	111
rect	198	111	199	112
rect	198	113	199	114
rect	198	114	199	115
rect	198	116	199	117
rect	198	117	199	118
rect	198	119	199	120
rect	198	120	199	121
rect	198	122	199	123
rect	198	123	199	124
rect	198	125	199	126
rect	198	126	199	127
rect	198	128	199	129
rect	198	129	199	130
rect	198	131	199	132
rect	198	132	199	133
rect	198	134	199	135
rect	198	135	199	136
rect	198	137	199	138
rect	198	138	199	139
rect	198	140	199	141
rect	198	141	199	142
rect	198	143	199	144
rect	198	144	199	145
rect	198	146	199	147
rect	198	147	199	148
rect	198	149	199	150
rect	198	150	199	151
rect	198	152	199	153
rect	198	153	199	154
rect	198	155	199	156
rect	198	156	199	157
rect	198	158	199	159
rect	198	159	199	160
rect	198	161	199	162
rect	198	162	199	163
rect	198	164	199	165
rect	198	165	199	166
rect	198	167	199	168
rect	198	168	199	169
rect	198	170	199	171
rect	198	171	199	172
rect	198	173	199	174
rect	198	174	199	175
rect	198	176	199	177
rect	198	177	199	178
rect	198	179	199	180
rect	198	180	199	181
rect	198	182	199	183
rect	198	183	199	184
rect	198	185	199	186
rect	198	186	199	187
rect	198	188	199	189
rect	198	189	199	190
rect	198	191	199	192
rect	198	192	199	193
rect	198	194	199	195
rect	198	195	199	196
rect	198	197	199	198
rect	198	198	199	199
rect	198	200	199	201
rect	198	201	199	202
rect	198	203	199	204
rect	198	204	199	205
rect	198	206	199	207
rect	198	207	199	208
rect	198	209	199	210
rect	198	210	199	211
rect	198	212	199	213
rect	198	213	199	214
rect	198	215	199	216
rect	198	216	199	217
rect	198	218	199	219
rect	198	219	199	220
rect	198	221	199	222
rect	198	222	199	223
rect	198	224	199	225
rect	198	225	199	226
rect	198	227	199	228
rect	198	228	199	229
rect	198	230	199	231
rect	198	231	199	232
rect	198	233	199	234
rect	198	234	199	235
rect	198	236	199	237
rect	198	237	199	238
rect	198	239	199	240
rect	198	240	199	241
rect	198	242	199	243
rect	198	243	199	244
rect	198	245	199	246
rect	198	246	199	247
rect	198	248	199	249
rect	198	249	199	250
rect	198	251	199	252
rect	198	252	199	253
rect	198	254	199	255
rect	198	255	199	256
rect	198	257	199	258
rect	198	258	199	259
rect	198	260	199	261
rect	198	261	199	262
rect	198	262	199	263
rect	198	263	199	264
rect	198	264	199	265
rect	198	266	199	267
rect	198	267	199	268
rect	198	269	199	270
rect	198	270	199	271
rect	198	272	199	273
rect	198	273	199	274
rect	198	275	199	276
rect	198	276	199	277
rect	198	278	199	279
rect	198	279	199	280
rect	198	281	199	282
rect	198	282	199	283
rect	198	284	199	285
rect	198	285	199	286
rect	198	287	199	288
rect	198	288	199	289
rect	198	290	199	291
rect	198	291	199	292
rect	198	293	199	294
rect	198	294	199	295
rect	198	296	199	297
rect	198	297	199	298
rect	198	299	199	300
rect	198	300	199	301
rect	198	302	199	303
rect	198	303	199	304
rect	198	304	199	305
rect	198	305	199	306
rect	198	306	199	307
rect	198	308	199	309
rect	198	309	199	310
rect	198	311	199	312
rect	198	312	199	313
rect	198	314	199	315
rect	198	315	199	316
rect	198	317	199	318
rect	198	318	199	319
rect	198	319	199	320
rect	198	320	199	321
rect	198	321	199	322
rect	198	322	199	323
rect	198	323	199	324
rect	198	324	199	325
rect	198	325	199	326
rect	198	326	199	327
rect	198	327	199	328
rect	198	328	199	329
rect	198	329	199	330
rect	198	330	199	331
rect	198	332	199	333
rect	198	333	199	334
rect	198	335	199	336
rect	198	336	199	337
rect	198	337	199	338
rect	198	338	199	339
rect	198	339	199	340
rect	198	340	199	341
rect	198	341	199	342
rect	198	342	199	343
rect	198	343	199	344
rect	198	344	199	345
rect	198	345	199	346
rect	198	347	199	348
rect	209	0	210	1
rect	209	1	210	2
rect	209	2	210	3
rect	209	3	210	4
rect	209	4	210	5
rect	209	5	210	6
rect	209	6	210	7
rect	209	8	210	9
rect	209	9	210	10
rect	209	11	210	12
rect	209	12	210	13
rect	209	14	210	15
rect	209	15	210	16
rect	209	17	210	18
rect	209	18	210	19
rect	209	20	210	21
rect	209	21	210	22
rect	209	23	210	24
rect	209	24	210	25
rect	209	26	210	27
rect	209	27	210	28
rect	209	29	210	30
rect	209	30	210	31
rect	209	32	210	33
rect	209	33	210	34
rect	209	35	210	36
rect	209	36	210	37
rect	209	38	210	39
rect	209	39	210	40
rect	209	41	210	42
rect	209	42	210	43
rect	209	44	210	45
rect	209	45	210	46
rect	209	47	210	48
rect	209	48	210	49
rect	209	50	210	51
rect	209	51	210	52
rect	209	53	210	54
rect	209	54	210	55
rect	209	56	210	57
rect	209	57	210	58
rect	209	59	210	60
rect	209	60	210	61
rect	209	62	210	63
rect	209	63	210	64
rect	209	65	210	66
rect	209	66	210	67
rect	209	68	210	69
rect	209	69	210	70
rect	209	71	210	72
rect	209	72	210	73
rect	209	74	210	75
rect	209	75	210	76
rect	209	77	210	78
rect	209	78	210	79
rect	209	80	210	81
rect	209	81	210	82
rect	209	83	210	84
rect	209	84	210	85
rect	209	86	210	87
rect	209	87	210	88
rect	209	89	210	90
rect	209	90	210	91
rect	209	92	210	93
rect	209	93	210	94
rect	209	95	210	96
rect	209	96	210	97
rect	209	98	210	99
rect	209	99	210	100
rect	209	101	210	102
rect	209	102	210	103
rect	209	104	210	105
rect	209	105	210	106
rect	209	107	210	108
rect	209	108	210	109
rect	209	110	210	111
rect	209	111	210	112
rect	209	113	210	114
rect	209	114	210	115
rect	209	116	210	117
rect	209	117	210	118
rect	209	119	210	120
rect	209	120	210	121
rect	209	122	210	123
rect	209	123	210	124
rect	209	125	210	126
rect	209	126	210	127
rect	209	128	210	129
rect	209	129	210	130
rect	209	131	210	132
rect	209	132	210	133
rect	209	134	210	135
rect	209	135	210	136
rect	209	137	210	138
rect	209	138	210	139
rect	209	140	210	141
rect	209	141	210	142
rect	209	143	210	144
rect	209	144	210	145
rect	209	146	210	147
rect	209	147	210	148
rect	209	149	210	150
rect	209	150	210	151
rect	209	152	210	153
rect	209	153	210	154
rect	209	155	210	156
rect	209	156	210	157
rect	209	158	210	159
rect	209	159	210	160
rect	209	161	210	162
rect	209	162	210	163
rect	209	164	210	165
rect	209	165	210	166
rect	209	167	210	168
rect	209	168	210	169
rect	209	170	210	171
rect	209	171	210	172
rect	209	173	210	174
rect	209	174	210	175
rect	209	176	210	177
rect	209	177	210	178
rect	209	179	210	180
rect	209	180	210	181
rect	209	182	210	183
rect	209	183	210	184
rect	209	185	210	186
rect	209	186	210	187
rect	209	188	210	189
rect	209	189	210	190
rect	209	191	210	192
rect	209	192	210	193
rect	209	194	210	195
rect	209	195	210	196
rect	209	197	210	198
rect	209	198	210	199
rect	209	200	210	201
rect	209	201	210	202
rect	209	203	210	204
rect	209	204	210	205
rect	209	206	210	207
rect	209	207	210	208
rect	209	209	210	210
rect	209	210	210	211
rect	209	212	210	213
rect	209	213	210	214
rect	209	215	210	216
rect	209	216	210	217
rect	209	218	210	219
rect	209	219	210	220
rect	209	221	210	222
rect	209	222	210	223
rect	209	224	210	225
rect	209	225	210	226
rect	209	227	210	228
rect	209	228	210	229
rect	209	230	210	231
rect	209	231	210	232
rect	209	233	210	234
rect	209	234	210	235
rect	209	236	210	237
rect	209	237	210	238
rect	209	239	210	240
rect	209	240	210	241
rect	209	242	210	243
rect	209	243	210	244
rect	209	245	210	246
rect	209	246	210	247
rect	209	248	210	249
rect	209	249	210	250
rect	209	251	210	252
rect	209	252	210	253
rect	209	253	210	254
rect	209	254	210	255
rect	209	255	210	256
rect	209	257	210	258
rect	209	258	210	259
rect	209	260	210	261
rect	209	261	210	262
rect	209	262	210	263
rect	209	263	210	264
rect	209	264	210	265
rect	209	266	210	267
rect	209	267	210	268
rect	209	269	210	270
rect	209	270	210	271
rect	209	272	210	273
rect	209	273	210	274
rect	209	275	210	276
rect	209	276	210	277
rect	209	278	210	279
rect	209	279	210	280
rect	209	280	210	281
rect	209	281	210	282
rect	209	282	210	283
rect	209	284	210	285
rect	209	285	210	286
rect	209	287	210	288
rect	209	288	210	289
rect	209	289	210	290
rect	209	290	210	291
rect	209	291	210	292
rect	209	293	210	294
rect	209	294	210	295
rect	209	295	210	296
rect	209	296	210	297
rect	209	297	210	298
rect	209	298	210	299
rect	209	299	210	300
rect	209	300	210	301
rect	209	301	210	302
rect	209	302	210	303
rect	209	303	210	304
rect	209	304	210	305
rect	209	305	210	306
rect	209	306	210	307
rect	209	308	210	309
rect	209	309	210	310
rect	209	311	210	312
rect	209	312	210	313
rect	209	313	210	314
rect	209	314	210	315
rect	209	315	210	316
rect	209	317	210	318
rect	209	318	210	319
rect	209	319	210	320
rect	209	320	210	321
rect	209	321	210	322
rect	209	322	210	323
rect	209	323	210	324
rect	209	324	210	325
rect	209	325	210	326
rect	209	326	210	327
rect	209	327	210	328
rect	209	328	210	329
rect	209	329	210	330
rect	209	330	210	331
rect	209	331	210	332
rect	209	332	210	333
rect	209	333	210	334
rect	209	334	210	335
rect	209	335	210	336
rect	209	336	210	337
rect	209	337	210	338
rect	209	338	210	339
rect	209	339	210	340
rect	209	340	210	341
rect	209	341	210	342
rect	209	342	210	343
rect	209	343	210	344
rect	209	344	210	345
rect	209	345	210	346
rect	209	346	210	347
rect	209	347	210	348
rect	211	0	212	1
rect	211	1	212	2
rect	211	2	212	3
rect	211	3	212	4
rect	211	4	212	5
rect	211	5	212	6
rect	211	6	212	7
rect	211	8	212	9
rect	211	9	212	10
rect	211	11	212	12
rect	211	12	212	13
rect	211	14	212	15
rect	211	15	212	16
rect	211	17	212	18
rect	211	18	212	19
rect	211	20	212	21
rect	211	21	212	22
rect	211	23	212	24
rect	211	24	212	25
rect	211	26	212	27
rect	211	27	212	28
rect	211	29	212	30
rect	211	30	212	31
rect	211	32	212	33
rect	211	33	212	34
rect	211	35	212	36
rect	211	36	212	37
rect	211	38	212	39
rect	211	39	212	40
rect	211	41	212	42
rect	211	42	212	43
rect	211	44	212	45
rect	211	45	212	46
rect	211	47	212	48
rect	211	48	212	49
rect	211	50	212	51
rect	211	51	212	52
rect	211	53	212	54
rect	211	54	212	55
rect	211	56	212	57
rect	211	57	212	58
rect	211	59	212	60
rect	211	60	212	61
rect	211	62	212	63
rect	211	63	212	64
rect	211	65	212	66
rect	211	66	212	67
rect	211	68	212	69
rect	211	69	212	70
rect	211	71	212	72
rect	211	72	212	73
rect	211	74	212	75
rect	211	75	212	76
rect	211	77	212	78
rect	211	78	212	79
rect	211	80	212	81
rect	211	81	212	82
rect	211	83	212	84
rect	211	84	212	85
rect	211	86	212	87
rect	211	87	212	88
rect	211	89	212	90
rect	211	90	212	91
rect	211	92	212	93
rect	211	93	212	94
rect	211	95	212	96
rect	211	96	212	97
rect	211	98	212	99
rect	211	99	212	100
rect	211	101	212	102
rect	211	102	212	103
rect	211	104	212	105
rect	211	105	212	106
rect	211	107	212	108
rect	211	108	212	109
rect	211	110	212	111
rect	211	111	212	112
rect	211	113	212	114
rect	211	114	212	115
rect	211	116	212	117
rect	211	117	212	118
rect	211	119	212	120
rect	211	120	212	121
rect	211	122	212	123
rect	211	123	212	124
rect	211	125	212	126
rect	211	126	212	127
rect	211	128	212	129
rect	211	129	212	130
rect	211	131	212	132
rect	211	132	212	133
rect	211	134	212	135
rect	211	135	212	136
rect	211	137	212	138
rect	211	138	212	139
rect	211	140	212	141
rect	211	141	212	142
rect	211	143	212	144
rect	211	144	212	145
rect	211	146	212	147
rect	211	147	212	148
rect	211	149	212	150
rect	211	150	212	151
rect	211	152	212	153
rect	211	153	212	154
rect	211	155	212	156
rect	211	156	212	157
rect	211	158	212	159
rect	211	159	212	160
rect	211	161	212	162
rect	211	162	212	163
rect	211	164	212	165
rect	211	165	212	166
rect	211	167	212	168
rect	211	168	212	169
rect	211	170	212	171
rect	211	171	212	172
rect	211	173	212	174
rect	211	174	212	175
rect	211	176	212	177
rect	211	177	212	178
rect	211	179	212	180
rect	211	180	212	181
rect	211	182	212	183
rect	211	183	212	184
rect	211	185	212	186
rect	211	186	212	187
rect	211	188	212	189
rect	211	189	212	190
rect	211	191	212	192
rect	211	192	212	193
rect	211	194	212	195
rect	211	195	212	196
rect	211	197	212	198
rect	211	198	212	199
rect	211	200	212	201
rect	211	201	212	202
rect	211	203	212	204
rect	211	204	212	205
rect	211	206	212	207
rect	211	207	212	208
rect	211	209	212	210
rect	211	210	212	211
rect	211	212	212	213
rect	211	213	212	214
rect	211	215	212	216
rect	211	216	212	217
rect	211	218	212	219
rect	211	219	212	220
rect	211	221	212	222
rect	211	222	212	223
rect	211	224	212	225
rect	211	225	212	226
rect	211	227	212	228
rect	211	228	212	229
rect	211	230	212	231
rect	211	231	212	232
rect	211	233	212	234
rect	211	234	212	235
rect	211	236	212	237
rect	211	237	212	238
rect	211	239	212	240
rect	211	240	212	241
rect	211	242	212	243
rect	211	243	212	244
rect	211	245	212	246
rect	211	246	212	247
rect	211	248	212	249
rect	211	249	212	250
rect	211	251	212	252
rect	211	252	212	253
rect	211	253	212	254
rect	211	254	212	255
rect	211	255	212	256
rect	211	257	212	258
rect	211	258	212	259
rect	211	260	212	261
rect	211	261	212	262
rect	211	262	212	263
rect	211	263	212	264
rect	211	264	212	265
rect	211	266	212	267
rect	211	267	212	268
rect	211	269	212	270
rect	211	270	212	271
rect	211	272	212	273
rect	211	273	212	274
rect	211	275	212	276
rect	211	276	212	277
rect	211	278	212	279
rect	211	279	212	280
rect	211	280	212	281
rect	211	281	212	282
rect	211	282	212	283
rect	211	284	212	285
rect	211	285	212	286
rect	211	287	212	288
rect	211	288	212	289
rect	211	289	212	290
rect	211	290	212	291
rect	211	291	212	292
rect	211	293	212	294
rect	211	294	212	295
rect	211	295	212	296
rect	211	296	212	297
rect	211	297	212	298
rect	211	298	212	299
rect	211	299	212	300
rect	211	300	212	301
rect	211	301	212	302
rect	211	302	212	303
rect	211	303	212	304
rect	211	304	212	305
rect	211	305	212	306
rect	211	306	212	307
rect	211	308	212	309
rect	211	309	212	310
rect	211	311	212	312
rect	211	312	212	313
rect	211	313	212	314
rect	211	314	212	315
rect	211	315	212	316
rect	211	317	212	318
rect	211	318	212	319
rect	211	319	212	320
rect	211	320	212	321
rect	212	0	213	1
rect	212	1	213	2
rect	212	2	213	3
rect	212	3	213	4
rect	212	4	213	5
rect	212	5	213	6
rect	212	6	213	7
rect	212	8	213	9
rect	212	9	213	10
rect	212	11	213	12
rect	212	12	213	13
rect	212	14	213	15
rect	212	15	213	16
rect	212	17	213	18
rect	212	18	213	19
rect	212	20	213	21
rect	212	21	213	22
rect	212	23	213	24
rect	212	24	213	25
rect	212	26	213	27
rect	212	27	213	28
rect	212	29	213	30
rect	212	30	213	31
rect	212	32	213	33
rect	212	33	213	34
rect	212	35	213	36
rect	212	36	213	37
rect	212	38	213	39
rect	212	39	213	40
rect	212	41	213	42
rect	212	42	213	43
rect	212	44	213	45
rect	212	45	213	46
rect	212	47	213	48
rect	212	48	213	49
rect	212	50	213	51
rect	212	51	213	52
rect	212	53	213	54
rect	212	54	213	55
rect	212	56	213	57
rect	212	57	213	58
rect	212	59	213	60
rect	212	60	213	61
rect	212	62	213	63
rect	212	63	213	64
rect	212	65	213	66
rect	212	66	213	67
rect	212	68	213	69
rect	212	69	213	70
rect	212	71	213	72
rect	212	72	213	73
rect	212	74	213	75
rect	212	75	213	76
rect	212	77	213	78
rect	212	78	213	79
rect	212	80	213	81
rect	212	81	213	82
rect	212	83	213	84
rect	212	84	213	85
rect	212	86	213	87
rect	212	87	213	88
rect	212	89	213	90
rect	212	90	213	91
rect	212	92	213	93
rect	212	93	213	94
rect	212	95	213	96
rect	212	96	213	97
rect	212	98	213	99
rect	212	99	213	100
rect	212	101	213	102
rect	212	102	213	103
rect	212	104	213	105
rect	212	105	213	106
rect	212	107	213	108
rect	212	108	213	109
rect	212	110	213	111
rect	212	111	213	112
rect	212	113	213	114
rect	212	114	213	115
rect	212	116	213	117
rect	212	117	213	118
rect	212	119	213	120
rect	212	120	213	121
rect	212	122	213	123
rect	212	123	213	124
rect	212	125	213	126
rect	212	126	213	127
rect	212	128	213	129
rect	212	129	213	130
rect	212	131	213	132
rect	212	132	213	133
rect	212	134	213	135
rect	212	135	213	136
rect	212	137	213	138
rect	212	138	213	139
rect	212	140	213	141
rect	212	141	213	142
rect	212	143	213	144
rect	212	144	213	145
rect	212	146	213	147
rect	212	147	213	148
rect	212	149	213	150
rect	212	150	213	151
rect	212	152	213	153
rect	212	153	213	154
rect	212	155	213	156
rect	212	156	213	157
rect	212	158	213	159
rect	212	159	213	160
rect	212	161	213	162
rect	212	162	213	163
rect	212	164	213	165
rect	212	165	213	166
rect	212	167	213	168
rect	212	168	213	169
rect	212	170	213	171
rect	212	171	213	172
rect	212	173	213	174
rect	212	174	213	175
rect	212	176	213	177
rect	212	177	213	178
rect	212	179	213	180
rect	212	180	213	181
rect	212	182	213	183
rect	212	183	213	184
rect	212	185	213	186
rect	212	186	213	187
rect	212	188	213	189
rect	212	189	213	190
rect	212	191	213	192
rect	212	192	213	193
rect	212	194	213	195
rect	212	195	213	196
rect	212	197	213	198
rect	212	198	213	199
rect	212	200	213	201
rect	212	201	213	202
rect	212	203	213	204
rect	212	204	213	205
rect	212	206	213	207
rect	212	207	213	208
rect	212	209	213	210
rect	212	210	213	211
rect	212	212	213	213
rect	212	213	213	214
rect	212	215	213	216
rect	212	216	213	217
rect	212	218	213	219
rect	212	219	213	220
rect	212	221	213	222
rect	212	222	213	223
rect	212	224	213	225
rect	212	225	213	226
rect	212	227	213	228
rect	212	228	213	229
rect	212	230	213	231
rect	212	231	213	232
rect	212	233	213	234
rect	212	234	213	235
rect	212	236	213	237
rect	212	237	213	238
rect	212	239	213	240
rect	212	240	213	241
rect	212	242	213	243
rect	212	243	213	244
rect	212	245	213	246
rect	212	246	213	247
rect	212	248	213	249
rect	212	249	213	250
rect	212	251	213	252
rect	212	252	213	253
rect	212	253	213	254
rect	212	254	213	255
rect	212	255	213	256
rect	212	257	213	258
rect	212	258	213	259
rect	212	260	213	261
rect	212	261	213	262
rect	212	262	213	263
rect	212	263	213	264
rect	212	264	213	265
rect	212	266	213	267
rect	212	267	213	268
rect	212	269	213	270
rect	212	270	213	271
rect	212	272	213	273
rect	212	273	213	274
rect	212	275	213	276
rect	212	276	213	277
rect	212	278	213	279
rect	212	279	213	280
rect	212	280	213	281
rect	212	281	213	282
rect	212	282	213	283
rect	212	284	213	285
rect	212	285	213	286
rect	212	287	213	288
rect	212	288	213	289
rect	212	289	213	290
rect	212	290	213	291
rect	212	291	213	292
rect	212	293	213	294
rect	212	294	213	295
rect	212	295	213	296
rect	212	296	213	297
rect	212	297	213	298
rect	212	298	213	299
rect	212	299	213	300
rect	212	300	213	301
rect	212	301	213	302
rect	212	302	213	303
rect	212	303	213	304
rect	212	304	213	305
rect	212	305	213	306
rect	212	306	213	307
rect	212	308	213	309
rect	212	309	213	310
rect	212	311	213	312
rect	212	312	213	313
rect	212	313	213	314
rect	212	314	213	315
rect	212	315	213	316
rect	212	317	213	318
rect	212	318	213	319
rect	212	319	213	320
rect	212	320	213	321
rect	213	0	214	1
rect	213	1	214	2
rect	213	2	214	3
rect	213	3	214	4
rect	213	4	214	5
rect	213	5	214	6
rect	213	6	214	7
rect	213	8	214	9
rect	213	9	214	10
rect	213	11	214	12
rect	213	12	214	13
rect	213	14	214	15
rect	213	15	214	16
rect	213	17	214	18
rect	213	18	214	19
rect	213	20	214	21
rect	213	21	214	22
rect	213	23	214	24
rect	213	24	214	25
rect	213	26	214	27
rect	213	27	214	28
rect	213	29	214	30
rect	213	30	214	31
rect	213	32	214	33
rect	213	33	214	34
rect	213	35	214	36
rect	213	36	214	37
rect	213	38	214	39
rect	213	39	214	40
rect	213	41	214	42
rect	213	42	214	43
rect	213	44	214	45
rect	213	45	214	46
rect	213	47	214	48
rect	213	48	214	49
rect	213	50	214	51
rect	213	51	214	52
rect	213	53	214	54
rect	213	54	214	55
rect	213	56	214	57
rect	213	57	214	58
rect	213	59	214	60
rect	213	60	214	61
rect	213	62	214	63
rect	213	63	214	64
rect	213	65	214	66
rect	213	66	214	67
rect	213	68	214	69
rect	213	69	214	70
rect	213	71	214	72
rect	213	72	214	73
rect	213	74	214	75
rect	213	75	214	76
rect	213	77	214	78
rect	213	78	214	79
rect	213	80	214	81
rect	213	81	214	82
rect	213	83	214	84
rect	213	84	214	85
rect	213	86	214	87
rect	213	87	214	88
rect	213	89	214	90
rect	213	90	214	91
rect	213	92	214	93
rect	213	93	214	94
rect	213	95	214	96
rect	213	96	214	97
rect	213	98	214	99
rect	213	99	214	100
rect	213	101	214	102
rect	213	102	214	103
rect	213	104	214	105
rect	213	105	214	106
rect	213	107	214	108
rect	213	108	214	109
rect	213	110	214	111
rect	213	111	214	112
rect	213	113	214	114
rect	213	114	214	115
rect	213	116	214	117
rect	213	117	214	118
rect	213	119	214	120
rect	213	120	214	121
rect	213	122	214	123
rect	213	123	214	124
rect	213	125	214	126
rect	213	126	214	127
rect	213	128	214	129
rect	213	129	214	130
rect	213	131	214	132
rect	213	132	214	133
rect	213	134	214	135
rect	213	135	214	136
rect	213	137	214	138
rect	213	138	214	139
rect	213	140	214	141
rect	213	141	214	142
rect	213	143	214	144
rect	213	144	214	145
rect	213	146	214	147
rect	213	147	214	148
rect	213	149	214	150
rect	213	150	214	151
rect	213	152	214	153
rect	213	153	214	154
rect	213	155	214	156
rect	213	156	214	157
rect	213	158	214	159
rect	213	159	214	160
rect	213	161	214	162
rect	213	162	214	163
rect	213	164	214	165
rect	213	165	214	166
rect	213	167	214	168
rect	213	168	214	169
rect	213	170	214	171
rect	213	171	214	172
rect	213	173	214	174
rect	213	174	214	175
rect	213	176	214	177
rect	213	177	214	178
rect	213	179	214	180
rect	213	180	214	181
rect	213	182	214	183
rect	213	183	214	184
rect	213	185	214	186
rect	213	186	214	187
rect	213	188	214	189
rect	213	189	214	190
rect	213	191	214	192
rect	213	192	214	193
rect	213	194	214	195
rect	213	195	214	196
rect	213	197	214	198
rect	213	198	214	199
rect	213	200	214	201
rect	213	201	214	202
rect	213	203	214	204
rect	213	204	214	205
rect	213	206	214	207
rect	213	207	214	208
rect	213	209	214	210
rect	213	210	214	211
rect	213	212	214	213
rect	213	213	214	214
rect	213	215	214	216
rect	213	216	214	217
rect	213	218	214	219
rect	213	219	214	220
rect	213	221	214	222
rect	213	222	214	223
rect	213	224	214	225
rect	213	225	214	226
rect	213	227	214	228
rect	213	228	214	229
rect	213	230	214	231
rect	213	231	214	232
rect	213	233	214	234
rect	213	234	214	235
rect	213	236	214	237
rect	213	237	214	238
rect	213	239	214	240
rect	213	240	214	241
rect	213	242	214	243
rect	213	243	214	244
rect	213	245	214	246
rect	213	246	214	247
rect	213	248	214	249
rect	213	249	214	250
rect	213	251	214	252
rect	213	252	214	253
rect	213	253	214	254
rect	213	254	214	255
rect	213	255	214	256
rect	213	257	214	258
rect	213	258	214	259
rect	213	260	214	261
rect	213	261	214	262
rect	213	262	214	263
rect	213	263	214	264
rect	213	264	214	265
rect	213	266	214	267
rect	213	267	214	268
rect	213	269	214	270
rect	213	270	214	271
rect	213	272	214	273
rect	213	273	214	274
rect	213	275	214	276
rect	213	276	214	277
rect	213	278	214	279
rect	213	279	214	280
rect	213	280	214	281
rect	213	281	214	282
rect	213	282	214	283
rect	213	284	214	285
rect	213	285	214	286
rect	213	287	214	288
rect	213	288	214	289
rect	213	289	214	290
rect	213	290	214	291
rect	213	291	214	292
rect	213	293	214	294
rect	213	294	214	295
rect	213	295	214	296
rect	213	296	214	297
rect	213	297	214	298
rect	213	298	214	299
rect	213	299	214	300
rect	213	300	214	301
rect	213	301	214	302
rect	213	302	214	303
rect	213	303	214	304
rect	213	304	214	305
rect	213	305	214	306
rect	213	306	214	307
rect	213	308	214	309
rect	213	309	214	310
rect	213	311	214	312
rect	213	312	214	313
rect	213	313	214	314
rect	213	314	214	315
rect	213	315	214	316
rect	213	317	214	318
rect	213	318	214	319
rect	213	319	214	320
rect	213	320	214	321
rect	214	0	215	1
rect	214	1	215	2
rect	214	2	215	3
rect	214	3	215	4
rect	214	4	215	5
rect	214	5	215	6
rect	214	6	215	7
rect	214	8	215	9
rect	214	9	215	10
rect	214	11	215	12
rect	214	12	215	13
rect	214	14	215	15
rect	214	15	215	16
rect	214	17	215	18
rect	214	18	215	19
rect	214	20	215	21
rect	214	21	215	22
rect	214	23	215	24
rect	214	24	215	25
rect	214	26	215	27
rect	214	27	215	28
rect	214	29	215	30
rect	214	30	215	31
rect	214	32	215	33
rect	214	33	215	34
rect	214	35	215	36
rect	214	36	215	37
rect	214	38	215	39
rect	214	39	215	40
rect	214	41	215	42
rect	214	42	215	43
rect	214	44	215	45
rect	214	45	215	46
rect	214	47	215	48
rect	214	48	215	49
rect	214	50	215	51
rect	214	51	215	52
rect	214	53	215	54
rect	214	54	215	55
rect	214	56	215	57
rect	214	57	215	58
rect	214	59	215	60
rect	214	60	215	61
rect	214	62	215	63
rect	214	63	215	64
rect	214	65	215	66
rect	214	66	215	67
rect	214	68	215	69
rect	214	69	215	70
rect	214	71	215	72
rect	214	72	215	73
rect	214	74	215	75
rect	214	75	215	76
rect	214	77	215	78
rect	214	78	215	79
rect	214	80	215	81
rect	214	81	215	82
rect	214	83	215	84
rect	214	84	215	85
rect	214	86	215	87
rect	214	87	215	88
rect	214	89	215	90
rect	214	90	215	91
rect	214	92	215	93
rect	214	93	215	94
rect	214	95	215	96
rect	214	96	215	97
rect	214	98	215	99
rect	214	99	215	100
rect	214	101	215	102
rect	214	102	215	103
rect	214	104	215	105
rect	214	105	215	106
rect	214	107	215	108
rect	214	108	215	109
rect	214	110	215	111
rect	214	111	215	112
rect	214	113	215	114
rect	214	114	215	115
rect	214	116	215	117
rect	214	117	215	118
rect	214	119	215	120
rect	214	120	215	121
rect	214	122	215	123
rect	214	123	215	124
rect	214	125	215	126
rect	214	126	215	127
rect	214	128	215	129
rect	214	129	215	130
rect	214	131	215	132
rect	214	132	215	133
rect	214	134	215	135
rect	214	135	215	136
rect	214	137	215	138
rect	214	138	215	139
rect	214	140	215	141
rect	214	141	215	142
rect	214	143	215	144
rect	214	144	215	145
rect	214	146	215	147
rect	214	147	215	148
rect	214	149	215	150
rect	214	150	215	151
rect	214	152	215	153
rect	214	153	215	154
rect	214	155	215	156
rect	214	156	215	157
rect	214	158	215	159
rect	214	159	215	160
rect	214	161	215	162
rect	214	162	215	163
rect	214	164	215	165
rect	214	165	215	166
rect	214	167	215	168
rect	214	168	215	169
rect	214	170	215	171
rect	214	171	215	172
rect	214	173	215	174
rect	214	174	215	175
rect	214	176	215	177
rect	214	177	215	178
rect	214	179	215	180
rect	214	180	215	181
rect	214	182	215	183
rect	214	183	215	184
rect	214	185	215	186
rect	214	186	215	187
rect	214	188	215	189
rect	214	189	215	190
rect	214	191	215	192
rect	214	192	215	193
rect	214	194	215	195
rect	214	195	215	196
rect	214	197	215	198
rect	214	198	215	199
rect	214	200	215	201
rect	214	201	215	202
rect	214	203	215	204
rect	214	204	215	205
rect	214	206	215	207
rect	214	207	215	208
rect	214	209	215	210
rect	214	210	215	211
rect	214	212	215	213
rect	214	213	215	214
rect	214	215	215	216
rect	214	216	215	217
rect	214	218	215	219
rect	214	219	215	220
rect	214	221	215	222
rect	214	222	215	223
rect	214	224	215	225
rect	214	225	215	226
rect	214	227	215	228
rect	214	228	215	229
rect	214	230	215	231
rect	214	231	215	232
rect	214	233	215	234
rect	214	234	215	235
rect	214	236	215	237
rect	214	237	215	238
rect	214	239	215	240
rect	214	240	215	241
rect	214	242	215	243
rect	214	243	215	244
rect	214	245	215	246
rect	214	246	215	247
rect	214	248	215	249
rect	214	249	215	250
rect	214	251	215	252
rect	214	252	215	253
rect	214	253	215	254
rect	214	254	215	255
rect	214	255	215	256
rect	214	257	215	258
rect	214	258	215	259
rect	214	260	215	261
rect	214	261	215	262
rect	214	262	215	263
rect	214	263	215	264
rect	214	264	215	265
rect	214	266	215	267
rect	214	267	215	268
rect	214	269	215	270
rect	214	270	215	271
rect	214	272	215	273
rect	214	273	215	274
rect	214	275	215	276
rect	214	276	215	277
rect	214	278	215	279
rect	214	279	215	280
rect	214	280	215	281
rect	214	281	215	282
rect	214	282	215	283
rect	214	284	215	285
rect	214	285	215	286
rect	214	287	215	288
rect	214	288	215	289
rect	214	289	215	290
rect	214	290	215	291
rect	214	291	215	292
rect	214	293	215	294
rect	214	294	215	295
rect	214	295	215	296
rect	214	296	215	297
rect	214	297	215	298
rect	214	298	215	299
rect	214	299	215	300
rect	214	300	215	301
rect	214	301	215	302
rect	214	302	215	303
rect	214	303	215	304
rect	214	304	215	305
rect	214	305	215	306
rect	214	306	215	307
rect	214	308	215	309
rect	214	309	215	310
rect	214	311	215	312
rect	214	312	215	313
rect	214	313	215	314
rect	214	314	215	315
rect	214	315	215	316
rect	214	317	215	318
rect	214	318	215	319
rect	214	319	215	320
rect	214	320	215	321
rect	215	0	216	1
rect	215	1	216	2
rect	215	2	216	3
rect	215	3	216	4
rect	215	4	216	5
rect	215	5	216	6
rect	215	6	216	7
rect	215	8	216	9
rect	215	9	216	10
rect	215	11	216	12
rect	215	12	216	13
rect	215	14	216	15
rect	215	15	216	16
rect	215	17	216	18
rect	215	18	216	19
rect	215	20	216	21
rect	215	21	216	22
rect	215	23	216	24
rect	215	24	216	25
rect	215	26	216	27
rect	215	27	216	28
rect	215	29	216	30
rect	215	30	216	31
rect	215	32	216	33
rect	215	33	216	34
rect	215	35	216	36
rect	215	36	216	37
rect	215	38	216	39
rect	215	39	216	40
rect	215	41	216	42
rect	215	42	216	43
rect	215	44	216	45
rect	215	45	216	46
rect	215	47	216	48
rect	215	48	216	49
rect	215	50	216	51
rect	215	51	216	52
rect	215	53	216	54
rect	215	54	216	55
rect	215	56	216	57
rect	215	57	216	58
rect	215	59	216	60
rect	215	60	216	61
rect	215	62	216	63
rect	215	63	216	64
rect	215	65	216	66
rect	215	66	216	67
rect	215	68	216	69
rect	215	69	216	70
rect	215	71	216	72
rect	215	72	216	73
rect	215	74	216	75
rect	215	75	216	76
rect	215	77	216	78
rect	215	78	216	79
rect	215	80	216	81
rect	215	81	216	82
rect	215	83	216	84
rect	215	84	216	85
rect	215	86	216	87
rect	215	87	216	88
rect	215	89	216	90
rect	215	90	216	91
rect	215	92	216	93
rect	215	93	216	94
rect	215	95	216	96
rect	215	96	216	97
rect	215	98	216	99
rect	215	99	216	100
rect	215	101	216	102
rect	215	102	216	103
rect	215	104	216	105
rect	215	105	216	106
rect	215	107	216	108
rect	215	108	216	109
rect	215	110	216	111
rect	215	111	216	112
rect	215	113	216	114
rect	215	114	216	115
rect	215	116	216	117
rect	215	117	216	118
rect	215	119	216	120
rect	215	120	216	121
rect	215	122	216	123
rect	215	123	216	124
rect	215	125	216	126
rect	215	126	216	127
rect	215	128	216	129
rect	215	129	216	130
rect	215	131	216	132
rect	215	132	216	133
rect	215	134	216	135
rect	215	135	216	136
rect	215	137	216	138
rect	215	138	216	139
rect	215	140	216	141
rect	215	141	216	142
rect	215	143	216	144
rect	215	144	216	145
rect	215	146	216	147
rect	215	147	216	148
rect	215	149	216	150
rect	215	150	216	151
rect	215	152	216	153
rect	215	153	216	154
rect	215	155	216	156
rect	215	156	216	157
rect	215	158	216	159
rect	215	159	216	160
rect	215	161	216	162
rect	215	162	216	163
rect	215	164	216	165
rect	215	165	216	166
rect	215	167	216	168
rect	215	168	216	169
rect	215	170	216	171
rect	215	171	216	172
rect	215	173	216	174
rect	215	174	216	175
rect	215	176	216	177
rect	215	177	216	178
rect	215	179	216	180
rect	215	180	216	181
rect	215	182	216	183
rect	215	183	216	184
rect	215	185	216	186
rect	215	186	216	187
rect	215	188	216	189
rect	215	189	216	190
rect	215	191	216	192
rect	215	192	216	193
rect	215	194	216	195
rect	215	195	216	196
rect	215	197	216	198
rect	215	198	216	199
rect	215	200	216	201
rect	215	201	216	202
rect	215	203	216	204
rect	215	204	216	205
rect	215	206	216	207
rect	215	207	216	208
rect	215	209	216	210
rect	215	210	216	211
rect	215	212	216	213
rect	215	213	216	214
rect	215	215	216	216
rect	215	216	216	217
rect	215	218	216	219
rect	215	219	216	220
rect	215	221	216	222
rect	215	222	216	223
rect	215	224	216	225
rect	215	225	216	226
rect	215	227	216	228
rect	215	228	216	229
rect	215	230	216	231
rect	215	231	216	232
rect	215	233	216	234
rect	215	234	216	235
rect	215	236	216	237
rect	215	237	216	238
rect	215	239	216	240
rect	215	240	216	241
rect	215	242	216	243
rect	215	243	216	244
rect	215	245	216	246
rect	215	246	216	247
rect	215	248	216	249
rect	215	249	216	250
rect	215	251	216	252
rect	215	252	216	253
rect	215	253	216	254
rect	215	254	216	255
rect	215	255	216	256
rect	215	257	216	258
rect	215	258	216	259
rect	215	260	216	261
rect	215	261	216	262
rect	215	262	216	263
rect	215	263	216	264
rect	215	264	216	265
rect	215	266	216	267
rect	215	267	216	268
rect	215	269	216	270
rect	215	270	216	271
rect	215	272	216	273
rect	215	273	216	274
rect	215	275	216	276
rect	215	276	216	277
rect	215	278	216	279
rect	215	279	216	280
rect	215	280	216	281
rect	215	281	216	282
rect	215	282	216	283
rect	215	283	216	284
rect	215	284	216	285
rect	215	285	216	286
rect	215	286	216	287
rect	215	287	216	288
rect	215	288	216	289
rect	215	289	216	290
rect	215	290	216	291
rect	215	291	216	292
rect	215	293	216	294
rect	215	294	216	295
rect	215	295	216	296
rect	215	296	216	297
rect	215	297	216	298
rect	215	298	216	299
rect	215	299	216	300
rect	215	300	216	301
rect	215	301	216	302
rect	215	302	216	303
rect	215	303	216	304
rect	215	304	216	305
rect	215	305	216	306
rect	215	306	216	307
rect	215	308	216	309
rect	215	309	216	310
rect	215	310	216	311
rect	215	311	216	312
rect	215	312	216	313
rect	215	313	216	314
rect	215	314	216	315
rect	215	315	216	316
rect	215	316	216	317
rect	215	317	216	318
rect	215	318	216	319
rect	215	319	216	320
rect	215	320	216	321
rect	220	0	221	1
rect	220	1	221	2
rect	220	2	221	3
rect	220	3	221	4
rect	220	4	221	5
rect	220	5	221	6
rect	220	6	221	7
rect	220	8	221	9
rect	220	9	221	10
rect	220	11	221	12
rect	220	12	221	13
rect	220	14	221	15
rect	220	15	221	16
rect	220	17	221	18
rect	220	18	221	19
rect	220	20	221	21
rect	220	21	221	22
rect	220	23	221	24
rect	220	24	221	25
rect	220	26	221	27
rect	220	27	221	28
rect	220	29	221	30
rect	220	30	221	31
rect	220	32	221	33
rect	220	33	221	34
rect	220	35	221	36
rect	220	36	221	37
rect	220	38	221	39
rect	220	39	221	40
rect	220	41	221	42
rect	220	42	221	43
rect	220	44	221	45
rect	220	45	221	46
rect	220	47	221	48
rect	220	48	221	49
rect	220	50	221	51
rect	220	51	221	52
rect	220	53	221	54
rect	220	54	221	55
rect	220	56	221	57
rect	220	57	221	58
rect	220	59	221	60
rect	220	60	221	61
rect	220	62	221	63
rect	220	63	221	64
rect	220	65	221	66
rect	220	66	221	67
rect	220	68	221	69
rect	220	69	221	70
rect	220	71	221	72
rect	220	72	221	73
rect	220	74	221	75
rect	220	75	221	76
rect	220	77	221	78
rect	220	78	221	79
rect	220	80	221	81
rect	220	81	221	82
rect	220	83	221	84
rect	220	84	221	85
rect	220	86	221	87
rect	220	87	221	88
rect	220	89	221	90
rect	220	90	221	91
rect	220	92	221	93
rect	220	93	221	94
rect	220	95	221	96
rect	220	96	221	97
rect	220	98	221	99
rect	220	99	221	100
rect	220	101	221	102
rect	220	102	221	103
rect	220	104	221	105
rect	220	105	221	106
rect	220	107	221	108
rect	220	108	221	109
rect	220	110	221	111
rect	220	111	221	112
rect	220	113	221	114
rect	220	114	221	115
rect	220	116	221	117
rect	220	117	221	118
rect	220	119	221	120
rect	220	120	221	121
rect	220	122	221	123
rect	220	123	221	124
rect	220	125	221	126
rect	220	126	221	127
rect	220	128	221	129
rect	220	129	221	130
rect	220	131	221	132
rect	220	132	221	133
rect	220	134	221	135
rect	220	135	221	136
rect	220	137	221	138
rect	220	138	221	139
rect	220	140	221	141
rect	220	141	221	142
rect	220	143	221	144
rect	220	144	221	145
rect	220	146	221	147
rect	220	147	221	148
rect	220	149	221	150
rect	220	150	221	151
rect	220	152	221	153
rect	220	153	221	154
rect	220	155	221	156
rect	220	156	221	157
rect	220	158	221	159
rect	220	159	221	160
rect	220	161	221	162
rect	220	162	221	163
rect	220	164	221	165
rect	220	165	221	166
rect	220	167	221	168
rect	220	168	221	169
rect	220	170	221	171
rect	220	171	221	172
rect	220	173	221	174
rect	220	174	221	175
rect	220	176	221	177
rect	220	177	221	178
rect	220	179	221	180
rect	220	180	221	181
rect	220	182	221	183
rect	220	183	221	184
rect	220	185	221	186
rect	220	186	221	187
rect	220	188	221	189
rect	220	189	221	190
rect	220	191	221	192
rect	220	192	221	193
rect	220	194	221	195
rect	220	195	221	196
rect	220	197	221	198
rect	220	198	221	199
rect	220	200	221	201
rect	220	201	221	202
rect	220	203	221	204
rect	220	204	221	205
rect	220	206	221	207
rect	220	207	221	208
rect	220	209	221	210
rect	220	210	221	211
rect	220	212	221	213
rect	220	213	221	214
rect	220	215	221	216
rect	220	216	221	217
rect	220	218	221	219
rect	220	219	221	220
rect	220	221	221	222
rect	220	222	221	223
rect	220	224	221	225
rect	220	225	221	226
rect	220	227	221	228
rect	220	228	221	229
rect	220	230	221	231
rect	220	231	221	232
rect	220	233	221	234
rect	220	234	221	235
rect	220	236	221	237
rect	220	237	221	238
rect	220	239	221	240
rect	220	240	221	241
rect	220	242	221	243
rect	220	243	221	244
rect	220	245	221	246
rect	220	246	221	247
rect	220	248	221	249
rect	220	249	221	250
rect	220	251	221	252
rect	220	252	221	253
rect	220	253	221	254
rect	220	254	221	255
rect	220	255	221	256
rect	220	257	221	258
rect	220	258	221	259
rect	220	260	221	261
rect	220	261	221	262
rect	220	262	221	263
rect	220	263	221	264
rect	220	264	221	265
rect	220	266	221	267
rect	220	267	221	268
rect	220	268	221	269
rect	220	269	221	270
rect	220	270	221	271
rect	220	271	221	272
rect	220	272	221	273
rect	220	273	221	274
rect	220	275	221	276
rect	220	276	221	277
rect	220	278	221	279
rect	220	279	221	280
rect	220	280	221	281
rect	220	281	221	282
rect	220	282	221	283
rect	220	283	221	284
rect	220	284	221	285
rect	220	285	221	286
rect	220	286	221	287
rect	220	287	221	288
rect	220	288	221	289
rect	220	289	221	290
rect	220	290	221	291
rect	220	291	221	292
rect	220	292	221	293
rect	220	293	221	294
rect	220	294	221	295
rect	220	295	221	296
rect	220	296	221	297
rect	220	297	221	298
rect	220	298	221	299
rect	220	299	221	300
rect	220	300	221	301
rect	220	301	221	302
rect	220	302	221	303
rect	220	303	221	304
rect	220	304	221	305
rect	220	305	221	306
rect	220	306	221	307
rect	220	307	221	308
rect	220	308	221	309
rect	220	309	221	310
rect	220	310	221	311
rect	220	311	221	312
rect	220	312	221	313
rect	220	313	221	314
rect	220	314	221	315
rect	220	315	221	316
rect	220	316	221	317
rect	220	317	221	318
rect	220	318	221	319
rect	220	319	221	320
rect	220	320	221	321
rect	222	0	223	1
rect	222	1	223	2
rect	222	2	223	3
rect	222	3	223	4
rect	222	4	223	5
rect	222	5	223	6
rect	222	6	223	7
rect	222	8	223	9
rect	222	9	223	10
rect	222	11	223	12
rect	222	12	223	13
rect	222	14	223	15
rect	222	15	223	16
rect	222	17	223	18
rect	222	18	223	19
rect	222	20	223	21
rect	222	21	223	22
rect	222	23	223	24
rect	222	24	223	25
rect	222	26	223	27
rect	222	27	223	28
rect	222	29	223	30
rect	222	30	223	31
rect	222	32	223	33
rect	222	33	223	34
rect	222	35	223	36
rect	222	36	223	37
rect	222	38	223	39
rect	222	39	223	40
rect	222	41	223	42
rect	222	42	223	43
rect	222	44	223	45
rect	222	45	223	46
rect	222	47	223	48
rect	222	48	223	49
rect	222	50	223	51
rect	222	51	223	52
rect	222	53	223	54
rect	222	54	223	55
rect	222	56	223	57
rect	222	57	223	58
rect	222	59	223	60
rect	222	60	223	61
rect	222	62	223	63
rect	222	63	223	64
rect	222	65	223	66
rect	222	66	223	67
rect	222	68	223	69
rect	222	69	223	70
rect	222	71	223	72
rect	222	72	223	73
rect	222	74	223	75
rect	222	75	223	76
rect	222	77	223	78
rect	222	78	223	79
rect	222	80	223	81
rect	222	81	223	82
rect	222	83	223	84
rect	222	84	223	85
rect	222	86	223	87
rect	222	87	223	88
rect	222	89	223	90
rect	222	90	223	91
rect	222	92	223	93
rect	222	93	223	94
rect	222	95	223	96
rect	222	96	223	97
rect	222	98	223	99
rect	222	99	223	100
rect	222	101	223	102
rect	222	102	223	103
rect	222	104	223	105
rect	222	105	223	106
rect	222	107	223	108
rect	222	108	223	109
rect	222	110	223	111
rect	222	111	223	112
rect	222	113	223	114
rect	222	114	223	115
rect	222	116	223	117
rect	222	117	223	118
rect	222	119	223	120
rect	222	120	223	121
rect	222	122	223	123
rect	222	123	223	124
rect	222	125	223	126
rect	222	126	223	127
rect	222	128	223	129
rect	222	129	223	130
rect	222	131	223	132
rect	222	132	223	133
rect	222	134	223	135
rect	222	135	223	136
rect	222	137	223	138
rect	222	138	223	139
rect	222	140	223	141
rect	222	141	223	142
rect	222	143	223	144
rect	222	144	223	145
rect	222	146	223	147
rect	222	147	223	148
rect	222	149	223	150
rect	222	150	223	151
rect	222	152	223	153
rect	222	153	223	154
rect	222	155	223	156
rect	222	156	223	157
rect	222	158	223	159
rect	222	159	223	160
rect	222	161	223	162
rect	222	162	223	163
rect	222	164	223	165
rect	222	165	223	166
rect	222	167	223	168
rect	222	168	223	169
rect	222	170	223	171
rect	222	171	223	172
rect	222	173	223	174
rect	222	174	223	175
rect	222	176	223	177
rect	222	177	223	178
rect	222	179	223	180
rect	222	180	223	181
rect	222	182	223	183
rect	222	183	223	184
rect	222	185	223	186
rect	222	186	223	187
rect	222	188	223	189
rect	222	189	223	190
rect	222	191	223	192
rect	222	192	223	193
rect	222	194	223	195
rect	222	195	223	196
rect	222	197	223	198
rect	222	198	223	199
rect	222	200	223	201
rect	222	201	223	202
rect	222	203	223	204
rect	222	204	223	205
rect	222	206	223	207
rect	222	207	223	208
rect	222	209	223	210
rect	222	210	223	211
rect	222	212	223	213
rect	222	213	223	214
rect	222	215	223	216
rect	222	216	223	217
rect	222	218	223	219
rect	222	219	223	220
rect	222	221	223	222
rect	222	222	223	223
rect	222	224	223	225
rect	222	225	223	226
rect	222	227	223	228
rect	222	228	223	229
rect	222	230	223	231
rect	222	231	223	232
rect	222	233	223	234
rect	222	234	223	235
rect	222	236	223	237
rect	222	237	223	238
rect	222	239	223	240
rect	222	240	223	241
rect	222	242	223	243
rect	222	243	223	244
rect	222	245	223	246
rect	222	246	223	247
rect	222	248	223	249
rect	222	249	223	250
rect	222	251	223	252
rect	222	252	223	253
rect	222	253	223	254
rect	222	254	223	255
rect	222	255	223	256
rect	222	257	223	258
rect	222	258	223	259
rect	222	260	223	261
rect	222	261	223	262
rect	222	262	223	263
rect	222	263	223	264
rect	222	264	223	265
rect	222	266	223	267
rect	222	267	223	268
rect	222	268	223	269
rect	222	269	223	270
rect	222	270	223	271
rect	222	271	223	272
rect	222	272	223	273
rect	222	273	223	274
rect	222	275	223	276
rect	222	276	223	277
rect	222	278	223	279
rect	222	279	223	280
rect	222	280	223	281
rect	222	281	223	282
rect	222	282	223	283
rect	222	283	223	284
rect	222	284	223	285
rect	222	285	223	286
rect	222	286	223	287
rect	222	287	223	288
rect	223	0	224	1
rect	223	1	224	2
rect	223	2	224	3
rect	223	3	224	4
rect	223	4	224	5
rect	223	5	224	6
rect	223	6	224	7
rect	223	8	224	9
rect	223	9	224	10
rect	223	11	224	12
rect	223	12	224	13
rect	223	14	224	15
rect	223	15	224	16
rect	223	17	224	18
rect	223	18	224	19
rect	223	20	224	21
rect	223	21	224	22
rect	223	23	224	24
rect	223	24	224	25
rect	223	26	224	27
rect	223	27	224	28
rect	223	29	224	30
rect	223	30	224	31
rect	223	32	224	33
rect	223	33	224	34
rect	223	35	224	36
rect	223	36	224	37
rect	223	38	224	39
rect	223	39	224	40
rect	223	41	224	42
rect	223	42	224	43
rect	223	44	224	45
rect	223	45	224	46
rect	223	47	224	48
rect	223	48	224	49
rect	223	50	224	51
rect	223	51	224	52
rect	223	53	224	54
rect	223	54	224	55
rect	223	56	224	57
rect	223	57	224	58
rect	223	59	224	60
rect	223	60	224	61
rect	223	62	224	63
rect	223	63	224	64
rect	223	65	224	66
rect	223	66	224	67
rect	223	68	224	69
rect	223	69	224	70
rect	223	71	224	72
rect	223	72	224	73
rect	223	74	224	75
rect	223	75	224	76
rect	223	77	224	78
rect	223	78	224	79
rect	223	80	224	81
rect	223	81	224	82
rect	223	83	224	84
rect	223	84	224	85
rect	223	86	224	87
rect	223	87	224	88
rect	223	89	224	90
rect	223	90	224	91
rect	223	92	224	93
rect	223	93	224	94
rect	223	95	224	96
rect	223	96	224	97
rect	223	98	224	99
rect	223	99	224	100
rect	223	101	224	102
rect	223	102	224	103
rect	223	104	224	105
rect	223	105	224	106
rect	223	107	224	108
rect	223	108	224	109
rect	223	110	224	111
rect	223	111	224	112
rect	223	113	224	114
rect	223	114	224	115
rect	223	116	224	117
rect	223	117	224	118
rect	223	119	224	120
rect	223	120	224	121
rect	223	122	224	123
rect	223	123	224	124
rect	223	125	224	126
rect	223	126	224	127
rect	223	128	224	129
rect	223	129	224	130
rect	223	131	224	132
rect	223	132	224	133
rect	223	134	224	135
rect	223	135	224	136
rect	223	137	224	138
rect	223	138	224	139
rect	223	140	224	141
rect	223	141	224	142
rect	223	143	224	144
rect	223	144	224	145
rect	223	146	224	147
rect	223	147	224	148
rect	223	149	224	150
rect	223	150	224	151
rect	223	152	224	153
rect	223	153	224	154
rect	223	155	224	156
rect	223	156	224	157
rect	223	158	224	159
rect	223	159	224	160
rect	223	161	224	162
rect	223	162	224	163
rect	223	164	224	165
rect	223	165	224	166
rect	223	167	224	168
rect	223	168	224	169
rect	223	170	224	171
rect	223	171	224	172
rect	223	173	224	174
rect	223	174	224	175
rect	223	176	224	177
rect	223	177	224	178
rect	223	179	224	180
rect	223	180	224	181
rect	223	182	224	183
rect	223	183	224	184
rect	223	185	224	186
rect	223	186	224	187
rect	223	188	224	189
rect	223	189	224	190
rect	223	191	224	192
rect	223	192	224	193
rect	223	194	224	195
rect	223	195	224	196
rect	223	197	224	198
rect	223	198	224	199
rect	223	200	224	201
rect	223	201	224	202
rect	223	203	224	204
rect	223	204	224	205
rect	223	206	224	207
rect	223	207	224	208
rect	223	209	224	210
rect	223	210	224	211
rect	223	212	224	213
rect	223	213	224	214
rect	223	215	224	216
rect	223	216	224	217
rect	223	218	224	219
rect	223	219	224	220
rect	223	221	224	222
rect	223	222	224	223
rect	223	224	224	225
rect	223	225	224	226
rect	223	227	224	228
rect	223	228	224	229
rect	223	230	224	231
rect	223	231	224	232
rect	223	233	224	234
rect	223	234	224	235
rect	223	236	224	237
rect	223	237	224	238
rect	223	239	224	240
rect	223	240	224	241
rect	223	242	224	243
rect	223	243	224	244
rect	223	245	224	246
rect	223	246	224	247
rect	223	248	224	249
rect	223	249	224	250
rect	223	251	224	252
rect	223	252	224	253
rect	223	253	224	254
rect	223	254	224	255
rect	223	255	224	256
rect	223	257	224	258
rect	223	258	224	259
rect	223	260	224	261
rect	223	261	224	262
rect	223	262	224	263
rect	223	263	224	264
rect	223	264	224	265
rect	223	266	224	267
rect	223	267	224	268
rect	223	268	224	269
rect	223	269	224	270
rect	223	270	224	271
rect	223	271	224	272
rect	223	272	224	273
rect	223	273	224	274
rect	223	275	224	276
rect	223	276	224	277
rect	223	278	224	279
rect	223	279	224	280
rect	223	280	224	281
rect	223	281	224	282
rect	223	282	224	283
rect	223	283	224	284
rect	223	284	224	285
rect	223	285	224	286
rect	223	286	224	287
rect	223	287	224	288
rect	224	0	225	1
rect	224	1	225	2
rect	224	2	225	3
rect	224	3	225	4
rect	224	4	225	5
rect	224	5	225	6
rect	224	6	225	7
rect	224	8	225	9
rect	224	9	225	10
rect	224	11	225	12
rect	224	12	225	13
rect	224	14	225	15
rect	224	15	225	16
rect	224	17	225	18
rect	224	18	225	19
rect	224	20	225	21
rect	224	21	225	22
rect	224	23	225	24
rect	224	24	225	25
rect	224	26	225	27
rect	224	27	225	28
rect	224	29	225	30
rect	224	30	225	31
rect	224	32	225	33
rect	224	33	225	34
rect	224	35	225	36
rect	224	36	225	37
rect	224	38	225	39
rect	224	39	225	40
rect	224	41	225	42
rect	224	42	225	43
rect	224	44	225	45
rect	224	45	225	46
rect	224	47	225	48
rect	224	48	225	49
rect	224	50	225	51
rect	224	51	225	52
rect	224	53	225	54
rect	224	54	225	55
rect	224	56	225	57
rect	224	57	225	58
rect	224	59	225	60
rect	224	60	225	61
rect	224	62	225	63
rect	224	63	225	64
rect	224	65	225	66
rect	224	66	225	67
rect	224	68	225	69
rect	224	69	225	70
rect	224	71	225	72
rect	224	72	225	73
rect	224	74	225	75
rect	224	75	225	76
rect	224	77	225	78
rect	224	78	225	79
rect	224	80	225	81
rect	224	81	225	82
rect	224	83	225	84
rect	224	84	225	85
rect	224	86	225	87
rect	224	87	225	88
rect	224	89	225	90
rect	224	90	225	91
rect	224	92	225	93
rect	224	93	225	94
rect	224	95	225	96
rect	224	96	225	97
rect	224	98	225	99
rect	224	99	225	100
rect	224	101	225	102
rect	224	102	225	103
rect	224	104	225	105
rect	224	105	225	106
rect	224	107	225	108
rect	224	108	225	109
rect	224	110	225	111
rect	224	111	225	112
rect	224	113	225	114
rect	224	114	225	115
rect	224	116	225	117
rect	224	117	225	118
rect	224	119	225	120
rect	224	120	225	121
rect	224	122	225	123
rect	224	123	225	124
rect	224	125	225	126
rect	224	126	225	127
rect	224	128	225	129
rect	224	129	225	130
rect	224	131	225	132
rect	224	132	225	133
rect	224	134	225	135
rect	224	135	225	136
rect	224	137	225	138
rect	224	138	225	139
rect	224	140	225	141
rect	224	141	225	142
rect	224	143	225	144
rect	224	144	225	145
rect	224	146	225	147
rect	224	147	225	148
rect	224	149	225	150
rect	224	150	225	151
rect	224	152	225	153
rect	224	153	225	154
rect	224	155	225	156
rect	224	156	225	157
rect	224	158	225	159
rect	224	159	225	160
rect	224	161	225	162
rect	224	162	225	163
rect	224	164	225	165
rect	224	165	225	166
rect	224	167	225	168
rect	224	168	225	169
rect	224	170	225	171
rect	224	171	225	172
rect	224	173	225	174
rect	224	174	225	175
rect	224	176	225	177
rect	224	177	225	178
rect	224	179	225	180
rect	224	180	225	181
rect	224	182	225	183
rect	224	183	225	184
rect	224	185	225	186
rect	224	186	225	187
rect	224	188	225	189
rect	224	189	225	190
rect	224	191	225	192
rect	224	192	225	193
rect	224	194	225	195
rect	224	195	225	196
rect	224	197	225	198
rect	224	198	225	199
rect	224	200	225	201
rect	224	201	225	202
rect	224	203	225	204
rect	224	204	225	205
rect	224	206	225	207
rect	224	207	225	208
rect	224	209	225	210
rect	224	210	225	211
rect	224	212	225	213
rect	224	213	225	214
rect	224	215	225	216
rect	224	216	225	217
rect	224	218	225	219
rect	224	219	225	220
rect	224	221	225	222
rect	224	222	225	223
rect	224	224	225	225
rect	224	225	225	226
rect	224	227	225	228
rect	224	228	225	229
rect	224	230	225	231
rect	224	231	225	232
rect	224	233	225	234
rect	224	234	225	235
rect	224	236	225	237
rect	224	237	225	238
rect	224	239	225	240
rect	224	240	225	241
rect	224	242	225	243
rect	224	243	225	244
rect	224	245	225	246
rect	224	246	225	247
rect	224	248	225	249
rect	224	249	225	250
rect	224	251	225	252
rect	224	252	225	253
rect	224	253	225	254
rect	224	254	225	255
rect	224	255	225	256
rect	224	257	225	258
rect	224	258	225	259
rect	224	260	225	261
rect	224	261	225	262
rect	224	262	225	263
rect	224	263	225	264
rect	224	264	225	265
rect	224	266	225	267
rect	224	267	225	268
rect	224	268	225	269
rect	224	269	225	270
rect	224	270	225	271
rect	224	271	225	272
rect	224	272	225	273
rect	224	273	225	274
rect	224	275	225	276
rect	224	276	225	277
rect	224	278	225	279
rect	224	279	225	280
rect	224	280	225	281
rect	224	281	225	282
rect	224	282	225	283
rect	224	283	225	284
rect	224	284	225	285
rect	224	285	225	286
rect	224	286	225	287
rect	224	287	225	288
rect	225	0	226	1
rect	225	1	226	2
rect	225	2	226	3
rect	225	3	226	4
rect	225	4	226	5
rect	225	5	226	6
rect	225	6	226	7
rect	225	8	226	9
rect	225	9	226	10
rect	225	11	226	12
rect	225	12	226	13
rect	225	14	226	15
rect	225	15	226	16
rect	225	17	226	18
rect	225	18	226	19
rect	225	20	226	21
rect	225	21	226	22
rect	225	23	226	24
rect	225	24	226	25
rect	225	26	226	27
rect	225	27	226	28
rect	225	29	226	30
rect	225	30	226	31
rect	225	32	226	33
rect	225	33	226	34
rect	225	35	226	36
rect	225	36	226	37
rect	225	38	226	39
rect	225	39	226	40
rect	225	41	226	42
rect	225	42	226	43
rect	225	44	226	45
rect	225	45	226	46
rect	225	47	226	48
rect	225	48	226	49
rect	225	50	226	51
rect	225	51	226	52
rect	225	53	226	54
rect	225	54	226	55
rect	225	56	226	57
rect	225	57	226	58
rect	225	59	226	60
rect	225	60	226	61
rect	225	62	226	63
rect	225	63	226	64
rect	225	65	226	66
rect	225	66	226	67
rect	225	68	226	69
rect	225	69	226	70
rect	225	71	226	72
rect	225	72	226	73
rect	225	74	226	75
rect	225	75	226	76
rect	225	77	226	78
rect	225	78	226	79
rect	225	80	226	81
rect	225	81	226	82
rect	225	83	226	84
rect	225	84	226	85
rect	225	86	226	87
rect	225	87	226	88
rect	225	89	226	90
rect	225	90	226	91
rect	225	92	226	93
rect	225	93	226	94
rect	225	95	226	96
rect	225	96	226	97
rect	225	98	226	99
rect	225	99	226	100
rect	225	101	226	102
rect	225	102	226	103
rect	225	104	226	105
rect	225	105	226	106
rect	225	107	226	108
rect	225	108	226	109
rect	225	110	226	111
rect	225	111	226	112
rect	225	113	226	114
rect	225	114	226	115
rect	225	116	226	117
rect	225	117	226	118
rect	225	119	226	120
rect	225	120	226	121
rect	225	122	226	123
rect	225	123	226	124
rect	225	125	226	126
rect	225	126	226	127
rect	225	128	226	129
rect	225	129	226	130
rect	225	131	226	132
rect	225	132	226	133
rect	225	134	226	135
rect	225	135	226	136
rect	225	137	226	138
rect	225	138	226	139
rect	225	140	226	141
rect	225	141	226	142
rect	225	143	226	144
rect	225	144	226	145
rect	225	146	226	147
rect	225	147	226	148
rect	225	149	226	150
rect	225	150	226	151
rect	225	152	226	153
rect	225	153	226	154
rect	225	155	226	156
rect	225	156	226	157
rect	225	158	226	159
rect	225	159	226	160
rect	225	161	226	162
rect	225	162	226	163
rect	225	164	226	165
rect	225	165	226	166
rect	225	167	226	168
rect	225	168	226	169
rect	225	170	226	171
rect	225	171	226	172
rect	225	173	226	174
rect	225	174	226	175
rect	225	176	226	177
rect	225	177	226	178
rect	225	179	226	180
rect	225	180	226	181
rect	225	182	226	183
rect	225	183	226	184
rect	225	185	226	186
rect	225	186	226	187
rect	225	188	226	189
rect	225	189	226	190
rect	225	191	226	192
rect	225	192	226	193
rect	225	194	226	195
rect	225	195	226	196
rect	225	197	226	198
rect	225	198	226	199
rect	225	200	226	201
rect	225	201	226	202
rect	225	203	226	204
rect	225	204	226	205
rect	225	206	226	207
rect	225	207	226	208
rect	225	209	226	210
rect	225	210	226	211
rect	225	212	226	213
rect	225	213	226	214
rect	225	215	226	216
rect	225	216	226	217
rect	225	218	226	219
rect	225	219	226	220
rect	225	221	226	222
rect	225	222	226	223
rect	225	224	226	225
rect	225	225	226	226
rect	225	227	226	228
rect	225	228	226	229
rect	225	230	226	231
rect	225	231	226	232
rect	225	233	226	234
rect	225	234	226	235
rect	225	236	226	237
rect	225	237	226	238
rect	225	239	226	240
rect	225	240	226	241
rect	225	242	226	243
rect	225	243	226	244
rect	225	245	226	246
rect	225	246	226	247
rect	225	248	226	249
rect	225	249	226	250
rect	225	251	226	252
rect	225	252	226	253
rect	225	253	226	254
rect	225	254	226	255
rect	225	255	226	256
rect	225	257	226	258
rect	225	258	226	259
rect	225	260	226	261
rect	225	261	226	262
rect	225	262	226	263
rect	225	263	226	264
rect	225	264	226	265
rect	225	266	226	267
rect	225	267	226	268
rect	225	268	226	269
rect	225	269	226	270
rect	225	270	226	271
rect	225	271	226	272
rect	225	272	226	273
rect	225	273	226	274
rect	225	275	226	276
rect	225	276	226	277
rect	225	278	226	279
rect	225	279	226	280
rect	225	280	226	281
rect	225	281	226	282
rect	225	282	226	283
rect	225	283	226	284
rect	225	284	226	285
rect	225	285	226	286
rect	225	286	226	287
rect	225	287	226	288
rect	226	0	227	1
rect	226	1	227	2
rect	226	2	227	3
rect	226	3	227	4
rect	226	4	227	5
rect	226	5	227	6
rect	226	6	227	7
rect	226	8	227	9
rect	226	9	227	10
rect	226	11	227	12
rect	226	12	227	13
rect	226	14	227	15
rect	226	15	227	16
rect	226	17	227	18
rect	226	18	227	19
rect	226	20	227	21
rect	226	21	227	22
rect	226	23	227	24
rect	226	24	227	25
rect	226	26	227	27
rect	226	27	227	28
rect	226	29	227	30
rect	226	30	227	31
rect	226	32	227	33
rect	226	33	227	34
rect	226	35	227	36
rect	226	36	227	37
rect	226	38	227	39
rect	226	39	227	40
rect	226	41	227	42
rect	226	42	227	43
rect	226	44	227	45
rect	226	45	227	46
rect	226	47	227	48
rect	226	48	227	49
rect	226	50	227	51
rect	226	51	227	52
rect	226	53	227	54
rect	226	54	227	55
rect	226	56	227	57
rect	226	57	227	58
rect	226	59	227	60
rect	226	60	227	61
rect	226	62	227	63
rect	226	63	227	64
rect	226	65	227	66
rect	226	66	227	67
rect	226	68	227	69
rect	226	69	227	70
rect	226	71	227	72
rect	226	72	227	73
rect	226	74	227	75
rect	226	75	227	76
rect	226	77	227	78
rect	226	78	227	79
rect	226	80	227	81
rect	226	81	227	82
rect	226	83	227	84
rect	226	84	227	85
rect	226	86	227	87
rect	226	87	227	88
rect	226	89	227	90
rect	226	90	227	91
rect	226	92	227	93
rect	226	93	227	94
rect	226	95	227	96
rect	226	96	227	97
rect	226	98	227	99
rect	226	99	227	100
rect	226	101	227	102
rect	226	102	227	103
rect	226	104	227	105
rect	226	105	227	106
rect	226	107	227	108
rect	226	108	227	109
rect	226	110	227	111
rect	226	111	227	112
rect	226	113	227	114
rect	226	114	227	115
rect	226	116	227	117
rect	226	117	227	118
rect	226	119	227	120
rect	226	120	227	121
rect	226	122	227	123
rect	226	123	227	124
rect	226	125	227	126
rect	226	126	227	127
rect	226	128	227	129
rect	226	129	227	130
rect	226	131	227	132
rect	226	132	227	133
rect	226	134	227	135
rect	226	135	227	136
rect	226	137	227	138
rect	226	138	227	139
rect	226	140	227	141
rect	226	141	227	142
rect	226	143	227	144
rect	226	144	227	145
rect	226	146	227	147
rect	226	147	227	148
rect	226	149	227	150
rect	226	150	227	151
rect	226	152	227	153
rect	226	153	227	154
rect	226	155	227	156
rect	226	156	227	157
rect	226	158	227	159
rect	226	159	227	160
rect	226	161	227	162
rect	226	162	227	163
rect	226	164	227	165
rect	226	165	227	166
rect	226	167	227	168
rect	226	168	227	169
rect	226	170	227	171
rect	226	171	227	172
rect	226	173	227	174
rect	226	174	227	175
rect	226	176	227	177
rect	226	177	227	178
rect	226	179	227	180
rect	226	180	227	181
rect	226	182	227	183
rect	226	183	227	184
rect	226	185	227	186
rect	226	186	227	187
rect	226	188	227	189
rect	226	189	227	190
rect	226	191	227	192
rect	226	192	227	193
rect	226	194	227	195
rect	226	195	227	196
rect	226	197	227	198
rect	226	198	227	199
rect	226	200	227	201
rect	226	201	227	202
rect	226	203	227	204
rect	226	204	227	205
rect	226	206	227	207
rect	226	207	227	208
rect	226	209	227	210
rect	226	210	227	211
rect	226	212	227	213
rect	226	213	227	214
rect	226	215	227	216
rect	226	216	227	217
rect	226	218	227	219
rect	226	219	227	220
rect	226	221	227	222
rect	226	222	227	223
rect	226	224	227	225
rect	226	225	227	226
rect	226	227	227	228
rect	226	228	227	229
rect	226	230	227	231
rect	226	231	227	232
rect	226	233	227	234
rect	226	234	227	235
rect	226	236	227	237
rect	226	237	227	238
rect	226	239	227	240
rect	226	240	227	241
rect	226	242	227	243
rect	226	243	227	244
rect	226	245	227	246
rect	226	246	227	247
rect	226	248	227	249
rect	226	249	227	250
rect	226	251	227	252
rect	226	252	227	253
rect	226	253	227	254
rect	226	254	227	255
rect	226	255	227	256
rect	226	257	227	258
rect	226	258	227	259
rect	226	260	227	261
rect	226	261	227	262
rect	226	262	227	263
rect	226	263	227	264
rect	226	264	227	265
rect	226	266	227	267
rect	226	267	227	268
rect	226	268	227	269
rect	226	269	227	270
rect	226	270	227	271
rect	226	271	227	272
rect	226	272	227	273
rect	226	273	227	274
rect	226	275	227	276
rect	226	276	227	277
rect	226	278	227	279
rect	226	279	227	280
rect	226	280	227	281
rect	226	281	227	282
rect	226	282	227	283
rect	226	283	227	284
rect	226	284	227	285
rect	226	285	227	286
rect	226	286	227	287
rect	226	287	227	288
rect	235	0	236	1
rect	235	1	236	2
rect	235	2	236	3
rect	235	3	236	4
rect	235	4	236	5
rect	235	5	236	6
rect	235	6	236	7
rect	235	8	236	9
rect	235	9	236	10
rect	235	11	236	12
rect	235	12	236	13
rect	235	14	236	15
rect	235	15	236	16
rect	235	17	236	18
rect	235	18	236	19
rect	235	20	236	21
rect	235	21	236	22
rect	235	23	236	24
rect	235	24	236	25
rect	235	26	236	27
rect	235	27	236	28
rect	235	29	236	30
rect	235	30	236	31
rect	235	32	236	33
rect	235	33	236	34
rect	235	35	236	36
rect	235	36	236	37
rect	235	38	236	39
rect	235	39	236	40
rect	235	41	236	42
rect	235	42	236	43
rect	235	44	236	45
rect	235	45	236	46
rect	235	47	236	48
rect	235	48	236	49
rect	235	50	236	51
rect	235	51	236	52
rect	235	53	236	54
rect	235	54	236	55
rect	235	56	236	57
rect	235	57	236	58
rect	235	59	236	60
rect	235	60	236	61
rect	235	62	236	63
rect	235	63	236	64
rect	235	65	236	66
rect	235	66	236	67
rect	235	68	236	69
rect	235	69	236	70
rect	235	71	236	72
rect	235	72	236	73
rect	235	74	236	75
rect	235	75	236	76
rect	235	77	236	78
rect	235	78	236	79
rect	235	80	236	81
rect	235	81	236	82
rect	235	83	236	84
rect	235	84	236	85
rect	235	86	236	87
rect	235	87	236	88
rect	235	89	236	90
rect	235	90	236	91
rect	235	91	236	92
rect	235	92	236	93
rect	235	93	236	94
rect	235	95	236	96
rect	235	96	236	97
rect	235	98	236	99
rect	235	99	236	100
rect	235	101	236	102
rect	235	102	236	103
rect	235	104	236	105
rect	235	105	236	106
rect	235	107	236	108
rect	235	108	236	109
rect	235	110	236	111
rect	235	111	236	112
rect	235	113	236	114
rect	235	114	236	115
rect	235	116	236	117
rect	235	117	236	118
rect	235	119	236	120
rect	235	120	236	121
rect	235	122	236	123
rect	235	123	236	124
rect	235	125	236	126
rect	235	126	236	127
rect	235	128	236	129
rect	235	129	236	130
rect	235	130	236	131
rect	235	131	236	132
rect	235	132	236	133
rect	235	134	236	135
rect	235	135	236	136
rect	235	137	236	138
rect	235	138	236	139
rect	235	140	236	141
rect	235	141	236	142
rect	235	143	236	144
rect	235	144	236	145
rect	235	146	236	147
rect	235	147	236	148
rect	235	149	236	150
rect	235	150	236	151
rect	235	152	236	153
rect	235	153	236	154
rect	235	155	236	156
rect	235	156	236	157
rect	235	158	236	159
rect	235	159	236	160
rect	235	161	236	162
rect	235	162	236	163
rect	235	164	236	165
rect	235	165	236	166
rect	235	167	236	168
rect	235	168	236	169
rect	235	170	236	171
rect	235	171	236	172
rect	235	173	236	174
rect	235	174	236	175
rect	235	176	236	177
rect	235	177	236	178
rect	235	179	236	180
rect	235	180	236	181
rect	235	182	236	183
rect	235	183	236	184
rect	235	185	236	186
rect	235	186	236	187
rect	235	188	236	189
rect	235	189	236	190
rect	235	190	236	191
rect	235	191	236	192
rect	235	192	236	193
rect	235	194	236	195
rect	235	195	236	196
rect	235	197	236	198
rect	235	198	236	199
rect	235	200	236	201
rect	235	201	236	202
rect	235	203	236	204
rect	235	204	236	205
rect	235	206	236	207
rect	235	207	236	208
rect	235	209	236	210
rect	235	210	236	211
rect	235	212	236	213
rect	235	213	236	214
rect	235	215	236	216
rect	235	216	236	217
rect	235	218	236	219
rect	235	219	236	220
rect	235	221	236	222
rect	235	222	236	223
rect	235	224	236	225
rect	235	225	236	226
rect	235	227	236	228
rect	235	228	236	229
rect	235	230	236	231
rect	235	231	236	232
rect	235	233	236	234
rect	235	234	236	235
rect	235	236	236	237
rect	235	237	236	238
rect	235	239	236	240
rect	235	240	236	241
rect	235	242	236	243
rect	235	243	236	244
rect	235	245	236	246
rect	235	246	236	247
rect	235	248	236	249
rect	235	249	236	250
rect	235	251	236	252
rect	235	252	236	253
rect	235	253	236	254
rect	235	254	236	255
rect	235	255	236	256
rect	235	257	236	258
rect	235	258	236	259
rect	235	260	236	261
rect	235	261	236	262
rect	235	262	236	263
rect	235	263	236	264
rect	235	264	236	265
rect	235	265	236	266
rect	235	266	236	267
rect	235	267	236	268
rect	235	268	236	269
rect	235	269	236	270
rect	235	270	236	271
rect	235	271	236	272
rect	235	272	236	273
rect	235	273	236	274
rect	235	274	236	275
rect	235	275	236	276
rect	235	276	236	277
rect	235	277	236	278
rect	235	278	236	279
rect	235	279	236	280
rect	235	280	236	281
rect	235	281	236	282
rect	235	282	236	283
rect	235	283	236	284
rect	235	284	236	285
rect	235	285	236	286
rect	235	286	236	287
rect	235	287	236	288
rect	237	0	238	1
rect	237	1	238	2
rect	237	2	238	3
rect	237	3	238	4
rect	237	4	238	5
rect	237	5	238	6
rect	237	6	238	7
rect	237	8	238	9
rect	237	9	238	10
rect	237	11	238	12
rect	237	12	238	13
rect	237	14	238	15
rect	237	15	238	16
rect	237	17	238	18
rect	237	18	238	19
rect	237	20	238	21
rect	237	21	238	22
rect	237	23	238	24
rect	237	24	238	25
rect	237	26	238	27
rect	237	27	238	28
rect	237	29	238	30
rect	237	30	238	31
rect	237	32	238	33
rect	237	33	238	34
rect	237	35	238	36
rect	237	36	238	37
rect	237	38	238	39
rect	237	39	238	40
rect	237	41	238	42
rect	237	42	238	43
rect	237	44	238	45
rect	237	45	238	46
rect	237	47	238	48
rect	237	48	238	49
rect	237	50	238	51
rect	237	51	238	52
rect	237	53	238	54
rect	237	54	238	55
rect	237	56	238	57
rect	237	57	238	58
rect	237	59	238	60
rect	237	60	238	61
rect	237	62	238	63
rect	237	63	238	64
rect	237	65	238	66
rect	237	66	238	67
rect	237	68	238	69
rect	237	69	238	70
rect	237	71	238	72
rect	237	72	238	73
rect	237	74	238	75
rect	237	75	238	76
rect	237	77	238	78
rect	237	78	238	79
rect	237	80	238	81
rect	237	81	238	82
rect	237	83	238	84
rect	237	84	238	85
rect	237	86	238	87
rect	237	87	238	88
rect	237	89	238	90
rect	237	90	238	91
rect	237	91	238	92
rect	237	92	238	93
rect	237	93	238	94
rect	237	95	238	96
rect	237	96	238	97
rect	237	98	238	99
rect	237	99	238	100
rect	237	101	238	102
rect	237	102	238	103
rect	237	104	238	105
rect	237	105	238	106
rect	237	107	238	108
rect	237	108	238	109
rect	237	110	238	111
rect	237	111	238	112
rect	237	113	238	114
rect	237	114	238	115
rect	237	116	238	117
rect	237	117	238	118
rect	237	119	238	120
rect	237	120	238	121
rect	237	122	238	123
rect	237	123	238	124
rect	237	125	238	126
rect	237	126	238	127
rect	237	128	238	129
rect	237	129	238	130
rect	237	130	238	131
rect	237	131	238	132
rect	237	132	238	133
rect	237	134	238	135
rect	237	135	238	136
rect	237	137	238	138
rect	237	138	238	139
rect	237	140	238	141
rect	237	141	238	142
rect	237	143	238	144
rect	237	144	238	145
rect	237	146	238	147
rect	237	147	238	148
rect	237	149	238	150
rect	237	150	238	151
rect	237	152	238	153
rect	237	153	238	154
rect	237	155	238	156
rect	237	156	238	157
rect	237	158	238	159
rect	237	159	238	160
rect	237	161	238	162
rect	237	162	238	163
rect	237	164	238	165
rect	237	165	238	166
rect	237	167	238	168
rect	237	168	238	169
rect	237	170	238	171
rect	237	171	238	172
rect	237	173	238	174
rect	237	174	238	175
rect	237	176	238	177
rect	237	177	238	178
rect	237	179	238	180
rect	237	180	238	181
rect	237	182	238	183
rect	237	183	238	184
rect	237	185	238	186
rect	237	186	238	187
rect	237	188	238	189
rect	237	189	238	190
rect	237	190	238	191
rect	237	191	238	192
rect	237	192	238	193
rect	237	194	238	195
rect	237	195	238	196
rect	237	197	238	198
rect	237	198	238	199
rect	237	200	238	201
rect	237	201	238	202
rect	237	203	238	204
rect	237	204	238	205
rect	237	206	238	207
rect	237	207	238	208
rect	237	209	238	210
rect	237	210	238	211
rect	237	212	238	213
rect	237	213	238	214
rect	237	215	238	216
rect	237	216	238	217
rect	237	218	238	219
rect	237	219	238	220
rect	237	221	238	222
rect	237	222	238	223
rect	237	224	238	225
rect	237	225	238	226
rect	237	227	238	228
rect	237	228	238	229
rect	237	230	238	231
rect	237	231	238	232
rect	237	233	238	234
rect	237	234	238	235
rect	237	236	238	237
rect	237	237	238	238
rect	237	239	238	240
rect	237	240	238	241
rect	237	242	238	243
rect	237	243	238	244
rect	237	245	238	246
rect	237	246	238	247
rect	237	248	238	249
rect	237	249	238	250
rect	237	251	238	252
rect	237	252	238	253
rect	237	253	238	254
rect	237	254	238	255
rect	237	255	238	256
rect	237	257	238	258
rect	237	258	238	259
rect	237	260	238	261
rect	237	261	238	262
rect	237	262	238	263
rect	237	263	238	264
rect	237	264	238	265
rect	237	265	238	266
rect	237	266	238	267
rect	237	267	238	268
rect	237	268	238	269
rect	237	269	238	270
rect	237	270	238	271
rect	237	271	238	272
rect	237	272	238	273
rect	237	273	238	274
rect	237	274	238	275
rect	237	275	238	276
rect	237	276	238	277
rect	237	277	238	278
rect	237	278	238	279
rect	237	279	238	280
rect	237	280	238	281
rect	237	281	238	282
rect	237	282	238	283
rect	237	283	238	284
rect	237	284	238	285
rect	238	0	239	1
rect	238	1	239	2
rect	238	2	239	3
rect	238	3	239	4
rect	238	4	239	5
rect	238	5	239	6
rect	238	6	239	7
rect	238	8	239	9
rect	238	9	239	10
rect	238	11	239	12
rect	238	12	239	13
rect	238	14	239	15
rect	238	15	239	16
rect	238	17	239	18
rect	238	18	239	19
rect	238	20	239	21
rect	238	21	239	22
rect	238	23	239	24
rect	238	24	239	25
rect	238	26	239	27
rect	238	27	239	28
rect	238	29	239	30
rect	238	30	239	31
rect	238	32	239	33
rect	238	33	239	34
rect	238	35	239	36
rect	238	36	239	37
rect	238	38	239	39
rect	238	39	239	40
rect	238	41	239	42
rect	238	42	239	43
rect	238	44	239	45
rect	238	45	239	46
rect	238	47	239	48
rect	238	48	239	49
rect	238	50	239	51
rect	238	51	239	52
rect	238	53	239	54
rect	238	54	239	55
rect	238	56	239	57
rect	238	57	239	58
rect	238	59	239	60
rect	238	60	239	61
rect	238	62	239	63
rect	238	63	239	64
rect	238	65	239	66
rect	238	66	239	67
rect	238	68	239	69
rect	238	69	239	70
rect	238	71	239	72
rect	238	72	239	73
rect	238	74	239	75
rect	238	75	239	76
rect	238	77	239	78
rect	238	78	239	79
rect	238	80	239	81
rect	238	81	239	82
rect	238	83	239	84
rect	238	84	239	85
rect	238	86	239	87
rect	238	87	239	88
rect	238	89	239	90
rect	238	90	239	91
rect	238	91	239	92
rect	238	92	239	93
rect	238	93	239	94
rect	238	95	239	96
rect	238	96	239	97
rect	238	98	239	99
rect	238	99	239	100
rect	238	101	239	102
rect	238	102	239	103
rect	238	104	239	105
rect	238	105	239	106
rect	238	107	239	108
rect	238	108	239	109
rect	238	110	239	111
rect	238	111	239	112
rect	238	113	239	114
rect	238	114	239	115
rect	238	116	239	117
rect	238	117	239	118
rect	238	119	239	120
rect	238	120	239	121
rect	238	122	239	123
rect	238	123	239	124
rect	238	125	239	126
rect	238	126	239	127
rect	238	128	239	129
rect	238	129	239	130
rect	238	130	239	131
rect	238	131	239	132
rect	238	132	239	133
rect	238	134	239	135
rect	238	135	239	136
rect	238	137	239	138
rect	238	138	239	139
rect	238	140	239	141
rect	238	141	239	142
rect	238	143	239	144
rect	238	144	239	145
rect	238	146	239	147
rect	238	147	239	148
rect	238	149	239	150
rect	238	150	239	151
rect	238	152	239	153
rect	238	153	239	154
rect	238	155	239	156
rect	238	156	239	157
rect	238	158	239	159
rect	238	159	239	160
rect	238	161	239	162
rect	238	162	239	163
rect	238	164	239	165
rect	238	165	239	166
rect	238	167	239	168
rect	238	168	239	169
rect	238	170	239	171
rect	238	171	239	172
rect	238	173	239	174
rect	238	174	239	175
rect	238	176	239	177
rect	238	177	239	178
rect	238	179	239	180
rect	238	180	239	181
rect	238	182	239	183
rect	238	183	239	184
rect	238	185	239	186
rect	238	186	239	187
rect	238	188	239	189
rect	238	189	239	190
rect	238	190	239	191
rect	238	191	239	192
rect	238	192	239	193
rect	238	194	239	195
rect	238	195	239	196
rect	238	197	239	198
rect	238	198	239	199
rect	238	200	239	201
rect	238	201	239	202
rect	238	203	239	204
rect	238	204	239	205
rect	238	206	239	207
rect	238	207	239	208
rect	238	209	239	210
rect	238	210	239	211
rect	238	212	239	213
rect	238	213	239	214
rect	238	215	239	216
rect	238	216	239	217
rect	238	218	239	219
rect	238	219	239	220
rect	238	221	239	222
rect	238	222	239	223
rect	238	224	239	225
rect	238	225	239	226
rect	238	227	239	228
rect	238	228	239	229
rect	238	230	239	231
rect	238	231	239	232
rect	238	233	239	234
rect	238	234	239	235
rect	238	236	239	237
rect	238	237	239	238
rect	238	239	239	240
rect	238	240	239	241
rect	238	242	239	243
rect	238	243	239	244
rect	238	245	239	246
rect	238	246	239	247
rect	238	248	239	249
rect	238	249	239	250
rect	238	251	239	252
rect	238	252	239	253
rect	238	253	239	254
rect	238	254	239	255
rect	238	255	239	256
rect	238	257	239	258
rect	238	258	239	259
rect	238	260	239	261
rect	238	261	239	262
rect	238	262	239	263
rect	238	263	239	264
rect	238	264	239	265
rect	238	265	239	266
rect	238	266	239	267
rect	238	267	239	268
rect	238	268	239	269
rect	238	269	239	270
rect	238	270	239	271
rect	238	271	239	272
rect	238	272	239	273
rect	238	273	239	274
rect	238	274	239	275
rect	238	275	239	276
rect	238	276	239	277
rect	238	277	239	278
rect	238	278	239	279
rect	238	279	239	280
rect	238	280	239	281
rect	238	281	239	282
rect	238	282	239	283
rect	238	283	239	284
rect	238	284	239	285
rect	239	0	240	1
rect	239	1	240	2
rect	239	2	240	3
rect	239	3	240	4
rect	239	4	240	5
rect	239	5	240	6
rect	239	6	240	7
rect	239	8	240	9
rect	239	9	240	10
rect	239	11	240	12
rect	239	12	240	13
rect	239	14	240	15
rect	239	15	240	16
rect	239	17	240	18
rect	239	18	240	19
rect	239	20	240	21
rect	239	21	240	22
rect	239	23	240	24
rect	239	24	240	25
rect	239	26	240	27
rect	239	27	240	28
rect	239	29	240	30
rect	239	30	240	31
rect	239	32	240	33
rect	239	33	240	34
rect	239	35	240	36
rect	239	36	240	37
rect	239	38	240	39
rect	239	39	240	40
rect	239	41	240	42
rect	239	42	240	43
rect	239	44	240	45
rect	239	45	240	46
rect	239	47	240	48
rect	239	48	240	49
rect	239	50	240	51
rect	239	51	240	52
rect	239	53	240	54
rect	239	54	240	55
rect	239	56	240	57
rect	239	57	240	58
rect	239	59	240	60
rect	239	60	240	61
rect	239	62	240	63
rect	239	63	240	64
rect	239	65	240	66
rect	239	66	240	67
rect	239	68	240	69
rect	239	69	240	70
rect	239	71	240	72
rect	239	72	240	73
rect	239	74	240	75
rect	239	75	240	76
rect	239	77	240	78
rect	239	78	240	79
rect	239	80	240	81
rect	239	81	240	82
rect	239	83	240	84
rect	239	84	240	85
rect	239	86	240	87
rect	239	87	240	88
rect	239	89	240	90
rect	239	90	240	91
rect	239	91	240	92
rect	239	92	240	93
rect	239	93	240	94
rect	239	95	240	96
rect	239	96	240	97
rect	239	98	240	99
rect	239	99	240	100
rect	239	101	240	102
rect	239	102	240	103
rect	239	104	240	105
rect	239	105	240	106
rect	239	107	240	108
rect	239	108	240	109
rect	239	110	240	111
rect	239	111	240	112
rect	239	113	240	114
rect	239	114	240	115
rect	239	116	240	117
rect	239	117	240	118
rect	239	119	240	120
rect	239	120	240	121
rect	239	122	240	123
rect	239	123	240	124
rect	239	125	240	126
rect	239	126	240	127
rect	239	128	240	129
rect	239	129	240	130
rect	239	130	240	131
rect	239	131	240	132
rect	239	132	240	133
rect	239	134	240	135
rect	239	135	240	136
rect	239	137	240	138
rect	239	138	240	139
rect	239	140	240	141
rect	239	141	240	142
rect	239	143	240	144
rect	239	144	240	145
rect	239	146	240	147
rect	239	147	240	148
rect	239	149	240	150
rect	239	150	240	151
rect	239	152	240	153
rect	239	153	240	154
rect	239	155	240	156
rect	239	156	240	157
rect	239	158	240	159
rect	239	159	240	160
rect	239	161	240	162
rect	239	162	240	163
rect	239	164	240	165
rect	239	165	240	166
rect	239	167	240	168
rect	239	168	240	169
rect	239	170	240	171
rect	239	171	240	172
rect	239	173	240	174
rect	239	174	240	175
rect	239	176	240	177
rect	239	177	240	178
rect	239	179	240	180
rect	239	180	240	181
rect	239	182	240	183
rect	239	183	240	184
rect	239	185	240	186
rect	239	186	240	187
rect	239	188	240	189
rect	239	189	240	190
rect	239	190	240	191
rect	239	191	240	192
rect	239	192	240	193
rect	239	194	240	195
rect	239	195	240	196
rect	239	197	240	198
rect	239	198	240	199
rect	239	200	240	201
rect	239	201	240	202
rect	239	203	240	204
rect	239	204	240	205
rect	239	206	240	207
rect	239	207	240	208
rect	239	209	240	210
rect	239	210	240	211
rect	239	212	240	213
rect	239	213	240	214
rect	239	215	240	216
rect	239	216	240	217
rect	239	218	240	219
rect	239	219	240	220
rect	239	221	240	222
rect	239	222	240	223
rect	239	224	240	225
rect	239	225	240	226
rect	239	227	240	228
rect	239	228	240	229
rect	239	230	240	231
rect	239	231	240	232
rect	239	233	240	234
rect	239	234	240	235
rect	239	236	240	237
rect	239	237	240	238
rect	239	239	240	240
rect	239	240	240	241
rect	239	242	240	243
rect	239	243	240	244
rect	239	245	240	246
rect	239	246	240	247
rect	239	248	240	249
rect	239	249	240	250
rect	239	251	240	252
rect	239	252	240	253
rect	239	253	240	254
rect	239	254	240	255
rect	239	255	240	256
rect	239	257	240	258
rect	239	258	240	259
rect	239	260	240	261
rect	239	261	240	262
rect	239	262	240	263
rect	239	263	240	264
rect	239	264	240	265
rect	239	265	240	266
rect	239	266	240	267
rect	239	267	240	268
rect	239	268	240	269
rect	239	269	240	270
rect	239	270	240	271
rect	239	271	240	272
rect	239	272	240	273
rect	239	273	240	274
rect	239	274	240	275
rect	239	275	240	276
rect	239	276	240	277
rect	239	277	240	278
rect	239	278	240	279
rect	239	279	240	280
rect	239	280	240	281
rect	239	281	240	282
rect	239	282	240	283
rect	239	283	240	284
rect	239	284	240	285
rect	240	0	241	1
rect	240	1	241	2
rect	240	2	241	3
rect	240	3	241	4
rect	240	4	241	5
rect	240	5	241	6
rect	240	6	241	7
rect	240	8	241	9
rect	240	9	241	10
rect	240	11	241	12
rect	240	12	241	13
rect	240	14	241	15
rect	240	15	241	16
rect	240	17	241	18
rect	240	18	241	19
rect	240	20	241	21
rect	240	21	241	22
rect	240	23	241	24
rect	240	24	241	25
rect	240	26	241	27
rect	240	27	241	28
rect	240	29	241	30
rect	240	30	241	31
rect	240	32	241	33
rect	240	33	241	34
rect	240	35	241	36
rect	240	36	241	37
rect	240	38	241	39
rect	240	39	241	40
rect	240	41	241	42
rect	240	42	241	43
rect	240	44	241	45
rect	240	45	241	46
rect	240	47	241	48
rect	240	48	241	49
rect	240	50	241	51
rect	240	51	241	52
rect	240	53	241	54
rect	240	54	241	55
rect	240	56	241	57
rect	240	57	241	58
rect	240	59	241	60
rect	240	60	241	61
rect	240	62	241	63
rect	240	63	241	64
rect	240	65	241	66
rect	240	66	241	67
rect	240	68	241	69
rect	240	69	241	70
rect	240	71	241	72
rect	240	72	241	73
rect	240	74	241	75
rect	240	75	241	76
rect	240	77	241	78
rect	240	78	241	79
rect	240	80	241	81
rect	240	81	241	82
rect	240	83	241	84
rect	240	84	241	85
rect	240	86	241	87
rect	240	87	241	88
rect	240	89	241	90
rect	240	90	241	91
rect	240	91	241	92
rect	240	92	241	93
rect	240	93	241	94
rect	240	95	241	96
rect	240	96	241	97
rect	240	98	241	99
rect	240	99	241	100
rect	240	101	241	102
rect	240	102	241	103
rect	240	104	241	105
rect	240	105	241	106
rect	240	107	241	108
rect	240	108	241	109
rect	240	110	241	111
rect	240	111	241	112
rect	240	113	241	114
rect	240	114	241	115
rect	240	116	241	117
rect	240	117	241	118
rect	240	119	241	120
rect	240	120	241	121
rect	240	122	241	123
rect	240	123	241	124
rect	240	125	241	126
rect	240	126	241	127
rect	240	128	241	129
rect	240	129	241	130
rect	240	130	241	131
rect	240	131	241	132
rect	240	132	241	133
rect	240	134	241	135
rect	240	135	241	136
rect	240	137	241	138
rect	240	138	241	139
rect	240	140	241	141
rect	240	141	241	142
rect	240	143	241	144
rect	240	144	241	145
rect	240	146	241	147
rect	240	147	241	148
rect	240	149	241	150
rect	240	150	241	151
rect	240	152	241	153
rect	240	153	241	154
rect	240	155	241	156
rect	240	156	241	157
rect	240	158	241	159
rect	240	159	241	160
rect	240	161	241	162
rect	240	162	241	163
rect	240	164	241	165
rect	240	165	241	166
rect	240	167	241	168
rect	240	168	241	169
rect	240	170	241	171
rect	240	171	241	172
rect	240	173	241	174
rect	240	174	241	175
rect	240	176	241	177
rect	240	177	241	178
rect	240	179	241	180
rect	240	180	241	181
rect	240	182	241	183
rect	240	183	241	184
rect	240	185	241	186
rect	240	186	241	187
rect	240	188	241	189
rect	240	189	241	190
rect	240	190	241	191
rect	240	191	241	192
rect	240	192	241	193
rect	240	194	241	195
rect	240	195	241	196
rect	240	197	241	198
rect	240	198	241	199
rect	240	200	241	201
rect	240	201	241	202
rect	240	203	241	204
rect	240	204	241	205
rect	240	206	241	207
rect	240	207	241	208
rect	240	209	241	210
rect	240	210	241	211
rect	240	212	241	213
rect	240	213	241	214
rect	240	215	241	216
rect	240	216	241	217
rect	240	218	241	219
rect	240	219	241	220
rect	240	221	241	222
rect	240	222	241	223
rect	240	224	241	225
rect	240	225	241	226
rect	240	227	241	228
rect	240	228	241	229
rect	240	230	241	231
rect	240	231	241	232
rect	240	233	241	234
rect	240	234	241	235
rect	240	236	241	237
rect	240	237	241	238
rect	240	239	241	240
rect	240	240	241	241
rect	240	242	241	243
rect	240	243	241	244
rect	240	245	241	246
rect	240	246	241	247
rect	240	248	241	249
rect	240	249	241	250
rect	240	251	241	252
rect	240	252	241	253
rect	240	253	241	254
rect	240	254	241	255
rect	240	255	241	256
rect	240	257	241	258
rect	240	258	241	259
rect	240	260	241	261
rect	240	261	241	262
rect	240	262	241	263
rect	240	263	241	264
rect	240	264	241	265
rect	240	265	241	266
rect	240	266	241	267
rect	240	267	241	268
rect	240	268	241	269
rect	240	269	241	270
rect	240	270	241	271
rect	240	271	241	272
rect	240	272	241	273
rect	240	273	241	274
rect	240	274	241	275
rect	240	275	241	276
rect	240	276	241	277
rect	240	277	241	278
rect	240	278	241	279
rect	240	279	241	280
rect	240	280	241	281
rect	240	281	241	282
rect	240	282	241	283
rect	240	283	241	284
rect	240	284	241	285
rect	241	0	242	1
rect	241	1	242	2
rect	241	2	242	3
rect	241	3	242	4
rect	241	4	242	5
rect	241	5	242	6
rect	241	6	242	7
rect	241	8	242	9
rect	241	9	242	10
rect	241	11	242	12
rect	241	12	242	13
rect	241	14	242	15
rect	241	15	242	16
rect	241	17	242	18
rect	241	18	242	19
rect	241	20	242	21
rect	241	21	242	22
rect	241	23	242	24
rect	241	24	242	25
rect	241	26	242	27
rect	241	27	242	28
rect	241	29	242	30
rect	241	30	242	31
rect	241	32	242	33
rect	241	33	242	34
rect	241	35	242	36
rect	241	36	242	37
rect	241	38	242	39
rect	241	39	242	40
rect	241	41	242	42
rect	241	42	242	43
rect	241	44	242	45
rect	241	45	242	46
rect	241	47	242	48
rect	241	48	242	49
rect	241	50	242	51
rect	241	51	242	52
rect	241	53	242	54
rect	241	54	242	55
rect	241	56	242	57
rect	241	57	242	58
rect	241	59	242	60
rect	241	60	242	61
rect	241	62	242	63
rect	241	63	242	64
rect	241	65	242	66
rect	241	66	242	67
rect	241	68	242	69
rect	241	69	242	70
rect	241	71	242	72
rect	241	72	242	73
rect	241	74	242	75
rect	241	75	242	76
rect	241	77	242	78
rect	241	78	242	79
rect	241	80	242	81
rect	241	81	242	82
rect	241	83	242	84
rect	241	84	242	85
rect	241	86	242	87
rect	241	87	242	88
rect	241	89	242	90
rect	241	90	242	91
rect	241	91	242	92
rect	241	92	242	93
rect	241	93	242	94
rect	241	95	242	96
rect	241	96	242	97
rect	241	98	242	99
rect	241	99	242	100
rect	241	101	242	102
rect	241	102	242	103
rect	241	104	242	105
rect	241	105	242	106
rect	241	107	242	108
rect	241	108	242	109
rect	241	110	242	111
rect	241	111	242	112
rect	241	113	242	114
rect	241	114	242	115
rect	241	116	242	117
rect	241	117	242	118
rect	241	119	242	120
rect	241	120	242	121
rect	241	121	242	122
rect	241	122	242	123
rect	241	123	242	124
rect	241	125	242	126
rect	241	126	242	127
rect	241	128	242	129
rect	241	129	242	130
rect	241	130	242	131
rect	241	131	242	132
rect	241	132	242	133
rect	241	134	242	135
rect	241	135	242	136
rect	241	137	242	138
rect	241	138	242	139
rect	241	140	242	141
rect	241	141	242	142
rect	241	143	242	144
rect	241	144	242	145
rect	241	146	242	147
rect	241	147	242	148
rect	241	149	242	150
rect	241	150	242	151
rect	241	152	242	153
rect	241	153	242	154
rect	241	155	242	156
rect	241	156	242	157
rect	241	158	242	159
rect	241	159	242	160
rect	241	161	242	162
rect	241	162	242	163
rect	241	164	242	165
rect	241	165	242	166
rect	241	167	242	168
rect	241	168	242	169
rect	241	170	242	171
rect	241	171	242	172
rect	241	173	242	174
rect	241	174	242	175
rect	241	176	242	177
rect	241	177	242	178
rect	241	179	242	180
rect	241	180	242	181
rect	241	182	242	183
rect	241	183	242	184
rect	241	185	242	186
rect	241	186	242	187
rect	241	188	242	189
rect	241	189	242	190
rect	241	190	242	191
rect	241	191	242	192
rect	241	192	242	193
rect	241	194	242	195
rect	241	195	242	196
rect	241	197	242	198
rect	241	198	242	199
rect	241	200	242	201
rect	241	201	242	202
rect	241	203	242	204
rect	241	204	242	205
rect	241	206	242	207
rect	241	207	242	208
rect	241	209	242	210
rect	241	210	242	211
rect	241	212	242	213
rect	241	213	242	214
rect	241	215	242	216
rect	241	216	242	217
rect	241	218	242	219
rect	241	219	242	220
rect	241	221	242	222
rect	241	222	242	223
rect	241	224	242	225
rect	241	225	242	226
rect	241	227	242	228
rect	241	228	242	229
rect	241	230	242	231
rect	241	231	242	232
rect	241	233	242	234
rect	241	234	242	235
rect	241	236	242	237
rect	241	237	242	238
rect	241	239	242	240
rect	241	240	242	241
rect	241	241	242	242
rect	241	242	242	243
rect	241	243	242	244
rect	241	245	242	246
rect	241	246	242	247
rect	241	248	242	249
rect	241	249	242	250
rect	241	251	242	252
rect	241	252	242	253
rect	241	253	242	254
rect	241	254	242	255
rect	241	255	242	256
rect	241	257	242	258
rect	241	258	242	259
rect	241	260	242	261
rect	241	261	242	262
rect	241	262	242	263
rect	241	263	242	264
rect	241	264	242	265
rect	241	265	242	266
rect	241	266	242	267
rect	241	267	242	268
rect	241	268	242	269
rect	241	269	242	270
rect	241	270	242	271
rect	241	271	242	272
rect	241	272	242	273
rect	241	273	242	274
rect	241	274	242	275
rect	241	275	242	276
rect	241	276	242	277
rect	241	277	242	278
rect	241	278	242	279
rect	241	279	242	280
rect	241	280	242	281
rect	241	281	242	282
rect	241	282	242	283
rect	241	283	242	284
rect	241	284	242	285
rect	246	0	247	1
rect	246	1	247	2
rect	246	2	247	3
rect	246	3	247	4
rect	246	4	247	5
rect	246	5	247	6
rect	246	6	247	7
rect	246	8	247	9
rect	246	9	247	10
rect	246	11	247	12
rect	246	12	247	13
rect	246	14	247	15
rect	246	15	247	16
rect	246	17	247	18
rect	246	18	247	19
rect	246	20	247	21
rect	246	21	247	22
rect	246	23	247	24
rect	246	24	247	25
rect	246	26	247	27
rect	246	27	247	28
rect	246	29	247	30
rect	246	30	247	31
rect	246	32	247	33
rect	246	33	247	34
rect	246	35	247	36
rect	246	36	247	37
rect	246	38	247	39
rect	246	39	247	40
rect	246	41	247	42
rect	246	42	247	43
rect	246	44	247	45
rect	246	45	247	46
rect	246	47	247	48
rect	246	48	247	49
rect	246	50	247	51
rect	246	51	247	52
rect	246	53	247	54
rect	246	54	247	55
rect	246	56	247	57
rect	246	57	247	58
rect	246	59	247	60
rect	246	60	247	61
rect	246	62	247	63
rect	246	63	247	64
rect	246	65	247	66
rect	246	66	247	67
rect	246	68	247	69
rect	246	69	247	70
rect	246	71	247	72
rect	246	72	247	73
rect	246	74	247	75
rect	246	75	247	76
rect	246	77	247	78
rect	246	78	247	79
rect	246	80	247	81
rect	246	81	247	82
rect	246	83	247	84
rect	246	84	247	85
rect	246	86	247	87
rect	246	87	247	88
rect	246	89	247	90
rect	246	90	247	91
rect	246	91	247	92
rect	246	92	247	93
rect	246	93	247	94
rect	246	95	247	96
rect	246	96	247	97
rect	246	98	247	99
rect	246	99	247	100
rect	246	101	247	102
rect	246	102	247	103
rect	246	104	247	105
rect	246	105	247	106
rect	246	107	247	108
rect	246	108	247	109
rect	246	110	247	111
rect	246	111	247	112
rect	246	112	247	113
rect	246	113	247	114
rect	246	114	247	115
rect	246	116	247	117
rect	246	117	247	118
rect	246	119	247	120
rect	246	120	247	121
rect	246	121	247	122
rect	246	122	247	123
rect	246	123	247	124
rect	246	125	247	126
rect	246	126	247	127
rect	246	128	247	129
rect	246	129	247	130
rect	246	130	247	131
rect	246	131	247	132
rect	246	132	247	133
rect	246	134	247	135
rect	246	135	247	136
rect	246	137	247	138
rect	246	138	247	139
rect	246	140	247	141
rect	246	141	247	142
rect	246	143	247	144
rect	246	144	247	145
rect	246	146	247	147
rect	246	147	247	148
rect	246	149	247	150
rect	246	150	247	151
rect	246	152	247	153
rect	246	153	247	154
rect	246	155	247	156
rect	246	156	247	157
rect	246	158	247	159
rect	246	159	247	160
rect	246	161	247	162
rect	246	162	247	163
rect	246	164	247	165
rect	246	165	247	166
rect	246	167	247	168
rect	246	168	247	169
rect	246	170	247	171
rect	246	171	247	172
rect	246	173	247	174
rect	246	174	247	175
rect	246	176	247	177
rect	246	177	247	178
rect	246	179	247	180
rect	246	180	247	181
rect	246	182	247	183
rect	246	183	247	184
rect	246	185	247	186
rect	246	186	247	187
rect	246	188	247	189
rect	246	189	247	190
rect	246	190	247	191
rect	246	191	247	192
rect	246	192	247	193
rect	246	194	247	195
rect	246	195	247	196
rect	246	197	247	198
rect	246	198	247	199
rect	246	200	247	201
rect	246	201	247	202
rect	246	203	247	204
rect	246	204	247	205
rect	246	206	247	207
rect	246	207	247	208
rect	246	209	247	210
rect	246	210	247	211
rect	246	212	247	213
rect	246	213	247	214
rect	246	215	247	216
rect	246	216	247	217
rect	246	218	247	219
rect	246	219	247	220
rect	246	221	247	222
rect	246	222	247	223
rect	246	224	247	225
rect	246	225	247	226
rect	246	227	247	228
rect	246	228	247	229
rect	246	230	247	231
rect	246	231	247	232
rect	246	232	247	233
rect	246	233	247	234
rect	246	234	247	235
rect	246	235	247	236
rect	246	236	247	237
rect	246	237	247	238
rect	246	239	247	240
rect	246	240	247	241
rect	246	241	247	242
rect	246	242	247	243
rect	246	243	247	244
rect	246	245	247	246
rect	246	246	247	247
rect	246	248	247	249
rect	246	249	247	250
rect	246	251	247	252
rect	246	252	247	253
rect	246	253	247	254
rect	246	254	247	255
rect	246	255	247	256
rect	246	256	247	257
rect	246	257	247	258
rect	246	258	247	259
rect	246	259	247	260
rect	246	260	247	261
rect	246	261	247	262
rect	246	262	247	263
rect	246	263	247	264
rect	246	264	247	265
rect	246	265	247	266
rect	246	266	247	267
rect	246	267	247	268
rect	246	268	247	269
rect	246	269	247	270
rect	246	270	247	271
rect	246	271	247	272
rect	246	272	247	273
rect	246	273	247	274
rect	246	274	247	275
rect	246	275	247	276
rect	246	276	247	277
rect	246	277	247	278
rect	246	278	247	279
rect	246	279	247	280
rect	246	280	247	281
rect	246	281	247	282
rect	246	282	247	283
rect	246	283	247	284
rect	246	284	247	285
rect	248	0	249	1
rect	248	1	249	2
rect	248	2	249	3
rect	248	3	249	4
rect	248	4	249	5
rect	248	5	249	6
rect	248	6	249	7
rect	248	8	249	9
rect	248	9	249	10
rect	248	11	249	12
rect	248	12	249	13
rect	248	14	249	15
rect	248	15	249	16
rect	248	17	249	18
rect	248	18	249	19
rect	248	20	249	21
rect	248	21	249	22
rect	248	23	249	24
rect	248	24	249	25
rect	248	26	249	27
rect	248	27	249	28
rect	248	29	249	30
rect	248	30	249	31
rect	248	32	249	33
rect	248	33	249	34
rect	248	35	249	36
rect	248	36	249	37
rect	248	38	249	39
rect	248	39	249	40
rect	248	41	249	42
rect	248	42	249	43
rect	248	44	249	45
rect	248	45	249	46
rect	248	47	249	48
rect	248	48	249	49
rect	248	50	249	51
rect	248	51	249	52
rect	248	53	249	54
rect	248	54	249	55
rect	248	56	249	57
rect	248	57	249	58
rect	248	59	249	60
rect	248	60	249	61
rect	248	62	249	63
rect	248	63	249	64
rect	248	65	249	66
rect	248	66	249	67
rect	248	68	249	69
rect	248	69	249	70
rect	248	71	249	72
rect	248	72	249	73
rect	248	74	249	75
rect	248	75	249	76
rect	248	77	249	78
rect	248	78	249	79
rect	248	80	249	81
rect	248	81	249	82
rect	248	83	249	84
rect	248	84	249	85
rect	248	86	249	87
rect	248	87	249	88
rect	248	89	249	90
rect	248	90	249	91
rect	248	91	249	92
rect	248	92	249	93
rect	248	93	249	94
rect	248	95	249	96
rect	248	96	249	97
rect	248	98	249	99
rect	248	99	249	100
rect	248	101	249	102
rect	248	102	249	103
rect	248	104	249	105
rect	248	105	249	106
rect	248	107	249	108
rect	248	108	249	109
rect	248	110	249	111
rect	248	111	249	112
rect	248	112	249	113
rect	248	113	249	114
rect	248	114	249	115
rect	248	116	249	117
rect	248	117	249	118
rect	248	119	249	120
rect	248	120	249	121
rect	248	121	249	122
rect	248	122	249	123
rect	248	123	249	124
rect	248	125	249	126
rect	248	126	249	127
rect	248	128	249	129
rect	248	129	249	130
rect	248	130	249	131
rect	248	131	249	132
rect	248	132	249	133
rect	248	134	249	135
rect	248	135	249	136
rect	248	137	249	138
rect	248	138	249	139
rect	248	140	249	141
rect	248	141	249	142
rect	248	143	249	144
rect	248	144	249	145
rect	248	146	249	147
rect	248	147	249	148
rect	248	149	249	150
rect	248	150	249	151
rect	248	152	249	153
rect	248	153	249	154
rect	248	155	249	156
rect	248	156	249	157
rect	248	158	249	159
rect	248	159	249	160
rect	248	161	249	162
rect	248	162	249	163
rect	248	164	249	165
rect	248	165	249	166
rect	248	167	249	168
rect	248	168	249	169
rect	248	170	249	171
rect	248	171	249	172
rect	248	173	249	174
rect	248	174	249	175
rect	248	176	249	177
rect	248	177	249	178
rect	248	179	249	180
rect	248	180	249	181
rect	248	182	249	183
rect	248	183	249	184
rect	248	185	249	186
rect	248	186	249	187
rect	248	188	249	189
rect	248	189	249	190
rect	248	190	249	191
rect	248	191	249	192
rect	248	192	249	193
rect	248	194	249	195
rect	248	195	249	196
rect	248	197	249	198
rect	248	198	249	199
rect	248	200	249	201
rect	248	201	249	202
rect	248	203	249	204
rect	248	204	249	205
rect	248	206	249	207
rect	248	207	249	208
rect	248	209	249	210
rect	248	210	249	211
rect	248	212	249	213
rect	248	213	249	214
rect	248	215	249	216
rect	248	216	249	217
rect	248	218	249	219
rect	248	219	249	220
rect	248	221	249	222
rect	248	222	249	223
rect	248	224	249	225
rect	248	225	249	226
rect	248	227	249	228
rect	248	228	249	229
rect	248	230	249	231
rect	248	231	249	232
rect	248	232	249	233
rect	248	233	249	234
rect	248	234	249	235
rect	248	235	249	236
rect	248	236	249	237
rect	248	237	249	238
rect	248	239	249	240
rect	248	240	249	241
rect	248	241	249	242
rect	248	242	249	243
rect	248	243	249	244
rect	248	245	249	246
rect	248	246	249	247
rect	248	248	249	249
rect	248	249	249	250
rect	248	251	249	252
rect	248	252	249	253
rect	248	253	249	254
rect	248	254	249	255
rect	248	255	249	256
rect	248	256	249	257
rect	248	257	249	258
rect	248	258	249	259
rect	248	259	249	260
rect	248	260	249	261
rect	248	261	249	262
rect	248	262	249	263
rect	248	263	249	264
rect	248	264	249	265
rect	248	265	249	266
rect	248	266	249	267
rect	248	267	249	268
rect	248	268	249	269
rect	248	269	249	270
rect	249	0	250	1
rect	249	1	250	2
rect	249	2	250	3
rect	249	3	250	4
rect	249	4	250	5
rect	249	5	250	6
rect	249	6	250	7
rect	249	8	250	9
rect	249	9	250	10
rect	249	11	250	12
rect	249	12	250	13
rect	249	14	250	15
rect	249	15	250	16
rect	249	17	250	18
rect	249	18	250	19
rect	249	20	250	21
rect	249	21	250	22
rect	249	23	250	24
rect	249	24	250	25
rect	249	26	250	27
rect	249	27	250	28
rect	249	29	250	30
rect	249	30	250	31
rect	249	32	250	33
rect	249	33	250	34
rect	249	35	250	36
rect	249	36	250	37
rect	249	38	250	39
rect	249	39	250	40
rect	249	41	250	42
rect	249	42	250	43
rect	249	44	250	45
rect	249	45	250	46
rect	249	47	250	48
rect	249	48	250	49
rect	249	50	250	51
rect	249	51	250	52
rect	249	53	250	54
rect	249	54	250	55
rect	249	56	250	57
rect	249	57	250	58
rect	249	59	250	60
rect	249	60	250	61
rect	249	62	250	63
rect	249	63	250	64
rect	249	65	250	66
rect	249	66	250	67
rect	249	68	250	69
rect	249	69	250	70
rect	249	71	250	72
rect	249	72	250	73
rect	249	74	250	75
rect	249	75	250	76
rect	249	77	250	78
rect	249	78	250	79
rect	249	80	250	81
rect	249	81	250	82
rect	249	83	250	84
rect	249	84	250	85
rect	249	86	250	87
rect	249	87	250	88
rect	249	89	250	90
rect	249	90	250	91
rect	249	91	250	92
rect	249	92	250	93
rect	249	93	250	94
rect	249	95	250	96
rect	249	96	250	97
rect	249	98	250	99
rect	249	99	250	100
rect	249	101	250	102
rect	249	102	250	103
rect	249	104	250	105
rect	249	105	250	106
rect	249	107	250	108
rect	249	108	250	109
rect	249	110	250	111
rect	249	111	250	112
rect	249	112	250	113
rect	249	113	250	114
rect	249	114	250	115
rect	249	116	250	117
rect	249	117	250	118
rect	249	119	250	120
rect	249	120	250	121
rect	249	121	250	122
rect	249	122	250	123
rect	249	123	250	124
rect	249	125	250	126
rect	249	126	250	127
rect	249	128	250	129
rect	249	129	250	130
rect	249	130	250	131
rect	249	131	250	132
rect	249	132	250	133
rect	249	134	250	135
rect	249	135	250	136
rect	249	137	250	138
rect	249	138	250	139
rect	249	140	250	141
rect	249	141	250	142
rect	249	143	250	144
rect	249	144	250	145
rect	249	146	250	147
rect	249	147	250	148
rect	249	149	250	150
rect	249	150	250	151
rect	249	152	250	153
rect	249	153	250	154
rect	249	155	250	156
rect	249	156	250	157
rect	249	158	250	159
rect	249	159	250	160
rect	249	161	250	162
rect	249	162	250	163
rect	249	164	250	165
rect	249	165	250	166
rect	249	167	250	168
rect	249	168	250	169
rect	249	170	250	171
rect	249	171	250	172
rect	249	173	250	174
rect	249	174	250	175
rect	249	176	250	177
rect	249	177	250	178
rect	249	179	250	180
rect	249	180	250	181
rect	249	182	250	183
rect	249	183	250	184
rect	249	185	250	186
rect	249	186	250	187
rect	249	188	250	189
rect	249	189	250	190
rect	249	190	250	191
rect	249	191	250	192
rect	249	192	250	193
rect	249	194	250	195
rect	249	195	250	196
rect	249	197	250	198
rect	249	198	250	199
rect	249	200	250	201
rect	249	201	250	202
rect	249	203	250	204
rect	249	204	250	205
rect	249	206	250	207
rect	249	207	250	208
rect	249	209	250	210
rect	249	210	250	211
rect	249	212	250	213
rect	249	213	250	214
rect	249	215	250	216
rect	249	216	250	217
rect	249	218	250	219
rect	249	219	250	220
rect	249	221	250	222
rect	249	222	250	223
rect	249	224	250	225
rect	249	225	250	226
rect	249	227	250	228
rect	249	228	250	229
rect	249	230	250	231
rect	249	231	250	232
rect	249	232	250	233
rect	249	233	250	234
rect	249	234	250	235
rect	249	235	250	236
rect	249	236	250	237
rect	249	237	250	238
rect	249	239	250	240
rect	249	240	250	241
rect	249	241	250	242
rect	249	242	250	243
rect	249	243	250	244
rect	249	245	250	246
rect	249	246	250	247
rect	249	248	250	249
rect	249	249	250	250
rect	249	251	250	252
rect	249	252	250	253
rect	249	253	250	254
rect	249	254	250	255
rect	249	255	250	256
rect	249	256	250	257
rect	249	257	250	258
rect	249	258	250	259
rect	249	259	250	260
rect	249	260	250	261
rect	249	261	250	262
rect	249	262	250	263
rect	249	263	250	264
rect	249	264	250	265
rect	249	265	250	266
rect	249	266	250	267
rect	249	267	250	268
rect	249	268	250	269
rect	249	269	250	270
rect	250	0	251	1
rect	250	1	251	2
rect	250	2	251	3
rect	250	3	251	4
rect	250	4	251	5
rect	250	5	251	6
rect	250	6	251	7
rect	250	8	251	9
rect	250	9	251	10
rect	250	11	251	12
rect	250	12	251	13
rect	250	14	251	15
rect	250	15	251	16
rect	250	17	251	18
rect	250	18	251	19
rect	250	20	251	21
rect	250	21	251	22
rect	250	23	251	24
rect	250	24	251	25
rect	250	26	251	27
rect	250	27	251	28
rect	250	29	251	30
rect	250	30	251	31
rect	250	32	251	33
rect	250	33	251	34
rect	250	35	251	36
rect	250	36	251	37
rect	250	38	251	39
rect	250	39	251	40
rect	250	41	251	42
rect	250	42	251	43
rect	250	44	251	45
rect	250	45	251	46
rect	250	47	251	48
rect	250	48	251	49
rect	250	50	251	51
rect	250	51	251	52
rect	250	53	251	54
rect	250	54	251	55
rect	250	56	251	57
rect	250	57	251	58
rect	250	59	251	60
rect	250	60	251	61
rect	250	62	251	63
rect	250	63	251	64
rect	250	65	251	66
rect	250	66	251	67
rect	250	68	251	69
rect	250	69	251	70
rect	250	71	251	72
rect	250	72	251	73
rect	250	74	251	75
rect	250	75	251	76
rect	250	77	251	78
rect	250	78	251	79
rect	250	80	251	81
rect	250	81	251	82
rect	250	83	251	84
rect	250	84	251	85
rect	250	86	251	87
rect	250	87	251	88
rect	250	89	251	90
rect	250	90	251	91
rect	250	91	251	92
rect	250	92	251	93
rect	250	93	251	94
rect	250	95	251	96
rect	250	96	251	97
rect	250	98	251	99
rect	250	99	251	100
rect	250	101	251	102
rect	250	102	251	103
rect	250	104	251	105
rect	250	105	251	106
rect	250	107	251	108
rect	250	108	251	109
rect	250	110	251	111
rect	250	111	251	112
rect	250	112	251	113
rect	250	113	251	114
rect	250	114	251	115
rect	250	116	251	117
rect	250	117	251	118
rect	250	119	251	120
rect	250	120	251	121
rect	250	121	251	122
rect	250	122	251	123
rect	250	123	251	124
rect	250	125	251	126
rect	250	126	251	127
rect	250	128	251	129
rect	250	129	251	130
rect	250	130	251	131
rect	250	131	251	132
rect	250	132	251	133
rect	250	134	251	135
rect	250	135	251	136
rect	250	137	251	138
rect	250	138	251	139
rect	250	140	251	141
rect	250	141	251	142
rect	250	143	251	144
rect	250	144	251	145
rect	250	146	251	147
rect	250	147	251	148
rect	250	149	251	150
rect	250	150	251	151
rect	250	152	251	153
rect	250	153	251	154
rect	250	154	251	155
rect	250	155	251	156
rect	250	156	251	157
rect	250	158	251	159
rect	250	159	251	160
rect	250	161	251	162
rect	250	162	251	163
rect	250	164	251	165
rect	250	165	251	166
rect	250	167	251	168
rect	250	168	251	169
rect	250	170	251	171
rect	250	171	251	172
rect	250	173	251	174
rect	250	174	251	175
rect	250	176	251	177
rect	250	177	251	178
rect	250	179	251	180
rect	250	180	251	181
rect	250	182	251	183
rect	250	183	251	184
rect	250	185	251	186
rect	250	186	251	187
rect	250	188	251	189
rect	250	189	251	190
rect	250	190	251	191
rect	250	191	251	192
rect	250	192	251	193
rect	250	194	251	195
rect	250	195	251	196
rect	250	197	251	198
rect	250	198	251	199
rect	250	200	251	201
rect	250	201	251	202
rect	250	203	251	204
rect	250	204	251	205
rect	250	206	251	207
rect	250	207	251	208
rect	250	209	251	210
rect	250	210	251	211
rect	250	212	251	213
rect	250	213	251	214
rect	250	215	251	216
rect	250	216	251	217
rect	250	218	251	219
rect	250	219	251	220
rect	250	221	251	222
rect	250	222	251	223
rect	250	224	251	225
rect	250	225	251	226
rect	250	227	251	228
rect	250	228	251	229
rect	250	230	251	231
rect	250	231	251	232
rect	250	232	251	233
rect	250	233	251	234
rect	250	234	251	235
rect	250	235	251	236
rect	250	236	251	237
rect	250	237	251	238
rect	250	239	251	240
rect	250	240	251	241
rect	250	241	251	242
rect	250	242	251	243
rect	250	243	251	244
rect	250	244	251	245
rect	250	245	251	246
rect	250	246	251	247
rect	250	248	251	249
rect	250	249	251	250
rect	250	250	251	251
rect	250	251	251	252
rect	250	252	251	253
rect	250	253	251	254
rect	250	254	251	255
rect	250	255	251	256
rect	250	256	251	257
rect	250	257	251	258
rect	250	258	251	259
rect	250	259	251	260
rect	250	260	251	261
rect	250	261	251	262
rect	250	262	251	263
rect	250	263	251	264
rect	250	264	251	265
rect	250	265	251	266
rect	250	266	251	267
rect	250	267	251	268
rect	250	268	251	269
rect	250	269	251	270
rect	251	0	252	1
rect	251	1	252	2
rect	251	2	252	3
rect	251	3	252	4
rect	251	4	252	5
rect	251	5	252	6
rect	251	6	252	7
rect	251	8	252	9
rect	251	9	252	10
rect	251	11	252	12
rect	251	12	252	13
rect	251	14	252	15
rect	251	15	252	16
rect	251	17	252	18
rect	251	18	252	19
rect	251	20	252	21
rect	251	21	252	22
rect	251	23	252	24
rect	251	24	252	25
rect	251	26	252	27
rect	251	27	252	28
rect	251	29	252	30
rect	251	30	252	31
rect	251	32	252	33
rect	251	33	252	34
rect	251	35	252	36
rect	251	36	252	37
rect	251	38	252	39
rect	251	39	252	40
rect	251	41	252	42
rect	251	42	252	43
rect	251	44	252	45
rect	251	45	252	46
rect	251	47	252	48
rect	251	48	252	49
rect	251	50	252	51
rect	251	51	252	52
rect	251	53	252	54
rect	251	54	252	55
rect	251	56	252	57
rect	251	57	252	58
rect	251	59	252	60
rect	251	60	252	61
rect	251	62	252	63
rect	251	63	252	64
rect	251	65	252	66
rect	251	66	252	67
rect	251	68	252	69
rect	251	69	252	70
rect	251	71	252	72
rect	251	72	252	73
rect	251	74	252	75
rect	251	75	252	76
rect	251	77	252	78
rect	251	78	252	79
rect	251	80	252	81
rect	251	81	252	82
rect	251	83	252	84
rect	251	84	252	85
rect	251	86	252	87
rect	251	87	252	88
rect	251	89	252	90
rect	251	90	252	91
rect	251	91	252	92
rect	251	92	252	93
rect	251	93	252	94
rect	251	95	252	96
rect	251	96	252	97
rect	251	98	252	99
rect	251	99	252	100
rect	251	101	252	102
rect	251	102	252	103
rect	251	104	252	105
rect	251	105	252	106
rect	251	107	252	108
rect	251	108	252	109
rect	251	110	252	111
rect	251	111	252	112
rect	251	112	252	113
rect	251	113	252	114
rect	251	114	252	115
rect	251	116	252	117
rect	251	117	252	118
rect	251	119	252	120
rect	251	120	252	121
rect	251	121	252	122
rect	251	122	252	123
rect	251	123	252	124
rect	251	125	252	126
rect	251	126	252	127
rect	251	128	252	129
rect	251	129	252	130
rect	251	130	252	131
rect	251	131	252	132
rect	251	132	252	133
rect	251	134	252	135
rect	251	135	252	136
rect	251	137	252	138
rect	251	138	252	139
rect	251	140	252	141
rect	251	141	252	142
rect	251	143	252	144
rect	251	144	252	145
rect	251	146	252	147
rect	251	147	252	148
rect	251	149	252	150
rect	251	150	252	151
rect	251	152	252	153
rect	251	153	252	154
rect	251	154	252	155
rect	251	155	252	156
rect	251	156	252	157
rect	251	158	252	159
rect	251	159	252	160
rect	251	161	252	162
rect	251	162	252	163
rect	251	164	252	165
rect	251	165	252	166
rect	251	167	252	168
rect	251	168	252	169
rect	251	170	252	171
rect	251	171	252	172
rect	251	173	252	174
rect	251	174	252	175
rect	251	176	252	177
rect	251	177	252	178
rect	251	179	252	180
rect	251	180	252	181
rect	251	182	252	183
rect	251	183	252	184
rect	251	185	252	186
rect	251	186	252	187
rect	251	188	252	189
rect	251	189	252	190
rect	251	190	252	191
rect	251	191	252	192
rect	251	192	252	193
rect	251	194	252	195
rect	251	195	252	196
rect	251	197	252	198
rect	251	198	252	199
rect	251	200	252	201
rect	251	201	252	202
rect	251	203	252	204
rect	251	204	252	205
rect	251	206	252	207
rect	251	207	252	208
rect	251	209	252	210
rect	251	210	252	211
rect	251	212	252	213
rect	251	213	252	214
rect	251	215	252	216
rect	251	216	252	217
rect	251	218	252	219
rect	251	219	252	220
rect	251	221	252	222
rect	251	222	252	223
rect	251	224	252	225
rect	251	225	252	226
rect	251	227	252	228
rect	251	228	252	229
rect	251	230	252	231
rect	251	231	252	232
rect	251	232	252	233
rect	251	233	252	234
rect	251	234	252	235
rect	251	236	252	237
rect	251	237	252	238
rect	251	239	252	240
rect	251	240	252	241
rect	251	241	252	242
rect	251	242	252	243
rect	251	243	252	244
rect	251	244	252	245
rect	251	245	252	246
rect	251	246	252	247
rect	251	248	252	249
rect	251	249	252	250
rect	251	250	252	251
rect	251	251	252	252
rect	251	252	252	253
rect	251	253	252	254
rect	251	254	252	255
rect	251	255	252	256
rect	251	256	252	257
rect	251	257	252	258
rect	251	258	252	259
rect	251	259	252	260
rect	251	260	252	261
rect	251	261	252	262
rect	251	262	252	263
rect	251	263	252	264
rect	251	264	252	265
rect	251	265	252	266
rect	251	266	252	267
rect	251	267	252	268
rect	251	268	252	269
rect	251	269	252	270
rect	252	0	253	1
rect	252	1	253	2
rect	252	2	253	3
rect	252	3	253	4
rect	252	4	253	5
rect	252	5	253	6
rect	252	6	253	7
rect	252	8	253	9
rect	252	9	253	10
rect	252	11	253	12
rect	252	12	253	13
rect	252	14	253	15
rect	252	15	253	16
rect	252	17	253	18
rect	252	18	253	19
rect	252	20	253	21
rect	252	21	253	22
rect	252	23	253	24
rect	252	24	253	25
rect	252	26	253	27
rect	252	27	253	28
rect	252	29	253	30
rect	252	30	253	31
rect	252	32	253	33
rect	252	33	253	34
rect	252	35	253	36
rect	252	36	253	37
rect	252	38	253	39
rect	252	39	253	40
rect	252	41	253	42
rect	252	42	253	43
rect	252	44	253	45
rect	252	45	253	46
rect	252	47	253	48
rect	252	48	253	49
rect	252	50	253	51
rect	252	51	253	52
rect	252	53	253	54
rect	252	54	253	55
rect	252	56	253	57
rect	252	57	253	58
rect	252	59	253	60
rect	252	60	253	61
rect	252	62	253	63
rect	252	63	253	64
rect	252	65	253	66
rect	252	66	253	67
rect	252	68	253	69
rect	252	69	253	70
rect	252	71	253	72
rect	252	72	253	73
rect	252	74	253	75
rect	252	75	253	76
rect	252	77	253	78
rect	252	78	253	79
rect	252	80	253	81
rect	252	81	253	82
rect	252	83	253	84
rect	252	84	253	85
rect	252	86	253	87
rect	252	87	253	88
rect	252	89	253	90
rect	252	90	253	91
rect	252	91	253	92
rect	252	92	253	93
rect	252	93	253	94
rect	252	95	253	96
rect	252	96	253	97
rect	252	98	253	99
rect	252	99	253	100
rect	252	101	253	102
rect	252	102	253	103
rect	252	104	253	105
rect	252	105	253	106
rect	252	107	253	108
rect	252	108	253	109
rect	252	110	253	111
rect	252	111	253	112
rect	252	112	253	113
rect	252	113	253	114
rect	252	114	253	115
rect	252	116	253	117
rect	252	117	253	118
rect	252	119	253	120
rect	252	120	253	121
rect	252	121	253	122
rect	252	122	253	123
rect	252	123	253	124
rect	252	125	253	126
rect	252	126	253	127
rect	252	128	253	129
rect	252	129	253	130
rect	252	130	253	131
rect	252	131	253	132
rect	252	132	253	133
rect	252	134	253	135
rect	252	135	253	136
rect	252	137	253	138
rect	252	138	253	139
rect	252	140	253	141
rect	252	141	253	142
rect	252	143	253	144
rect	252	144	253	145
rect	252	146	253	147
rect	252	147	253	148
rect	252	149	253	150
rect	252	150	253	151
rect	252	152	253	153
rect	252	153	253	154
rect	252	154	253	155
rect	252	155	253	156
rect	252	156	253	157
rect	252	158	253	159
rect	252	159	253	160
rect	252	161	253	162
rect	252	162	253	163
rect	252	164	253	165
rect	252	165	253	166
rect	252	167	253	168
rect	252	168	253	169
rect	252	170	253	171
rect	252	171	253	172
rect	252	173	253	174
rect	252	174	253	175
rect	252	176	253	177
rect	252	177	253	178
rect	252	179	253	180
rect	252	180	253	181
rect	252	182	253	183
rect	252	183	253	184
rect	252	185	253	186
rect	252	186	253	187
rect	252	188	253	189
rect	252	189	253	190
rect	252	190	253	191
rect	252	191	253	192
rect	252	192	253	193
rect	252	194	253	195
rect	252	195	253	196
rect	252	197	253	198
rect	252	198	253	199
rect	252	200	253	201
rect	252	201	253	202
rect	252	203	253	204
rect	252	204	253	205
rect	252	206	253	207
rect	252	207	253	208
rect	252	209	253	210
rect	252	210	253	211
rect	252	212	253	213
rect	252	213	253	214
rect	252	215	253	216
rect	252	216	253	217
rect	252	218	253	219
rect	252	219	253	220
rect	252	221	253	222
rect	252	222	253	223
rect	252	224	253	225
rect	252	225	253	226
rect	252	227	253	228
rect	252	228	253	229
rect	252	230	253	231
rect	252	231	253	232
rect	252	232	253	233
rect	252	233	253	234
rect	252	234	253	235
rect	252	236	253	237
rect	252	237	253	238
rect	252	239	253	240
rect	252	240	253	241
rect	252	241	253	242
rect	252	242	253	243
rect	252	243	253	244
rect	252	244	253	245
rect	252	245	253	246
rect	252	246	253	247
rect	252	248	253	249
rect	252	249	253	250
rect	252	250	253	251
rect	252	251	253	252
rect	252	252	253	253
rect	252	253	253	254
rect	252	254	253	255
rect	252	255	253	256
rect	252	256	253	257
rect	252	257	253	258
rect	252	258	253	259
rect	252	259	253	260
rect	252	260	253	261
rect	252	261	253	262
rect	252	262	253	263
rect	252	263	253	264
rect	252	264	253	265
rect	252	265	253	266
rect	252	266	253	267
rect	252	267	253	268
rect	252	268	253	269
rect	252	269	253	270
rect	255	0	256	1
rect	255	1	256	2
rect	255	2	256	3
rect	255	3	256	4
rect	255	4	256	5
rect	255	5	256	6
rect	255	6	256	7
rect	255	8	256	9
rect	255	9	256	10
rect	255	11	256	12
rect	255	12	256	13
rect	255	14	256	15
rect	255	15	256	16
rect	255	17	256	18
rect	255	18	256	19
rect	255	20	256	21
rect	255	21	256	22
rect	255	23	256	24
rect	255	24	256	25
rect	255	26	256	27
rect	255	27	256	28
rect	255	29	256	30
rect	255	30	256	31
rect	255	32	256	33
rect	255	33	256	34
rect	255	35	256	36
rect	255	36	256	37
rect	255	38	256	39
rect	255	39	256	40
rect	255	41	256	42
rect	255	42	256	43
rect	255	44	256	45
rect	255	45	256	46
rect	255	47	256	48
rect	255	48	256	49
rect	255	50	256	51
rect	255	51	256	52
rect	255	53	256	54
rect	255	54	256	55
rect	255	56	256	57
rect	255	57	256	58
rect	255	59	256	60
rect	255	60	256	61
rect	255	62	256	63
rect	255	63	256	64
rect	255	65	256	66
rect	255	66	256	67
rect	255	68	256	69
rect	255	69	256	70
rect	255	70	256	71
rect	255	71	256	72
rect	255	72	256	73
rect	255	73	256	74
rect	255	74	256	75
rect	255	75	256	76
rect	255	76	256	77
rect	255	77	256	78
rect	255	78	256	79
rect	255	80	256	81
rect	255	81	256	82
rect	255	83	256	84
rect	255	84	256	85
rect	255	86	256	87
rect	255	87	256	88
rect	255	89	256	90
rect	255	90	256	91
rect	255	91	256	92
rect	255	92	256	93
rect	255	93	256	94
rect	255	94	256	95
rect	255	95	256	96
rect	255	96	256	97
rect	255	98	256	99
rect	255	99	256	100
rect	255	101	256	102
rect	255	102	256	103
rect	255	104	256	105
rect	255	105	256	106
rect	255	106	256	107
rect	255	107	256	108
rect	255	108	256	109
rect	255	110	256	111
rect	255	111	256	112
rect	255	112	256	113
rect	255	113	256	114
rect	255	114	256	115
rect	255	116	256	117
rect	255	117	256	118
rect	255	119	256	120
rect	255	120	256	121
rect	255	121	256	122
rect	255	122	256	123
rect	255	123	256	124
rect	255	125	256	126
rect	255	126	256	127
rect	255	128	256	129
rect	255	129	256	130
rect	255	130	256	131
rect	255	131	256	132
rect	255	132	256	133
rect	255	134	256	135
rect	255	135	256	136
rect	255	137	256	138
rect	255	138	256	139
rect	255	140	256	141
rect	255	141	256	142
rect	255	143	256	144
rect	255	144	256	145
rect	255	145	256	146
rect	255	146	256	147
rect	255	147	256	148
rect	255	149	256	150
rect	255	150	256	151
rect	255	152	256	153
rect	255	153	256	154
rect	255	154	256	155
rect	255	155	256	156
rect	255	156	256	157
rect	255	158	256	159
rect	255	159	256	160
rect	255	161	256	162
rect	255	162	256	163
rect	255	164	256	165
rect	255	165	256	166
rect	255	167	256	168
rect	255	168	256	169
rect	255	170	256	171
rect	255	171	256	172
rect	255	173	256	174
rect	255	174	256	175
rect	255	176	256	177
rect	255	177	256	178
rect	255	179	256	180
rect	255	180	256	181
rect	255	182	256	183
rect	255	183	256	184
rect	255	185	256	186
rect	255	186	256	187
rect	255	188	256	189
rect	255	189	256	190
rect	255	190	256	191
rect	255	191	256	192
rect	255	192	256	193
rect	255	194	256	195
rect	255	195	256	196
rect	255	197	256	198
rect	255	198	256	199
rect	255	200	256	201
rect	255	201	256	202
rect	255	203	256	204
rect	255	204	256	205
rect	255	206	256	207
rect	255	207	256	208
rect	255	209	256	210
rect	255	210	256	211
rect	255	212	256	213
rect	255	213	256	214
rect	255	214	256	215
rect	255	215	256	216
rect	255	216	256	217
rect	255	218	256	219
rect	255	219	256	220
rect	255	221	256	222
rect	255	222	256	223
rect	255	224	256	225
rect	255	225	256	226
rect	255	226	256	227
rect	255	227	256	228
rect	255	228	256	229
rect	255	229	256	230
rect	255	230	256	231
rect	255	231	256	232
rect	255	232	256	233
rect	255	233	256	234
rect	255	234	256	235
rect	255	235	256	236
rect	255	236	256	237
rect	255	237	256	238
rect	255	239	256	240
rect	255	240	256	241
rect	255	241	256	242
rect	255	242	256	243
rect	255	243	256	244
rect	255	244	256	245
rect	255	245	256	246
rect	255	246	256	247
rect	255	247	256	248
rect	255	248	256	249
rect	255	249	256	250
rect	255	250	256	251
rect	255	251	256	252
rect	255	252	256	253
rect	255	253	256	254
rect	255	254	256	255
rect	255	255	256	256
rect	255	256	256	257
rect	255	257	256	258
rect	255	258	256	259
rect	255	259	256	260
rect	255	260	256	261
rect	255	261	256	262
rect	255	262	256	263
rect	255	263	256	264
rect	255	264	256	265
rect	255	265	256	266
rect	255	266	256	267
rect	255	267	256	268
rect	255	268	256	269
rect	255	269	256	270
rect	257	0	258	1
rect	257	1	258	2
rect	257	2	258	3
rect	257	3	258	4
rect	257	4	258	5
rect	257	5	258	6
rect	257	6	258	7
rect	257	8	258	9
rect	257	9	258	10
rect	257	11	258	12
rect	257	12	258	13
rect	257	14	258	15
rect	257	15	258	16
rect	257	17	258	18
rect	257	18	258	19
rect	257	20	258	21
rect	257	21	258	22
rect	257	23	258	24
rect	257	24	258	25
rect	257	26	258	27
rect	257	27	258	28
rect	257	29	258	30
rect	257	30	258	31
rect	257	32	258	33
rect	257	33	258	34
rect	257	35	258	36
rect	257	36	258	37
rect	257	38	258	39
rect	257	39	258	40
rect	257	41	258	42
rect	257	42	258	43
rect	257	44	258	45
rect	257	45	258	46
rect	257	47	258	48
rect	257	48	258	49
rect	257	50	258	51
rect	257	51	258	52
rect	257	53	258	54
rect	257	54	258	55
rect	257	56	258	57
rect	257	57	258	58
rect	257	59	258	60
rect	257	60	258	61
rect	257	62	258	63
rect	257	63	258	64
rect	257	65	258	66
rect	257	66	258	67
rect	257	68	258	69
rect	257	69	258	70
rect	257	70	258	71
rect	257	71	258	72
rect	257	72	258	73
rect	257	73	258	74
rect	257	74	258	75
rect	257	75	258	76
rect	257	76	258	77
rect	257	77	258	78
rect	257	78	258	79
rect	257	80	258	81
rect	257	81	258	82
rect	257	83	258	84
rect	257	84	258	85
rect	257	86	258	87
rect	257	87	258	88
rect	257	89	258	90
rect	257	90	258	91
rect	257	91	258	92
rect	257	92	258	93
rect	257	93	258	94
rect	257	94	258	95
rect	257	95	258	96
rect	257	96	258	97
rect	257	98	258	99
rect	257	99	258	100
rect	257	101	258	102
rect	257	102	258	103
rect	257	104	258	105
rect	257	105	258	106
rect	257	106	258	107
rect	257	107	258	108
rect	257	108	258	109
rect	257	110	258	111
rect	257	111	258	112
rect	257	112	258	113
rect	257	113	258	114
rect	257	114	258	115
rect	257	116	258	117
rect	257	117	258	118
rect	257	119	258	120
rect	257	120	258	121
rect	257	121	258	122
rect	257	122	258	123
rect	257	123	258	124
rect	257	125	258	126
rect	257	126	258	127
rect	257	128	258	129
rect	257	129	258	130
rect	257	130	258	131
rect	257	131	258	132
rect	257	132	258	133
rect	257	134	258	135
rect	257	135	258	136
rect	257	137	258	138
rect	257	138	258	139
rect	257	140	258	141
rect	257	141	258	142
rect	257	143	258	144
rect	257	144	258	145
rect	257	145	258	146
rect	257	146	258	147
rect	257	147	258	148
rect	257	149	258	150
rect	257	150	258	151
rect	257	152	258	153
rect	257	153	258	154
rect	257	154	258	155
rect	257	155	258	156
rect	257	156	258	157
rect	257	158	258	159
rect	257	159	258	160
rect	257	161	258	162
rect	257	162	258	163
rect	257	164	258	165
rect	257	165	258	166
rect	257	167	258	168
rect	257	168	258	169
rect	257	170	258	171
rect	257	171	258	172
rect	257	173	258	174
rect	257	174	258	175
rect	257	176	258	177
rect	257	177	258	178
rect	257	179	258	180
rect	257	180	258	181
rect	257	182	258	183
rect	257	183	258	184
rect	257	185	258	186
rect	257	186	258	187
rect	257	188	258	189
rect	257	189	258	190
rect	257	190	258	191
rect	257	191	258	192
rect	257	192	258	193
rect	257	194	258	195
rect	257	195	258	196
rect	257	197	258	198
rect	257	198	258	199
rect	257	200	258	201
rect	257	201	258	202
rect	257	203	258	204
rect	257	204	258	205
rect	257	206	258	207
rect	257	207	258	208
rect	257	209	258	210
rect	257	210	258	211
rect	257	212	258	213
rect	257	213	258	214
rect	257	214	258	215
rect	257	215	258	216
rect	257	216	258	217
rect	257	218	258	219
rect	257	219	258	220
rect	257	221	258	222
rect	257	222	258	223
rect	257	224	258	225
rect	257	225	258	226
rect	257	226	258	227
rect	257	227	258	228
rect	257	228	258	229
rect	257	229	258	230
rect	257	230	258	231
rect	257	231	258	232
rect	257	232	258	233
rect	257	233	258	234
rect	257	234	258	235
rect	257	235	258	236
rect	257	236	258	237
rect	257	237	258	238
rect	257	239	258	240
rect	257	240	258	241
rect	257	241	258	242
rect	257	242	258	243
rect	257	243	258	244
rect	257	244	258	245
rect	257	245	258	246
rect	257	246	258	247
rect	257	247	258	248
rect	257	248	258	249
rect	257	249	258	250
rect	257	250	258	251
rect	257	251	258	252
rect	258	0	259	1
rect	258	1	259	2
rect	258	2	259	3
rect	258	3	259	4
rect	258	4	259	5
rect	258	5	259	6
rect	258	6	259	7
rect	258	8	259	9
rect	258	9	259	10
rect	258	11	259	12
rect	258	12	259	13
rect	258	14	259	15
rect	258	15	259	16
rect	258	17	259	18
rect	258	18	259	19
rect	258	20	259	21
rect	258	21	259	22
rect	258	23	259	24
rect	258	24	259	25
rect	258	26	259	27
rect	258	27	259	28
rect	258	29	259	30
rect	258	30	259	31
rect	258	32	259	33
rect	258	33	259	34
rect	258	35	259	36
rect	258	36	259	37
rect	258	38	259	39
rect	258	39	259	40
rect	258	41	259	42
rect	258	42	259	43
rect	258	44	259	45
rect	258	45	259	46
rect	258	47	259	48
rect	258	48	259	49
rect	258	50	259	51
rect	258	51	259	52
rect	258	53	259	54
rect	258	54	259	55
rect	258	56	259	57
rect	258	57	259	58
rect	258	59	259	60
rect	258	60	259	61
rect	258	62	259	63
rect	258	63	259	64
rect	258	65	259	66
rect	258	66	259	67
rect	258	68	259	69
rect	258	69	259	70
rect	258	70	259	71
rect	258	71	259	72
rect	258	72	259	73
rect	258	73	259	74
rect	258	74	259	75
rect	258	75	259	76
rect	258	76	259	77
rect	258	77	259	78
rect	258	78	259	79
rect	258	80	259	81
rect	258	81	259	82
rect	258	83	259	84
rect	258	84	259	85
rect	258	86	259	87
rect	258	87	259	88
rect	258	89	259	90
rect	258	90	259	91
rect	258	91	259	92
rect	258	92	259	93
rect	258	93	259	94
rect	258	94	259	95
rect	258	95	259	96
rect	258	96	259	97
rect	258	98	259	99
rect	258	99	259	100
rect	258	101	259	102
rect	258	102	259	103
rect	258	104	259	105
rect	258	105	259	106
rect	258	106	259	107
rect	258	107	259	108
rect	258	108	259	109
rect	258	110	259	111
rect	258	111	259	112
rect	258	112	259	113
rect	258	113	259	114
rect	258	114	259	115
rect	258	116	259	117
rect	258	117	259	118
rect	258	119	259	120
rect	258	120	259	121
rect	258	121	259	122
rect	258	122	259	123
rect	258	123	259	124
rect	258	125	259	126
rect	258	126	259	127
rect	258	128	259	129
rect	258	129	259	130
rect	258	130	259	131
rect	258	131	259	132
rect	258	132	259	133
rect	258	134	259	135
rect	258	135	259	136
rect	258	137	259	138
rect	258	138	259	139
rect	258	140	259	141
rect	258	141	259	142
rect	258	143	259	144
rect	258	144	259	145
rect	258	145	259	146
rect	258	146	259	147
rect	258	147	259	148
rect	258	149	259	150
rect	258	150	259	151
rect	258	152	259	153
rect	258	153	259	154
rect	258	154	259	155
rect	258	155	259	156
rect	258	156	259	157
rect	258	158	259	159
rect	258	159	259	160
rect	258	161	259	162
rect	258	162	259	163
rect	258	164	259	165
rect	258	165	259	166
rect	258	167	259	168
rect	258	168	259	169
rect	258	170	259	171
rect	258	171	259	172
rect	258	173	259	174
rect	258	174	259	175
rect	258	176	259	177
rect	258	177	259	178
rect	258	179	259	180
rect	258	180	259	181
rect	258	182	259	183
rect	258	183	259	184
rect	258	185	259	186
rect	258	186	259	187
rect	258	188	259	189
rect	258	189	259	190
rect	258	190	259	191
rect	258	191	259	192
rect	258	192	259	193
rect	258	194	259	195
rect	258	195	259	196
rect	258	197	259	198
rect	258	198	259	199
rect	258	200	259	201
rect	258	201	259	202
rect	258	203	259	204
rect	258	204	259	205
rect	258	206	259	207
rect	258	207	259	208
rect	258	209	259	210
rect	258	210	259	211
rect	258	212	259	213
rect	258	213	259	214
rect	258	214	259	215
rect	258	215	259	216
rect	258	216	259	217
rect	258	218	259	219
rect	258	219	259	220
rect	258	221	259	222
rect	258	222	259	223
rect	258	224	259	225
rect	258	225	259	226
rect	258	226	259	227
rect	258	227	259	228
rect	258	228	259	229
rect	258	229	259	230
rect	258	230	259	231
rect	258	231	259	232
rect	258	232	259	233
rect	258	233	259	234
rect	258	234	259	235
rect	258	235	259	236
rect	258	236	259	237
rect	258	237	259	238
rect	258	239	259	240
rect	258	240	259	241
rect	258	241	259	242
rect	258	242	259	243
rect	258	243	259	244
rect	258	244	259	245
rect	258	245	259	246
rect	258	246	259	247
rect	258	247	259	248
rect	258	248	259	249
rect	258	249	259	250
rect	258	250	259	251
rect	258	251	259	252
rect	259	0	260	1
rect	259	1	260	2
rect	259	2	260	3
rect	259	3	260	4
rect	259	4	260	5
rect	259	5	260	6
rect	259	6	260	7
rect	259	8	260	9
rect	259	9	260	10
rect	259	11	260	12
rect	259	12	260	13
rect	259	14	260	15
rect	259	15	260	16
rect	259	17	260	18
rect	259	18	260	19
rect	259	20	260	21
rect	259	21	260	22
rect	259	23	260	24
rect	259	24	260	25
rect	259	26	260	27
rect	259	27	260	28
rect	259	29	260	30
rect	259	30	260	31
rect	259	32	260	33
rect	259	33	260	34
rect	259	35	260	36
rect	259	36	260	37
rect	259	38	260	39
rect	259	39	260	40
rect	259	41	260	42
rect	259	42	260	43
rect	259	44	260	45
rect	259	45	260	46
rect	259	47	260	48
rect	259	48	260	49
rect	259	50	260	51
rect	259	51	260	52
rect	259	53	260	54
rect	259	54	260	55
rect	259	56	260	57
rect	259	57	260	58
rect	259	59	260	60
rect	259	60	260	61
rect	259	62	260	63
rect	259	63	260	64
rect	259	65	260	66
rect	259	66	260	67
rect	259	68	260	69
rect	259	69	260	70
rect	259	70	260	71
rect	259	71	260	72
rect	259	72	260	73
rect	259	73	260	74
rect	259	74	260	75
rect	259	75	260	76
rect	259	76	260	77
rect	259	77	260	78
rect	259	78	260	79
rect	259	80	260	81
rect	259	81	260	82
rect	259	83	260	84
rect	259	84	260	85
rect	259	86	260	87
rect	259	87	260	88
rect	259	89	260	90
rect	259	90	260	91
rect	259	91	260	92
rect	259	92	260	93
rect	259	93	260	94
rect	259	94	260	95
rect	259	95	260	96
rect	259	96	260	97
rect	259	97	260	98
rect	259	98	260	99
rect	259	99	260	100
rect	259	101	260	102
rect	259	102	260	103
rect	259	104	260	105
rect	259	105	260	106
rect	259	106	260	107
rect	259	107	260	108
rect	259	108	260	109
rect	259	110	260	111
rect	259	111	260	112
rect	259	112	260	113
rect	259	113	260	114
rect	259	114	260	115
rect	259	116	260	117
rect	259	117	260	118
rect	259	119	260	120
rect	259	120	260	121
rect	259	121	260	122
rect	259	122	260	123
rect	259	123	260	124
rect	259	125	260	126
rect	259	126	260	127
rect	259	128	260	129
rect	259	129	260	130
rect	259	130	260	131
rect	259	131	260	132
rect	259	132	260	133
rect	259	134	260	135
rect	259	135	260	136
rect	259	137	260	138
rect	259	138	260	139
rect	259	140	260	141
rect	259	141	260	142
rect	259	143	260	144
rect	259	144	260	145
rect	259	145	260	146
rect	259	146	260	147
rect	259	147	260	148
rect	259	149	260	150
rect	259	150	260	151
rect	259	152	260	153
rect	259	153	260	154
rect	259	154	260	155
rect	259	155	260	156
rect	259	156	260	157
rect	259	158	260	159
rect	259	159	260	160
rect	259	161	260	162
rect	259	162	260	163
rect	259	164	260	165
rect	259	165	260	166
rect	259	167	260	168
rect	259	168	260	169
rect	259	170	260	171
rect	259	171	260	172
rect	259	173	260	174
rect	259	174	260	175
rect	259	176	260	177
rect	259	177	260	178
rect	259	179	260	180
rect	259	180	260	181
rect	259	182	260	183
rect	259	183	260	184
rect	259	185	260	186
rect	259	186	260	187
rect	259	188	260	189
rect	259	189	260	190
rect	259	190	260	191
rect	259	191	260	192
rect	259	192	260	193
rect	259	194	260	195
rect	259	195	260	196
rect	259	197	260	198
rect	259	198	260	199
rect	259	200	260	201
rect	259	201	260	202
rect	259	203	260	204
rect	259	204	260	205
rect	259	206	260	207
rect	259	207	260	208
rect	259	209	260	210
rect	259	210	260	211
rect	259	212	260	213
rect	259	213	260	214
rect	259	214	260	215
rect	259	215	260	216
rect	259	216	260	217
rect	259	218	260	219
rect	259	219	260	220
rect	259	220	260	221
rect	259	221	260	222
rect	259	222	260	223
rect	259	224	260	225
rect	259	225	260	226
rect	259	226	260	227
rect	259	227	260	228
rect	259	228	260	229
rect	259	229	260	230
rect	259	230	260	231
rect	259	231	260	232
rect	259	232	260	233
rect	259	233	260	234
rect	259	234	260	235
rect	259	235	260	236
rect	259	236	260	237
rect	259	237	260	238
rect	259	239	260	240
rect	259	240	260	241
rect	259	241	260	242
rect	259	242	260	243
rect	259	243	260	244
rect	259	244	260	245
rect	259	245	260	246
rect	259	246	260	247
rect	259	247	260	248
rect	259	248	260	249
rect	259	249	260	250
rect	259	250	260	251
rect	259	251	260	252
rect	260	0	261	1
rect	260	1	261	2
rect	260	2	261	3
rect	260	3	261	4
rect	260	4	261	5
rect	260	5	261	6
rect	260	6	261	7
rect	260	8	261	9
rect	260	9	261	10
rect	260	11	261	12
rect	260	12	261	13
rect	260	14	261	15
rect	260	15	261	16
rect	260	17	261	18
rect	260	18	261	19
rect	260	20	261	21
rect	260	21	261	22
rect	260	23	261	24
rect	260	24	261	25
rect	260	26	261	27
rect	260	27	261	28
rect	260	29	261	30
rect	260	30	261	31
rect	260	32	261	33
rect	260	33	261	34
rect	260	35	261	36
rect	260	36	261	37
rect	260	38	261	39
rect	260	39	261	40
rect	260	41	261	42
rect	260	42	261	43
rect	260	44	261	45
rect	260	45	261	46
rect	260	47	261	48
rect	260	48	261	49
rect	260	50	261	51
rect	260	51	261	52
rect	260	53	261	54
rect	260	54	261	55
rect	260	56	261	57
rect	260	57	261	58
rect	260	59	261	60
rect	260	60	261	61
rect	260	62	261	63
rect	260	63	261	64
rect	260	65	261	66
rect	260	66	261	67
rect	260	68	261	69
rect	260	69	261	70
rect	260	70	261	71
rect	260	71	261	72
rect	260	72	261	73
rect	260	73	261	74
rect	260	74	261	75
rect	260	75	261	76
rect	260	76	261	77
rect	260	77	261	78
rect	260	78	261	79
rect	260	80	261	81
rect	260	81	261	82
rect	260	83	261	84
rect	260	84	261	85
rect	260	86	261	87
rect	260	87	261	88
rect	260	89	261	90
rect	260	90	261	91
rect	260	91	261	92
rect	260	92	261	93
rect	260	93	261	94
rect	260	94	261	95
rect	260	95	261	96
rect	260	96	261	97
rect	260	97	261	98
rect	260	98	261	99
rect	260	99	261	100
rect	260	101	261	102
rect	260	102	261	103
rect	260	104	261	105
rect	260	105	261	106
rect	260	106	261	107
rect	260	107	261	108
rect	260	108	261	109
rect	260	110	261	111
rect	260	111	261	112
rect	260	112	261	113
rect	260	113	261	114
rect	260	114	261	115
rect	260	116	261	117
rect	260	117	261	118
rect	260	119	261	120
rect	260	120	261	121
rect	260	121	261	122
rect	260	122	261	123
rect	260	123	261	124
rect	260	125	261	126
rect	260	126	261	127
rect	260	128	261	129
rect	260	129	261	130
rect	260	130	261	131
rect	260	131	261	132
rect	260	132	261	133
rect	260	134	261	135
rect	260	135	261	136
rect	260	137	261	138
rect	260	138	261	139
rect	260	140	261	141
rect	260	141	261	142
rect	260	143	261	144
rect	260	144	261	145
rect	260	145	261	146
rect	260	146	261	147
rect	260	147	261	148
rect	260	149	261	150
rect	260	150	261	151
rect	260	152	261	153
rect	260	153	261	154
rect	260	154	261	155
rect	260	155	261	156
rect	260	156	261	157
rect	260	158	261	159
rect	260	159	261	160
rect	260	161	261	162
rect	260	162	261	163
rect	260	164	261	165
rect	260	165	261	166
rect	260	167	261	168
rect	260	168	261	169
rect	260	170	261	171
rect	260	171	261	172
rect	260	173	261	174
rect	260	174	261	175
rect	260	176	261	177
rect	260	177	261	178
rect	260	179	261	180
rect	260	180	261	181
rect	260	182	261	183
rect	260	183	261	184
rect	260	185	261	186
rect	260	186	261	187
rect	260	188	261	189
rect	260	189	261	190
rect	260	190	261	191
rect	260	191	261	192
rect	260	192	261	193
rect	260	194	261	195
rect	260	195	261	196
rect	260	197	261	198
rect	260	198	261	199
rect	260	200	261	201
rect	260	201	261	202
rect	260	203	261	204
rect	260	204	261	205
rect	260	206	261	207
rect	260	207	261	208
rect	260	209	261	210
rect	260	210	261	211
rect	260	212	261	213
rect	260	213	261	214
rect	260	214	261	215
rect	260	215	261	216
rect	260	216	261	217
rect	260	218	261	219
rect	260	219	261	220
rect	260	220	261	221
rect	260	221	261	222
rect	260	222	261	223
rect	260	224	261	225
rect	260	225	261	226
rect	260	226	261	227
rect	260	227	261	228
rect	260	228	261	229
rect	260	229	261	230
rect	260	230	261	231
rect	260	231	261	232
rect	260	232	261	233
rect	260	233	261	234
rect	260	234	261	235
rect	260	235	261	236
rect	260	236	261	237
rect	260	237	261	238
rect	260	239	261	240
rect	260	240	261	241
rect	260	241	261	242
rect	260	242	261	243
rect	260	243	261	244
rect	260	244	261	245
rect	260	245	261	246
rect	260	246	261	247
rect	260	247	261	248
rect	260	248	261	249
rect	260	249	261	250
rect	260	250	261	251
rect	260	251	261	252
rect	261	0	262	1
rect	261	1	262	2
rect	261	2	262	3
rect	261	3	262	4
rect	261	4	262	5
rect	261	5	262	6
rect	261	6	262	7
rect	261	8	262	9
rect	261	9	262	10
rect	261	11	262	12
rect	261	12	262	13
rect	261	14	262	15
rect	261	15	262	16
rect	261	17	262	18
rect	261	18	262	19
rect	261	20	262	21
rect	261	21	262	22
rect	261	23	262	24
rect	261	24	262	25
rect	261	26	262	27
rect	261	27	262	28
rect	261	29	262	30
rect	261	30	262	31
rect	261	32	262	33
rect	261	33	262	34
rect	261	35	262	36
rect	261	36	262	37
rect	261	38	262	39
rect	261	39	262	40
rect	261	41	262	42
rect	261	42	262	43
rect	261	44	262	45
rect	261	45	262	46
rect	261	47	262	48
rect	261	48	262	49
rect	261	50	262	51
rect	261	51	262	52
rect	261	53	262	54
rect	261	54	262	55
rect	261	56	262	57
rect	261	57	262	58
rect	261	59	262	60
rect	261	60	262	61
rect	261	62	262	63
rect	261	63	262	64
rect	261	65	262	66
rect	261	66	262	67
rect	261	68	262	69
rect	261	69	262	70
rect	261	70	262	71
rect	261	71	262	72
rect	261	72	262	73
rect	261	73	262	74
rect	261	74	262	75
rect	261	75	262	76
rect	261	76	262	77
rect	261	77	262	78
rect	261	78	262	79
rect	261	80	262	81
rect	261	81	262	82
rect	261	83	262	84
rect	261	84	262	85
rect	261	86	262	87
rect	261	87	262	88
rect	261	89	262	90
rect	261	90	262	91
rect	261	91	262	92
rect	261	92	262	93
rect	261	93	262	94
rect	261	94	262	95
rect	261	95	262	96
rect	261	96	262	97
rect	261	97	262	98
rect	261	98	262	99
rect	261	99	262	100
rect	261	101	262	102
rect	261	102	262	103
rect	261	104	262	105
rect	261	105	262	106
rect	261	106	262	107
rect	261	107	262	108
rect	261	108	262	109
rect	261	110	262	111
rect	261	111	262	112
rect	261	112	262	113
rect	261	113	262	114
rect	261	114	262	115
rect	261	116	262	117
rect	261	117	262	118
rect	261	119	262	120
rect	261	120	262	121
rect	261	121	262	122
rect	261	122	262	123
rect	261	123	262	124
rect	261	125	262	126
rect	261	126	262	127
rect	261	128	262	129
rect	261	129	262	130
rect	261	130	262	131
rect	261	131	262	132
rect	261	132	262	133
rect	261	134	262	135
rect	261	135	262	136
rect	261	137	262	138
rect	261	138	262	139
rect	261	140	262	141
rect	261	141	262	142
rect	261	143	262	144
rect	261	144	262	145
rect	261	145	262	146
rect	261	146	262	147
rect	261	147	262	148
rect	261	149	262	150
rect	261	150	262	151
rect	261	152	262	153
rect	261	153	262	154
rect	261	154	262	155
rect	261	155	262	156
rect	261	156	262	157
rect	261	158	262	159
rect	261	159	262	160
rect	261	161	262	162
rect	261	162	262	163
rect	261	164	262	165
rect	261	165	262	166
rect	261	167	262	168
rect	261	168	262	169
rect	261	170	262	171
rect	261	171	262	172
rect	261	173	262	174
rect	261	174	262	175
rect	261	176	262	177
rect	261	177	262	178
rect	261	179	262	180
rect	261	180	262	181
rect	261	182	262	183
rect	261	183	262	184
rect	261	185	262	186
rect	261	186	262	187
rect	261	188	262	189
rect	261	189	262	190
rect	261	190	262	191
rect	261	191	262	192
rect	261	192	262	193
rect	261	194	262	195
rect	261	195	262	196
rect	261	197	262	198
rect	261	198	262	199
rect	261	200	262	201
rect	261	201	262	202
rect	261	203	262	204
rect	261	204	262	205
rect	261	206	262	207
rect	261	207	262	208
rect	261	209	262	210
rect	261	210	262	211
rect	261	212	262	213
rect	261	213	262	214
rect	261	214	262	215
rect	261	215	262	216
rect	261	216	262	217
rect	261	218	262	219
rect	261	219	262	220
rect	261	220	262	221
rect	261	221	262	222
rect	261	222	262	223
rect	261	224	262	225
rect	261	225	262	226
rect	261	226	262	227
rect	261	227	262	228
rect	261	228	262	229
rect	261	229	262	230
rect	261	230	262	231
rect	261	231	262	232
rect	261	232	262	233
rect	261	233	262	234
rect	261	234	262	235
rect	261	235	262	236
rect	261	236	262	237
rect	261	237	262	238
rect	261	239	262	240
rect	261	240	262	241
rect	261	241	262	242
rect	261	242	262	243
rect	261	243	262	244
rect	261	244	262	245
rect	261	245	262	246
rect	261	246	262	247
rect	261	247	262	248
rect	261	248	262	249
rect	261	249	262	250
rect	261	250	262	251
rect	261	251	262	252
rect	264	0	265	1
rect	264	1	265	2
rect	264	2	265	3
rect	264	3	265	4
rect	264	4	265	5
rect	264	5	265	6
rect	264	6	265	7
rect	264	8	265	9
rect	264	9	265	10
rect	264	11	265	12
rect	264	12	265	13
rect	264	14	265	15
rect	264	15	265	16
rect	264	17	265	18
rect	264	18	265	19
rect	264	20	265	21
rect	264	21	265	22
rect	264	23	265	24
rect	264	24	265	25
rect	264	26	265	27
rect	264	27	265	28
rect	264	29	265	30
rect	264	30	265	31
rect	264	32	265	33
rect	264	33	265	34
rect	264	35	265	36
rect	264	36	265	37
rect	264	38	265	39
rect	264	39	265	40
rect	264	41	265	42
rect	264	42	265	43
rect	264	44	265	45
rect	264	45	265	46
rect	264	47	265	48
rect	264	48	265	49
rect	264	50	265	51
rect	264	51	265	52
rect	264	53	265	54
rect	264	54	265	55
rect	264	56	265	57
rect	264	57	265	58
rect	264	59	265	60
rect	264	60	265	61
rect	264	62	265	63
rect	264	63	265	64
rect	264	65	265	66
rect	264	66	265	67
rect	264	67	265	68
rect	264	68	265	69
rect	264	69	265	70
rect	264	70	265	71
rect	264	71	265	72
rect	264	72	265	73
rect	264	73	265	74
rect	264	74	265	75
rect	264	75	265	76
rect	264	76	265	77
rect	264	77	265	78
rect	264	78	265	79
rect	264	80	265	81
rect	264	81	265	82
rect	264	83	265	84
rect	264	84	265	85
rect	264	86	265	87
rect	264	87	265	88
rect	264	89	265	90
rect	264	90	265	91
rect	264	91	265	92
rect	264	92	265	93
rect	264	93	265	94
rect	264	94	265	95
rect	264	95	265	96
rect	264	96	265	97
rect	264	97	265	98
rect	264	98	265	99
rect	264	99	265	100
rect	264	100	265	101
rect	264	101	265	102
rect	264	102	265	103
rect	264	104	265	105
rect	264	105	265	106
rect	264	106	265	107
rect	264	107	265	108
rect	264	108	265	109
rect	264	110	265	111
rect	264	111	265	112
rect	264	112	265	113
rect	264	113	265	114
rect	264	114	265	115
rect	264	116	265	117
rect	264	117	265	118
rect	264	119	265	120
rect	264	120	265	121
rect	264	121	265	122
rect	264	122	265	123
rect	264	123	265	124
rect	264	125	265	126
rect	264	126	265	127
rect	264	128	265	129
rect	264	129	265	130
rect	264	130	265	131
rect	264	131	265	132
rect	264	132	265	133
rect	264	134	265	135
rect	264	135	265	136
rect	264	137	265	138
rect	264	138	265	139
rect	264	140	265	141
rect	264	141	265	142
rect	264	143	265	144
rect	264	144	265	145
rect	264	145	265	146
rect	264	146	265	147
rect	264	147	265	148
rect	264	149	265	150
rect	264	150	265	151
rect	264	152	265	153
rect	264	153	265	154
rect	264	154	265	155
rect	264	155	265	156
rect	264	156	265	157
rect	264	158	265	159
rect	264	159	265	160
rect	264	161	265	162
rect	264	162	265	163
rect	264	164	265	165
rect	264	165	265	166
rect	264	167	265	168
rect	264	168	265	169
rect	264	170	265	171
rect	264	171	265	172
rect	264	173	265	174
rect	264	174	265	175
rect	264	176	265	177
rect	264	177	265	178
rect	264	179	265	180
rect	264	180	265	181
rect	264	182	265	183
rect	264	183	265	184
rect	264	185	265	186
rect	264	186	265	187
rect	264	188	265	189
rect	264	189	265	190
rect	264	190	265	191
rect	264	191	265	192
rect	264	192	265	193
rect	264	194	265	195
rect	264	195	265	196
rect	264	197	265	198
rect	264	198	265	199
rect	264	200	265	201
rect	264	201	265	202
rect	264	203	265	204
rect	264	204	265	205
rect	264	205	265	206
rect	264	206	265	207
rect	264	207	265	208
rect	264	208	265	209
rect	264	209	265	210
rect	264	210	265	211
rect	264	212	265	213
rect	264	213	265	214
rect	264	214	265	215
rect	264	215	265	216
rect	264	216	265	217
rect	264	218	265	219
rect	264	219	265	220
rect	264	220	265	221
rect	264	221	265	222
rect	264	222	265	223
rect	264	223	265	224
rect	264	224	265	225
rect	264	225	265	226
rect	264	226	265	227
rect	264	227	265	228
rect	264	228	265	229
rect	264	229	265	230
rect	264	230	265	231
rect	264	231	265	232
rect	264	232	265	233
rect	264	233	265	234
rect	264	234	265	235
rect	264	235	265	236
rect	264	236	265	237
rect	264	237	265	238
rect	264	239	265	240
rect	264	240	265	241
rect	264	241	265	242
rect	264	242	265	243
rect	264	243	265	244
rect	264	244	265	245
rect	264	245	265	246
rect	264	246	265	247
rect	264	247	265	248
rect	264	248	265	249
rect	264	249	265	250
rect	264	250	265	251
rect	264	251	265	252
rect	266	0	267	1
rect	266	1	267	2
rect	266	2	267	3
rect	266	3	267	4
rect	266	4	267	5
rect	266	5	267	6
rect	266	6	267	7
rect	266	8	267	9
rect	266	9	267	10
rect	266	11	267	12
rect	266	12	267	13
rect	266	14	267	15
rect	266	15	267	16
rect	266	17	267	18
rect	266	18	267	19
rect	266	20	267	21
rect	266	21	267	22
rect	266	23	267	24
rect	266	24	267	25
rect	266	26	267	27
rect	266	27	267	28
rect	266	29	267	30
rect	266	30	267	31
rect	266	32	267	33
rect	266	33	267	34
rect	266	35	267	36
rect	266	36	267	37
rect	266	38	267	39
rect	266	39	267	40
rect	266	41	267	42
rect	266	42	267	43
rect	266	44	267	45
rect	266	45	267	46
rect	266	47	267	48
rect	266	48	267	49
rect	266	50	267	51
rect	266	51	267	52
rect	266	53	267	54
rect	266	54	267	55
rect	266	56	267	57
rect	266	57	267	58
rect	266	59	267	60
rect	266	60	267	61
rect	266	62	267	63
rect	266	63	267	64
rect	266	65	267	66
rect	266	66	267	67
rect	266	67	267	68
rect	266	68	267	69
rect	266	69	267	70
rect	266	70	267	71
rect	266	71	267	72
rect	266	72	267	73
rect	266	73	267	74
rect	266	74	267	75
rect	266	75	267	76
rect	266	76	267	77
rect	266	77	267	78
rect	266	78	267	79
rect	266	80	267	81
rect	266	81	267	82
rect	266	83	267	84
rect	266	84	267	85
rect	266	86	267	87
rect	266	87	267	88
rect	266	89	267	90
rect	266	90	267	91
rect	266	91	267	92
rect	266	92	267	93
rect	266	93	267	94
rect	266	94	267	95
rect	266	95	267	96
rect	266	96	267	97
rect	266	97	267	98
rect	266	98	267	99
rect	266	99	267	100
rect	266	100	267	101
rect	266	101	267	102
rect	266	102	267	103
rect	266	104	267	105
rect	266	105	267	106
rect	266	106	267	107
rect	266	107	267	108
rect	266	108	267	109
rect	266	110	267	111
rect	266	111	267	112
rect	266	112	267	113
rect	266	113	267	114
rect	266	114	267	115
rect	266	116	267	117
rect	266	117	267	118
rect	266	119	267	120
rect	266	120	267	121
rect	266	121	267	122
rect	266	122	267	123
rect	266	123	267	124
rect	266	125	267	126
rect	266	126	267	127
rect	266	128	267	129
rect	266	129	267	130
rect	266	130	267	131
rect	266	131	267	132
rect	266	132	267	133
rect	266	134	267	135
rect	266	135	267	136
rect	266	137	267	138
rect	266	138	267	139
rect	266	140	267	141
rect	266	141	267	142
rect	266	143	267	144
rect	266	144	267	145
rect	266	145	267	146
rect	266	146	267	147
rect	266	147	267	148
rect	266	149	267	150
rect	266	150	267	151
rect	266	152	267	153
rect	266	153	267	154
rect	266	154	267	155
rect	266	155	267	156
rect	266	156	267	157
rect	266	158	267	159
rect	266	159	267	160
rect	266	161	267	162
rect	266	162	267	163
rect	266	164	267	165
rect	266	165	267	166
rect	266	167	267	168
rect	266	168	267	169
rect	266	170	267	171
rect	266	171	267	172
rect	266	173	267	174
rect	266	174	267	175
rect	266	176	267	177
rect	266	177	267	178
rect	266	179	267	180
rect	266	180	267	181
rect	266	182	267	183
rect	266	183	267	184
rect	266	185	267	186
rect	266	186	267	187
rect	266	188	267	189
rect	266	189	267	190
rect	266	190	267	191
rect	266	191	267	192
rect	266	192	267	193
rect	266	194	267	195
rect	266	195	267	196
rect	266	197	267	198
rect	266	198	267	199
rect	266	200	267	201
rect	266	201	267	202
rect	266	203	267	204
rect	266	204	267	205
rect	266	205	267	206
rect	266	206	267	207
rect	266	207	267	208
rect	266	208	267	209
rect	266	209	267	210
rect	266	210	267	211
rect	266	212	267	213
rect	266	213	267	214
rect	266	214	267	215
rect	266	215	267	216
rect	266	216	267	217
rect	266	218	267	219
rect	266	219	267	220
rect	266	220	267	221
rect	266	221	267	222
rect	266	222	267	223
rect	266	223	267	224
rect	266	224	267	225
rect	266	225	267	226
rect	266	226	267	227
rect	266	227	267	228
rect	266	228	267	229
rect	266	229	267	230
rect	266	230	267	231
rect	266	231	267	232
rect	266	232	267	233
rect	266	233	267	234
rect	266	234	267	235
rect	266	235	267	236
rect	266	236	267	237
rect	266	237	267	238
rect	266	239	267	240
rect	267	0	268	1
rect	267	1	268	2
rect	267	2	268	3
rect	267	3	268	4
rect	267	4	268	5
rect	267	5	268	6
rect	267	6	268	7
rect	267	8	268	9
rect	267	9	268	10
rect	267	11	268	12
rect	267	12	268	13
rect	267	14	268	15
rect	267	15	268	16
rect	267	17	268	18
rect	267	18	268	19
rect	267	20	268	21
rect	267	21	268	22
rect	267	23	268	24
rect	267	24	268	25
rect	267	26	268	27
rect	267	27	268	28
rect	267	29	268	30
rect	267	30	268	31
rect	267	32	268	33
rect	267	33	268	34
rect	267	35	268	36
rect	267	36	268	37
rect	267	38	268	39
rect	267	39	268	40
rect	267	41	268	42
rect	267	42	268	43
rect	267	44	268	45
rect	267	45	268	46
rect	267	47	268	48
rect	267	48	268	49
rect	267	50	268	51
rect	267	51	268	52
rect	267	53	268	54
rect	267	54	268	55
rect	267	56	268	57
rect	267	57	268	58
rect	267	59	268	60
rect	267	60	268	61
rect	267	62	268	63
rect	267	63	268	64
rect	267	65	268	66
rect	267	66	268	67
rect	267	67	268	68
rect	267	68	268	69
rect	267	69	268	70
rect	267	70	268	71
rect	267	71	268	72
rect	267	72	268	73
rect	267	73	268	74
rect	267	74	268	75
rect	267	75	268	76
rect	267	76	268	77
rect	267	77	268	78
rect	267	78	268	79
rect	267	80	268	81
rect	267	81	268	82
rect	267	83	268	84
rect	267	84	268	85
rect	267	86	268	87
rect	267	87	268	88
rect	267	89	268	90
rect	267	90	268	91
rect	267	91	268	92
rect	267	92	268	93
rect	267	93	268	94
rect	267	94	268	95
rect	267	95	268	96
rect	267	96	268	97
rect	267	97	268	98
rect	267	98	268	99
rect	267	99	268	100
rect	267	100	268	101
rect	267	101	268	102
rect	267	102	268	103
rect	267	104	268	105
rect	267	105	268	106
rect	267	106	268	107
rect	267	107	268	108
rect	267	108	268	109
rect	267	110	268	111
rect	267	111	268	112
rect	267	112	268	113
rect	267	113	268	114
rect	267	114	268	115
rect	267	116	268	117
rect	267	117	268	118
rect	267	119	268	120
rect	267	120	268	121
rect	267	121	268	122
rect	267	122	268	123
rect	267	123	268	124
rect	267	125	268	126
rect	267	126	268	127
rect	267	128	268	129
rect	267	129	268	130
rect	267	130	268	131
rect	267	131	268	132
rect	267	132	268	133
rect	267	134	268	135
rect	267	135	268	136
rect	267	137	268	138
rect	267	138	268	139
rect	267	140	268	141
rect	267	141	268	142
rect	267	143	268	144
rect	267	144	268	145
rect	267	145	268	146
rect	267	146	268	147
rect	267	147	268	148
rect	267	149	268	150
rect	267	150	268	151
rect	267	152	268	153
rect	267	153	268	154
rect	267	154	268	155
rect	267	155	268	156
rect	267	156	268	157
rect	267	158	268	159
rect	267	159	268	160
rect	267	161	268	162
rect	267	162	268	163
rect	267	164	268	165
rect	267	165	268	166
rect	267	167	268	168
rect	267	168	268	169
rect	267	170	268	171
rect	267	171	268	172
rect	267	173	268	174
rect	267	174	268	175
rect	267	176	268	177
rect	267	177	268	178
rect	267	179	268	180
rect	267	180	268	181
rect	267	182	268	183
rect	267	183	268	184
rect	267	185	268	186
rect	267	186	268	187
rect	267	188	268	189
rect	267	189	268	190
rect	267	190	268	191
rect	267	191	268	192
rect	267	192	268	193
rect	267	194	268	195
rect	267	195	268	196
rect	267	197	268	198
rect	267	198	268	199
rect	267	200	268	201
rect	267	201	268	202
rect	267	203	268	204
rect	267	204	268	205
rect	267	205	268	206
rect	267	206	268	207
rect	267	207	268	208
rect	267	208	268	209
rect	267	209	268	210
rect	267	210	268	211
rect	267	212	268	213
rect	267	213	268	214
rect	267	214	268	215
rect	267	215	268	216
rect	267	216	268	217
rect	267	218	268	219
rect	267	219	268	220
rect	267	220	268	221
rect	267	221	268	222
rect	267	222	268	223
rect	267	223	268	224
rect	267	224	268	225
rect	267	225	268	226
rect	267	226	268	227
rect	267	227	268	228
rect	267	228	268	229
rect	267	229	268	230
rect	267	230	268	231
rect	267	231	268	232
rect	267	232	268	233
rect	267	233	268	234
rect	267	234	268	235
rect	267	235	268	236
rect	267	236	268	237
rect	267	237	268	238
rect	267	239	268	240
rect	268	0	269	1
rect	268	1	269	2
rect	268	2	269	3
rect	268	3	269	4
rect	268	4	269	5
rect	268	5	269	6
rect	268	6	269	7
rect	268	8	269	9
rect	268	9	269	10
rect	268	11	269	12
rect	268	12	269	13
rect	268	14	269	15
rect	268	15	269	16
rect	268	17	269	18
rect	268	18	269	19
rect	268	20	269	21
rect	268	21	269	22
rect	268	23	269	24
rect	268	24	269	25
rect	268	26	269	27
rect	268	27	269	28
rect	268	29	269	30
rect	268	30	269	31
rect	268	32	269	33
rect	268	33	269	34
rect	268	35	269	36
rect	268	36	269	37
rect	268	38	269	39
rect	268	39	269	40
rect	268	41	269	42
rect	268	42	269	43
rect	268	44	269	45
rect	268	45	269	46
rect	268	47	269	48
rect	268	48	269	49
rect	268	50	269	51
rect	268	51	269	52
rect	268	53	269	54
rect	268	54	269	55
rect	268	56	269	57
rect	268	57	269	58
rect	268	59	269	60
rect	268	60	269	61
rect	268	62	269	63
rect	268	63	269	64
rect	268	65	269	66
rect	268	66	269	67
rect	268	67	269	68
rect	268	68	269	69
rect	268	69	269	70
rect	268	70	269	71
rect	268	71	269	72
rect	268	72	269	73
rect	268	73	269	74
rect	268	74	269	75
rect	268	75	269	76
rect	268	76	269	77
rect	268	77	269	78
rect	268	78	269	79
rect	268	80	269	81
rect	268	81	269	82
rect	268	83	269	84
rect	268	84	269	85
rect	268	86	269	87
rect	268	87	269	88
rect	268	89	269	90
rect	268	90	269	91
rect	268	91	269	92
rect	268	92	269	93
rect	268	93	269	94
rect	268	94	269	95
rect	268	95	269	96
rect	268	96	269	97
rect	268	97	269	98
rect	268	98	269	99
rect	268	99	269	100
rect	268	100	269	101
rect	268	101	269	102
rect	268	102	269	103
rect	268	104	269	105
rect	268	105	269	106
rect	268	106	269	107
rect	268	107	269	108
rect	268	108	269	109
rect	268	110	269	111
rect	268	111	269	112
rect	268	112	269	113
rect	268	113	269	114
rect	268	114	269	115
rect	268	116	269	117
rect	268	117	269	118
rect	268	119	269	120
rect	268	120	269	121
rect	268	121	269	122
rect	268	122	269	123
rect	268	123	269	124
rect	268	125	269	126
rect	268	126	269	127
rect	268	128	269	129
rect	268	129	269	130
rect	268	130	269	131
rect	268	131	269	132
rect	268	132	269	133
rect	268	134	269	135
rect	268	135	269	136
rect	268	137	269	138
rect	268	138	269	139
rect	268	140	269	141
rect	268	141	269	142
rect	268	143	269	144
rect	268	144	269	145
rect	268	145	269	146
rect	268	146	269	147
rect	268	147	269	148
rect	268	149	269	150
rect	268	150	269	151
rect	268	152	269	153
rect	268	153	269	154
rect	268	154	269	155
rect	268	155	269	156
rect	268	156	269	157
rect	268	158	269	159
rect	268	159	269	160
rect	268	161	269	162
rect	268	162	269	163
rect	268	164	269	165
rect	268	165	269	166
rect	268	167	269	168
rect	268	168	269	169
rect	268	170	269	171
rect	268	171	269	172
rect	268	173	269	174
rect	268	174	269	175
rect	268	176	269	177
rect	268	177	269	178
rect	268	179	269	180
rect	268	180	269	181
rect	268	182	269	183
rect	268	183	269	184
rect	268	185	269	186
rect	268	186	269	187
rect	268	188	269	189
rect	268	189	269	190
rect	268	190	269	191
rect	268	191	269	192
rect	268	192	269	193
rect	268	194	269	195
rect	268	195	269	196
rect	268	197	269	198
rect	268	198	269	199
rect	268	200	269	201
rect	268	201	269	202
rect	268	203	269	204
rect	268	204	269	205
rect	268	205	269	206
rect	268	206	269	207
rect	268	207	269	208
rect	268	208	269	209
rect	268	209	269	210
rect	268	210	269	211
rect	268	212	269	213
rect	268	213	269	214
rect	268	214	269	215
rect	268	215	269	216
rect	268	216	269	217
rect	268	218	269	219
rect	268	219	269	220
rect	268	220	269	221
rect	268	221	269	222
rect	268	222	269	223
rect	268	223	269	224
rect	268	224	269	225
rect	268	225	269	226
rect	268	226	269	227
rect	268	227	269	228
rect	268	228	269	229
rect	268	229	269	230
rect	268	230	269	231
rect	268	231	269	232
rect	268	232	269	233
rect	268	233	269	234
rect	268	234	269	235
rect	268	235	269	236
rect	268	236	269	237
rect	268	237	269	238
rect	268	239	269	240
rect	269	0	270	1
rect	269	1	270	2
rect	269	2	270	3
rect	269	3	270	4
rect	269	4	270	5
rect	269	5	270	6
rect	269	6	270	7
rect	269	8	270	9
rect	269	9	270	10
rect	269	11	270	12
rect	269	12	270	13
rect	269	14	270	15
rect	269	15	270	16
rect	269	17	270	18
rect	269	18	270	19
rect	269	20	270	21
rect	269	21	270	22
rect	269	23	270	24
rect	269	24	270	25
rect	269	26	270	27
rect	269	27	270	28
rect	269	29	270	30
rect	269	30	270	31
rect	269	32	270	33
rect	269	33	270	34
rect	269	35	270	36
rect	269	36	270	37
rect	269	38	270	39
rect	269	39	270	40
rect	269	41	270	42
rect	269	42	270	43
rect	269	44	270	45
rect	269	45	270	46
rect	269	47	270	48
rect	269	48	270	49
rect	269	50	270	51
rect	269	51	270	52
rect	269	53	270	54
rect	269	54	270	55
rect	269	56	270	57
rect	269	57	270	58
rect	269	59	270	60
rect	269	60	270	61
rect	269	62	270	63
rect	269	63	270	64
rect	269	65	270	66
rect	269	66	270	67
rect	269	67	270	68
rect	269	68	270	69
rect	269	69	270	70
rect	269	70	270	71
rect	269	71	270	72
rect	269	72	270	73
rect	269	73	270	74
rect	269	74	270	75
rect	269	75	270	76
rect	269	76	270	77
rect	269	77	270	78
rect	269	78	270	79
rect	269	80	270	81
rect	269	81	270	82
rect	269	83	270	84
rect	269	84	270	85
rect	269	86	270	87
rect	269	87	270	88
rect	269	89	270	90
rect	269	90	270	91
rect	269	91	270	92
rect	269	92	270	93
rect	269	93	270	94
rect	269	94	270	95
rect	269	95	270	96
rect	269	96	270	97
rect	269	97	270	98
rect	269	98	270	99
rect	269	99	270	100
rect	269	100	270	101
rect	269	101	270	102
rect	269	102	270	103
rect	269	104	270	105
rect	269	105	270	106
rect	269	106	270	107
rect	269	107	270	108
rect	269	108	270	109
rect	269	110	270	111
rect	269	111	270	112
rect	269	112	270	113
rect	269	113	270	114
rect	269	114	270	115
rect	269	116	270	117
rect	269	117	270	118
rect	269	119	270	120
rect	269	120	270	121
rect	269	121	270	122
rect	269	122	270	123
rect	269	123	270	124
rect	269	125	270	126
rect	269	126	270	127
rect	269	128	270	129
rect	269	129	270	130
rect	269	130	270	131
rect	269	131	270	132
rect	269	132	270	133
rect	269	134	270	135
rect	269	135	270	136
rect	269	137	270	138
rect	269	138	270	139
rect	269	140	270	141
rect	269	141	270	142
rect	269	143	270	144
rect	269	144	270	145
rect	269	145	270	146
rect	269	146	270	147
rect	269	147	270	148
rect	269	149	270	150
rect	269	150	270	151
rect	269	152	270	153
rect	269	153	270	154
rect	269	154	270	155
rect	269	155	270	156
rect	269	156	270	157
rect	269	158	270	159
rect	269	159	270	160
rect	269	161	270	162
rect	269	162	270	163
rect	269	164	270	165
rect	269	165	270	166
rect	269	167	270	168
rect	269	168	270	169
rect	269	170	270	171
rect	269	171	270	172
rect	269	173	270	174
rect	269	174	270	175
rect	269	176	270	177
rect	269	177	270	178
rect	269	179	270	180
rect	269	180	270	181
rect	269	182	270	183
rect	269	183	270	184
rect	269	185	270	186
rect	269	186	270	187
rect	269	188	270	189
rect	269	189	270	190
rect	269	190	270	191
rect	269	191	270	192
rect	269	192	270	193
rect	269	194	270	195
rect	269	195	270	196
rect	269	197	270	198
rect	269	198	270	199
rect	269	200	270	201
rect	269	201	270	202
rect	269	203	270	204
rect	269	204	270	205
rect	269	205	270	206
rect	269	206	270	207
rect	269	207	270	208
rect	269	208	270	209
rect	269	209	270	210
rect	269	210	270	211
rect	269	212	270	213
rect	269	213	270	214
rect	269	214	270	215
rect	269	215	270	216
rect	269	216	270	217
rect	269	218	270	219
rect	269	219	270	220
rect	269	220	270	221
rect	269	221	270	222
rect	269	222	270	223
rect	269	223	270	224
rect	269	224	270	225
rect	269	225	270	226
rect	269	226	270	227
rect	269	227	270	228
rect	269	228	270	229
rect	269	229	270	230
rect	269	230	270	231
rect	269	231	270	232
rect	269	232	270	233
rect	269	233	270	234
rect	269	234	270	235
rect	269	235	270	236
rect	269	236	270	237
rect	269	237	270	238
rect	269	239	270	240
rect	270	0	271	1
rect	270	1	271	2
rect	270	2	271	3
rect	270	3	271	4
rect	270	4	271	5
rect	270	5	271	6
rect	270	6	271	7
rect	270	8	271	9
rect	270	9	271	10
rect	270	11	271	12
rect	270	12	271	13
rect	270	14	271	15
rect	270	15	271	16
rect	270	17	271	18
rect	270	18	271	19
rect	270	20	271	21
rect	270	21	271	22
rect	270	23	271	24
rect	270	24	271	25
rect	270	26	271	27
rect	270	27	271	28
rect	270	29	271	30
rect	270	30	271	31
rect	270	32	271	33
rect	270	33	271	34
rect	270	35	271	36
rect	270	36	271	37
rect	270	38	271	39
rect	270	39	271	40
rect	270	41	271	42
rect	270	42	271	43
rect	270	44	271	45
rect	270	45	271	46
rect	270	47	271	48
rect	270	48	271	49
rect	270	50	271	51
rect	270	51	271	52
rect	270	52	271	53
rect	270	53	271	54
rect	270	54	271	55
rect	270	56	271	57
rect	270	57	271	58
rect	270	59	271	60
rect	270	60	271	61
rect	270	62	271	63
rect	270	63	271	64
rect	270	65	271	66
rect	270	66	271	67
rect	270	67	271	68
rect	270	68	271	69
rect	270	69	271	70
rect	270	70	271	71
rect	270	71	271	72
rect	270	72	271	73
rect	270	73	271	74
rect	270	74	271	75
rect	270	75	271	76
rect	270	76	271	77
rect	270	77	271	78
rect	270	78	271	79
rect	270	80	271	81
rect	270	81	271	82
rect	270	83	271	84
rect	270	84	271	85
rect	270	86	271	87
rect	270	87	271	88
rect	270	89	271	90
rect	270	90	271	91
rect	270	91	271	92
rect	270	92	271	93
rect	270	93	271	94
rect	270	94	271	95
rect	270	95	271	96
rect	270	96	271	97
rect	270	97	271	98
rect	270	98	271	99
rect	270	99	271	100
rect	270	100	271	101
rect	270	101	271	102
rect	270	102	271	103
rect	270	104	271	105
rect	270	105	271	106
rect	270	106	271	107
rect	270	107	271	108
rect	270	108	271	109
rect	270	110	271	111
rect	270	111	271	112
rect	270	112	271	113
rect	270	113	271	114
rect	270	114	271	115
rect	270	116	271	117
rect	270	117	271	118
rect	270	119	271	120
rect	270	120	271	121
rect	270	121	271	122
rect	270	122	271	123
rect	270	123	271	124
rect	270	125	271	126
rect	270	126	271	127
rect	270	128	271	129
rect	270	129	271	130
rect	270	130	271	131
rect	270	131	271	132
rect	270	132	271	133
rect	270	134	271	135
rect	270	135	271	136
rect	270	137	271	138
rect	270	138	271	139
rect	270	140	271	141
rect	270	141	271	142
rect	270	143	271	144
rect	270	144	271	145
rect	270	145	271	146
rect	270	146	271	147
rect	270	147	271	148
rect	270	149	271	150
rect	270	150	271	151
rect	270	152	271	153
rect	270	153	271	154
rect	270	154	271	155
rect	270	155	271	156
rect	270	156	271	157
rect	270	158	271	159
rect	270	159	271	160
rect	270	161	271	162
rect	270	162	271	163
rect	270	164	271	165
rect	270	165	271	166
rect	270	167	271	168
rect	270	168	271	169
rect	270	170	271	171
rect	270	171	271	172
rect	270	173	271	174
rect	270	174	271	175
rect	270	176	271	177
rect	270	177	271	178
rect	270	179	271	180
rect	270	180	271	181
rect	270	182	271	183
rect	270	183	271	184
rect	270	185	271	186
rect	270	186	271	187
rect	270	188	271	189
rect	270	189	271	190
rect	270	190	271	191
rect	270	191	271	192
rect	270	192	271	193
rect	270	193	271	194
rect	270	194	271	195
rect	270	195	271	196
rect	270	197	271	198
rect	270	198	271	199
rect	270	200	271	201
rect	270	201	271	202
rect	270	203	271	204
rect	270	204	271	205
rect	270	205	271	206
rect	270	206	271	207
rect	270	207	271	208
rect	270	208	271	209
rect	270	209	271	210
rect	270	210	271	211
rect	270	211	271	212
rect	270	212	271	213
rect	270	213	271	214
rect	270	214	271	215
rect	270	215	271	216
rect	270	216	271	217
rect	270	218	271	219
rect	270	219	271	220
rect	270	220	271	221
rect	270	221	271	222
rect	270	222	271	223
rect	270	223	271	224
rect	270	224	271	225
rect	270	225	271	226
rect	270	226	271	227
rect	270	227	271	228
rect	270	228	271	229
rect	270	229	271	230
rect	270	230	271	231
rect	270	231	271	232
rect	270	232	271	233
rect	270	233	271	234
rect	270	234	271	235
rect	270	235	271	236
rect	270	236	271	237
rect	270	237	271	238
rect	270	239	271	240
rect	275	0	276	1
rect	275	1	276	2
rect	275	2	276	3
rect	275	3	276	4
rect	275	4	276	5
rect	275	5	276	6
rect	275	6	276	7
rect	275	8	276	9
rect	275	9	276	10
rect	275	11	276	12
rect	275	12	276	13
rect	275	14	276	15
rect	275	15	276	16
rect	275	17	276	18
rect	275	18	276	19
rect	275	20	276	21
rect	275	21	276	22
rect	275	23	276	24
rect	275	24	276	25
rect	275	26	276	27
rect	275	27	276	28
rect	275	29	276	30
rect	275	30	276	31
rect	275	32	276	33
rect	275	33	276	34
rect	275	35	276	36
rect	275	36	276	37
rect	275	38	276	39
rect	275	39	276	40
rect	275	41	276	42
rect	275	42	276	43
rect	275	44	276	45
rect	275	45	276	46
rect	275	47	276	48
rect	275	48	276	49
rect	275	50	276	51
rect	275	51	276	52
rect	275	52	276	53
rect	275	53	276	54
rect	275	54	276	55
rect	275	56	276	57
rect	275	57	276	58
rect	275	58	276	59
rect	275	59	276	60
rect	275	60	276	61
rect	275	62	276	63
rect	275	63	276	64
rect	275	65	276	66
rect	275	66	276	67
rect	275	67	276	68
rect	275	68	276	69
rect	275	69	276	70
rect	275	70	276	71
rect	275	71	276	72
rect	275	72	276	73
rect	275	73	276	74
rect	275	74	276	75
rect	275	75	276	76
rect	275	76	276	77
rect	275	77	276	78
rect	275	78	276	79
rect	275	80	276	81
rect	275	81	276	82
rect	275	83	276	84
rect	275	84	276	85
rect	275	86	276	87
rect	275	87	276	88
rect	275	89	276	90
rect	275	90	276	91
rect	275	91	276	92
rect	275	92	276	93
rect	275	93	276	94
rect	275	94	276	95
rect	275	95	276	96
rect	275	96	276	97
rect	275	97	276	98
rect	275	98	276	99
rect	275	99	276	100
rect	275	100	276	101
rect	275	101	276	102
rect	275	102	276	103
rect	275	103	276	104
rect	275	104	276	105
rect	275	105	276	106
rect	275	106	276	107
rect	275	107	276	108
rect	275	108	276	109
rect	275	110	276	111
rect	275	111	276	112
rect	275	112	276	113
rect	275	113	276	114
rect	275	114	276	115
rect	275	116	276	117
rect	275	117	276	118
rect	275	119	276	120
rect	275	120	276	121
rect	275	121	276	122
rect	275	122	276	123
rect	275	123	276	124
rect	275	125	276	126
rect	275	126	276	127
rect	275	127	276	128
rect	275	128	276	129
rect	275	129	276	130
rect	275	130	276	131
rect	275	131	276	132
rect	275	132	276	133
rect	275	134	276	135
rect	275	135	276	136
rect	275	137	276	138
rect	275	138	276	139
rect	275	140	276	141
rect	275	141	276	142
rect	275	142	276	143
rect	275	143	276	144
rect	275	144	276	145
rect	275	145	276	146
rect	275	146	276	147
rect	275	147	276	148
rect	275	149	276	150
rect	275	150	276	151
rect	275	152	276	153
rect	275	153	276	154
rect	275	154	276	155
rect	275	155	276	156
rect	275	156	276	157
rect	275	158	276	159
rect	275	159	276	160
rect	275	161	276	162
rect	275	162	276	163
rect	275	164	276	165
rect	275	165	276	166
rect	275	167	276	168
rect	275	168	276	169
rect	275	170	276	171
rect	275	171	276	172
rect	275	173	276	174
rect	275	174	276	175
rect	275	176	276	177
rect	275	177	276	178
rect	275	179	276	180
rect	275	180	276	181
rect	275	181	276	182
rect	275	182	276	183
rect	275	183	276	184
rect	275	185	276	186
rect	275	186	276	187
rect	275	188	276	189
rect	275	189	276	190
rect	275	190	276	191
rect	275	191	276	192
rect	275	192	276	193
rect	275	193	276	194
rect	275	194	276	195
rect	275	195	276	196
rect	275	197	276	198
rect	275	198	276	199
rect	275	199	276	200
rect	275	200	276	201
rect	275	201	276	202
rect	275	202	276	203
rect	275	203	276	204
rect	275	204	276	205
rect	275	205	276	206
rect	275	206	276	207
rect	275	207	276	208
rect	275	208	276	209
rect	275	209	276	210
rect	275	210	276	211
rect	275	211	276	212
rect	275	212	276	213
rect	275	213	276	214
rect	275	214	276	215
rect	275	215	276	216
rect	275	216	276	217
rect	275	218	276	219
rect	275	219	276	220
rect	275	220	276	221
rect	275	221	276	222
rect	275	222	276	223
rect	275	223	276	224
rect	275	224	276	225
rect	275	225	276	226
rect	275	226	276	227
rect	275	227	276	228
rect	275	228	276	229
rect	275	229	276	230
rect	275	230	276	231
rect	275	231	276	232
rect	275	232	276	233
rect	275	233	276	234
rect	275	234	276	235
rect	275	235	276	236
rect	275	236	276	237
rect	275	237	276	238
rect	275	238	276	239
rect	275	239	276	240
rect	277	0	278	1
rect	277	1	278	2
rect	277	2	278	3
rect	277	3	278	4
rect	277	4	278	5
rect	277	5	278	6
rect	277	6	278	7
rect	277	8	278	9
rect	277	9	278	10
rect	277	11	278	12
rect	277	12	278	13
rect	277	14	278	15
rect	277	15	278	16
rect	277	17	278	18
rect	277	18	278	19
rect	277	20	278	21
rect	277	21	278	22
rect	277	23	278	24
rect	277	24	278	25
rect	277	26	278	27
rect	277	27	278	28
rect	277	29	278	30
rect	277	30	278	31
rect	277	32	278	33
rect	277	33	278	34
rect	277	35	278	36
rect	277	36	278	37
rect	277	38	278	39
rect	277	39	278	40
rect	277	41	278	42
rect	277	42	278	43
rect	277	44	278	45
rect	277	45	278	46
rect	277	47	278	48
rect	277	48	278	49
rect	277	50	278	51
rect	277	51	278	52
rect	277	52	278	53
rect	277	53	278	54
rect	277	54	278	55
rect	277	56	278	57
rect	277	57	278	58
rect	277	58	278	59
rect	277	59	278	60
rect	277	60	278	61
rect	277	62	278	63
rect	277	63	278	64
rect	277	65	278	66
rect	277	66	278	67
rect	277	67	278	68
rect	277	68	278	69
rect	277	69	278	70
rect	277	70	278	71
rect	277	71	278	72
rect	277	72	278	73
rect	277	73	278	74
rect	277	74	278	75
rect	277	75	278	76
rect	277	76	278	77
rect	277	77	278	78
rect	277	78	278	79
rect	277	80	278	81
rect	277	81	278	82
rect	277	83	278	84
rect	277	84	278	85
rect	277	86	278	87
rect	277	87	278	88
rect	277	89	278	90
rect	277	90	278	91
rect	277	91	278	92
rect	277	92	278	93
rect	277	93	278	94
rect	277	94	278	95
rect	277	95	278	96
rect	277	96	278	97
rect	277	97	278	98
rect	277	98	278	99
rect	277	99	278	100
rect	277	100	278	101
rect	277	101	278	102
rect	277	102	278	103
rect	277	103	278	104
rect	277	104	278	105
rect	277	105	278	106
rect	277	106	278	107
rect	277	107	278	108
rect	277	108	278	109
rect	277	110	278	111
rect	277	111	278	112
rect	277	112	278	113
rect	277	113	278	114
rect	277	114	278	115
rect	277	116	278	117
rect	277	117	278	118
rect	277	119	278	120
rect	277	120	278	121
rect	277	121	278	122
rect	277	122	278	123
rect	277	123	278	124
rect	277	125	278	126
rect	277	126	278	127
rect	277	127	278	128
rect	277	128	278	129
rect	277	129	278	130
rect	277	130	278	131
rect	277	131	278	132
rect	277	132	278	133
rect	277	134	278	135
rect	277	135	278	136
rect	277	137	278	138
rect	277	138	278	139
rect	277	140	278	141
rect	277	141	278	142
rect	277	142	278	143
rect	277	143	278	144
rect	277	144	278	145
rect	277	145	278	146
rect	277	146	278	147
rect	277	147	278	148
rect	277	149	278	150
rect	277	150	278	151
rect	277	152	278	153
rect	277	153	278	154
rect	277	154	278	155
rect	277	155	278	156
rect	277	156	278	157
rect	277	158	278	159
rect	277	159	278	160
rect	277	161	278	162
rect	277	162	278	163
rect	277	164	278	165
rect	277	165	278	166
rect	277	167	278	168
rect	277	168	278	169
rect	277	170	278	171
rect	277	171	278	172
rect	277	173	278	174
rect	277	174	278	175
rect	277	176	278	177
rect	277	177	278	178
rect	277	179	278	180
rect	277	180	278	181
rect	277	181	278	182
rect	277	182	278	183
rect	277	183	278	184
rect	277	185	278	186
rect	277	186	278	187
rect	277	188	278	189
rect	277	189	278	190
rect	277	190	278	191
rect	277	191	278	192
rect	277	192	278	193
rect	277	193	278	194
rect	277	194	278	195
rect	277	195	278	196
rect	277	197	278	198
rect	277	198	278	199
rect	277	199	278	200
rect	277	200	278	201
rect	277	201	278	202
rect	277	202	278	203
rect	277	203	278	204
rect	277	204	278	205
rect	277	205	278	206
rect	277	206	278	207
rect	277	207	278	208
rect	277	208	278	209
rect	277	209	278	210
rect	277	210	278	211
rect	277	211	278	212
rect	277	212	278	213
rect	277	213	278	214
rect	277	214	278	215
rect	277	215	278	216
rect	277	216	278	217
rect	277	218	278	219
rect	278	0	279	1
rect	278	1	279	2
rect	278	2	279	3
rect	278	3	279	4
rect	278	4	279	5
rect	278	5	279	6
rect	278	6	279	7
rect	278	8	279	9
rect	278	9	279	10
rect	278	11	279	12
rect	278	12	279	13
rect	278	14	279	15
rect	278	15	279	16
rect	278	17	279	18
rect	278	18	279	19
rect	278	20	279	21
rect	278	21	279	22
rect	278	23	279	24
rect	278	24	279	25
rect	278	26	279	27
rect	278	27	279	28
rect	278	29	279	30
rect	278	30	279	31
rect	278	32	279	33
rect	278	33	279	34
rect	278	35	279	36
rect	278	36	279	37
rect	278	38	279	39
rect	278	39	279	40
rect	278	41	279	42
rect	278	42	279	43
rect	278	44	279	45
rect	278	45	279	46
rect	278	47	279	48
rect	278	48	279	49
rect	278	50	279	51
rect	278	51	279	52
rect	278	52	279	53
rect	278	53	279	54
rect	278	54	279	55
rect	278	56	279	57
rect	278	57	279	58
rect	278	58	279	59
rect	278	59	279	60
rect	278	60	279	61
rect	278	62	279	63
rect	278	63	279	64
rect	278	65	279	66
rect	278	66	279	67
rect	278	67	279	68
rect	278	68	279	69
rect	278	69	279	70
rect	278	70	279	71
rect	278	71	279	72
rect	278	72	279	73
rect	278	73	279	74
rect	278	74	279	75
rect	278	75	279	76
rect	278	76	279	77
rect	278	77	279	78
rect	278	78	279	79
rect	278	80	279	81
rect	278	81	279	82
rect	278	83	279	84
rect	278	84	279	85
rect	278	86	279	87
rect	278	87	279	88
rect	278	89	279	90
rect	278	90	279	91
rect	278	91	279	92
rect	278	92	279	93
rect	278	93	279	94
rect	278	94	279	95
rect	278	95	279	96
rect	278	96	279	97
rect	278	97	279	98
rect	278	98	279	99
rect	278	99	279	100
rect	278	100	279	101
rect	278	101	279	102
rect	278	102	279	103
rect	278	103	279	104
rect	278	104	279	105
rect	278	105	279	106
rect	278	106	279	107
rect	278	107	279	108
rect	278	108	279	109
rect	278	110	279	111
rect	278	111	279	112
rect	278	112	279	113
rect	278	113	279	114
rect	278	114	279	115
rect	278	116	279	117
rect	278	117	279	118
rect	278	119	279	120
rect	278	120	279	121
rect	278	121	279	122
rect	278	122	279	123
rect	278	123	279	124
rect	278	125	279	126
rect	278	126	279	127
rect	278	127	279	128
rect	278	128	279	129
rect	278	129	279	130
rect	278	130	279	131
rect	278	131	279	132
rect	278	132	279	133
rect	278	134	279	135
rect	278	135	279	136
rect	278	137	279	138
rect	278	138	279	139
rect	278	140	279	141
rect	278	141	279	142
rect	278	142	279	143
rect	278	143	279	144
rect	278	144	279	145
rect	278	145	279	146
rect	278	146	279	147
rect	278	147	279	148
rect	278	149	279	150
rect	278	150	279	151
rect	278	152	279	153
rect	278	153	279	154
rect	278	154	279	155
rect	278	155	279	156
rect	278	156	279	157
rect	278	158	279	159
rect	278	159	279	160
rect	278	161	279	162
rect	278	162	279	163
rect	278	164	279	165
rect	278	165	279	166
rect	278	167	279	168
rect	278	168	279	169
rect	278	170	279	171
rect	278	171	279	172
rect	278	173	279	174
rect	278	174	279	175
rect	278	176	279	177
rect	278	177	279	178
rect	278	179	279	180
rect	278	180	279	181
rect	278	181	279	182
rect	278	182	279	183
rect	278	183	279	184
rect	278	185	279	186
rect	278	186	279	187
rect	278	188	279	189
rect	278	189	279	190
rect	278	190	279	191
rect	278	191	279	192
rect	278	192	279	193
rect	278	193	279	194
rect	278	194	279	195
rect	278	195	279	196
rect	278	197	279	198
rect	278	198	279	199
rect	278	199	279	200
rect	278	200	279	201
rect	278	201	279	202
rect	278	202	279	203
rect	278	203	279	204
rect	278	204	279	205
rect	278	205	279	206
rect	278	206	279	207
rect	278	207	279	208
rect	278	208	279	209
rect	278	209	279	210
rect	278	210	279	211
rect	278	211	279	212
rect	278	212	279	213
rect	278	213	279	214
rect	278	214	279	215
rect	278	215	279	216
rect	278	216	279	217
rect	278	218	279	219
rect	279	0	280	1
rect	279	1	280	2
rect	279	2	280	3
rect	279	3	280	4
rect	279	4	280	5
rect	279	5	280	6
rect	279	6	280	7
rect	279	8	280	9
rect	279	9	280	10
rect	279	11	280	12
rect	279	12	280	13
rect	279	14	280	15
rect	279	15	280	16
rect	279	17	280	18
rect	279	18	280	19
rect	279	20	280	21
rect	279	21	280	22
rect	279	23	280	24
rect	279	24	280	25
rect	279	26	280	27
rect	279	27	280	28
rect	279	29	280	30
rect	279	30	280	31
rect	279	32	280	33
rect	279	33	280	34
rect	279	35	280	36
rect	279	36	280	37
rect	279	38	280	39
rect	279	39	280	40
rect	279	41	280	42
rect	279	42	280	43
rect	279	44	280	45
rect	279	45	280	46
rect	279	47	280	48
rect	279	48	280	49
rect	279	50	280	51
rect	279	51	280	52
rect	279	52	280	53
rect	279	53	280	54
rect	279	54	280	55
rect	279	56	280	57
rect	279	57	280	58
rect	279	58	280	59
rect	279	59	280	60
rect	279	60	280	61
rect	279	62	280	63
rect	279	63	280	64
rect	279	65	280	66
rect	279	66	280	67
rect	279	67	280	68
rect	279	68	280	69
rect	279	69	280	70
rect	279	70	280	71
rect	279	71	280	72
rect	279	72	280	73
rect	279	73	280	74
rect	279	74	280	75
rect	279	75	280	76
rect	279	76	280	77
rect	279	77	280	78
rect	279	78	280	79
rect	279	80	280	81
rect	279	81	280	82
rect	279	83	280	84
rect	279	84	280	85
rect	279	86	280	87
rect	279	87	280	88
rect	279	89	280	90
rect	279	90	280	91
rect	279	91	280	92
rect	279	92	280	93
rect	279	93	280	94
rect	279	94	280	95
rect	279	95	280	96
rect	279	96	280	97
rect	279	97	280	98
rect	279	98	280	99
rect	279	99	280	100
rect	279	100	280	101
rect	279	101	280	102
rect	279	102	280	103
rect	279	103	280	104
rect	279	104	280	105
rect	279	105	280	106
rect	279	106	280	107
rect	279	107	280	108
rect	279	108	280	109
rect	279	110	280	111
rect	279	111	280	112
rect	279	112	280	113
rect	279	113	280	114
rect	279	114	280	115
rect	279	116	280	117
rect	279	117	280	118
rect	279	119	280	120
rect	279	120	280	121
rect	279	121	280	122
rect	279	122	280	123
rect	279	123	280	124
rect	279	125	280	126
rect	279	126	280	127
rect	279	127	280	128
rect	279	128	280	129
rect	279	129	280	130
rect	279	130	280	131
rect	279	131	280	132
rect	279	132	280	133
rect	279	134	280	135
rect	279	135	280	136
rect	279	137	280	138
rect	279	138	280	139
rect	279	140	280	141
rect	279	141	280	142
rect	279	142	280	143
rect	279	143	280	144
rect	279	144	280	145
rect	279	145	280	146
rect	279	146	280	147
rect	279	147	280	148
rect	279	149	280	150
rect	279	150	280	151
rect	279	152	280	153
rect	279	153	280	154
rect	279	154	280	155
rect	279	155	280	156
rect	279	156	280	157
rect	279	158	280	159
rect	279	159	280	160
rect	279	161	280	162
rect	279	162	280	163
rect	279	164	280	165
rect	279	165	280	166
rect	279	167	280	168
rect	279	168	280	169
rect	279	170	280	171
rect	279	171	280	172
rect	279	173	280	174
rect	279	174	280	175
rect	279	176	280	177
rect	279	177	280	178
rect	279	179	280	180
rect	279	180	280	181
rect	279	181	280	182
rect	279	182	280	183
rect	279	183	280	184
rect	279	185	280	186
rect	279	186	280	187
rect	279	188	280	189
rect	279	189	280	190
rect	279	190	280	191
rect	279	191	280	192
rect	279	192	280	193
rect	279	193	280	194
rect	279	194	280	195
rect	279	195	280	196
rect	279	197	280	198
rect	279	198	280	199
rect	279	199	280	200
rect	279	200	280	201
rect	279	201	280	202
rect	279	202	280	203
rect	279	203	280	204
rect	279	204	280	205
rect	279	205	280	206
rect	279	206	280	207
rect	279	207	280	208
rect	279	208	280	209
rect	279	209	280	210
rect	279	210	280	211
rect	279	211	280	212
rect	279	212	280	213
rect	279	213	280	214
rect	279	214	280	215
rect	279	215	280	216
rect	279	216	280	217
rect	279	218	280	219
rect	280	0	281	1
rect	280	1	281	2
rect	280	2	281	3
rect	280	3	281	4
rect	280	4	281	5
rect	280	5	281	6
rect	280	6	281	7
rect	280	8	281	9
rect	280	9	281	10
rect	280	11	281	12
rect	280	12	281	13
rect	280	14	281	15
rect	280	15	281	16
rect	280	17	281	18
rect	280	18	281	19
rect	280	20	281	21
rect	280	21	281	22
rect	280	23	281	24
rect	280	24	281	25
rect	280	26	281	27
rect	280	27	281	28
rect	280	29	281	30
rect	280	30	281	31
rect	280	32	281	33
rect	280	33	281	34
rect	280	35	281	36
rect	280	36	281	37
rect	280	38	281	39
rect	280	39	281	40
rect	280	41	281	42
rect	280	42	281	43
rect	280	44	281	45
rect	280	45	281	46
rect	280	47	281	48
rect	280	48	281	49
rect	280	50	281	51
rect	280	51	281	52
rect	280	52	281	53
rect	280	53	281	54
rect	280	54	281	55
rect	280	56	281	57
rect	280	57	281	58
rect	280	58	281	59
rect	280	59	281	60
rect	280	60	281	61
rect	280	62	281	63
rect	280	63	281	64
rect	280	65	281	66
rect	280	66	281	67
rect	280	67	281	68
rect	280	68	281	69
rect	280	69	281	70
rect	280	70	281	71
rect	280	71	281	72
rect	280	72	281	73
rect	280	73	281	74
rect	280	74	281	75
rect	280	75	281	76
rect	280	76	281	77
rect	280	77	281	78
rect	280	78	281	79
rect	280	80	281	81
rect	280	81	281	82
rect	280	83	281	84
rect	280	84	281	85
rect	280	86	281	87
rect	280	87	281	88
rect	280	89	281	90
rect	280	90	281	91
rect	280	91	281	92
rect	280	92	281	93
rect	280	93	281	94
rect	280	94	281	95
rect	280	95	281	96
rect	280	96	281	97
rect	280	97	281	98
rect	280	98	281	99
rect	280	99	281	100
rect	280	100	281	101
rect	280	101	281	102
rect	280	102	281	103
rect	280	103	281	104
rect	280	104	281	105
rect	280	105	281	106
rect	280	106	281	107
rect	280	107	281	108
rect	280	108	281	109
rect	280	110	281	111
rect	280	111	281	112
rect	280	112	281	113
rect	280	113	281	114
rect	280	114	281	115
rect	280	116	281	117
rect	280	117	281	118
rect	280	119	281	120
rect	280	120	281	121
rect	280	121	281	122
rect	280	122	281	123
rect	280	123	281	124
rect	280	125	281	126
rect	280	126	281	127
rect	280	127	281	128
rect	280	128	281	129
rect	280	129	281	130
rect	280	130	281	131
rect	280	131	281	132
rect	280	132	281	133
rect	280	134	281	135
rect	280	135	281	136
rect	280	137	281	138
rect	280	138	281	139
rect	280	140	281	141
rect	280	141	281	142
rect	280	142	281	143
rect	280	143	281	144
rect	280	144	281	145
rect	280	145	281	146
rect	280	146	281	147
rect	280	147	281	148
rect	280	149	281	150
rect	280	150	281	151
rect	280	152	281	153
rect	280	153	281	154
rect	280	154	281	155
rect	280	155	281	156
rect	280	156	281	157
rect	280	158	281	159
rect	280	159	281	160
rect	280	161	281	162
rect	280	162	281	163
rect	280	164	281	165
rect	280	165	281	166
rect	280	167	281	168
rect	280	168	281	169
rect	280	170	281	171
rect	280	171	281	172
rect	280	173	281	174
rect	280	174	281	175
rect	280	176	281	177
rect	280	177	281	178
rect	280	179	281	180
rect	280	180	281	181
rect	280	181	281	182
rect	280	182	281	183
rect	280	183	281	184
rect	280	185	281	186
rect	280	186	281	187
rect	280	188	281	189
rect	280	189	281	190
rect	280	190	281	191
rect	280	191	281	192
rect	280	192	281	193
rect	280	193	281	194
rect	280	194	281	195
rect	280	195	281	196
rect	280	197	281	198
rect	280	198	281	199
rect	280	199	281	200
rect	280	200	281	201
rect	280	201	281	202
rect	280	202	281	203
rect	280	203	281	204
rect	280	204	281	205
rect	280	205	281	206
rect	280	206	281	207
rect	280	207	281	208
rect	280	208	281	209
rect	280	209	281	210
rect	280	210	281	211
rect	280	211	281	212
rect	280	212	281	213
rect	280	213	281	214
rect	280	214	281	215
rect	280	215	281	216
rect	280	216	281	217
rect	280	218	281	219
rect	281	0	282	1
rect	281	1	282	2
rect	281	2	282	3
rect	281	3	282	4
rect	281	4	282	5
rect	281	5	282	6
rect	281	6	282	7
rect	281	8	282	9
rect	281	9	282	10
rect	281	11	282	12
rect	281	12	282	13
rect	281	14	282	15
rect	281	15	282	16
rect	281	17	282	18
rect	281	18	282	19
rect	281	20	282	21
rect	281	21	282	22
rect	281	23	282	24
rect	281	24	282	25
rect	281	26	282	27
rect	281	27	282	28
rect	281	29	282	30
rect	281	30	282	31
rect	281	32	282	33
rect	281	33	282	34
rect	281	35	282	36
rect	281	36	282	37
rect	281	38	282	39
rect	281	39	282	40
rect	281	41	282	42
rect	281	42	282	43
rect	281	44	282	45
rect	281	45	282	46
rect	281	47	282	48
rect	281	48	282	49
rect	281	50	282	51
rect	281	51	282	52
rect	281	52	282	53
rect	281	53	282	54
rect	281	54	282	55
rect	281	56	282	57
rect	281	57	282	58
rect	281	58	282	59
rect	281	59	282	60
rect	281	60	282	61
rect	281	62	282	63
rect	281	63	282	64
rect	281	65	282	66
rect	281	66	282	67
rect	281	67	282	68
rect	281	68	282	69
rect	281	69	282	70
rect	281	70	282	71
rect	281	71	282	72
rect	281	72	282	73
rect	281	73	282	74
rect	281	74	282	75
rect	281	75	282	76
rect	281	76	282	77
rect	281	77	282	78
rect	281	78	282	79
rect	281	80	282	81
rect	281	81	282	82
rect	281	83	282	84
rect	281	84	282	85
rect	281	86	282	87
rect	281	87	282	88
rect	281	89	282	90
rect	281	90	282	91
rect	281	91	282	92
rect	281	92	282	93
rect	281	93	282	94
rect	281	94	282	95
rect	281	95	282	96
rect	281	96	282	97
rect	281	97	282	98
rect	281	98	282	99
rect	281	99	282	100
rect	281	100	282	101
rect	281	101	282	102
rect	281	102	282	103
rect	281	103	282	104
rect	281	104	282	105
rect	281	105	282	106
rect	281	106	282	107
rect	281	107	282	108
rect	281	108	282	109
rect	281	110	282	111
rect	281	111	282	112
rect	281	112	282	113
rect	281	113	282	114
rect	281	114	282	115
rect	281	116	282	117
rect	281	117	282	118
rect	281	119	282	120
rect	281	120	282	121
rect	281	121	282	122
rect	281	122	282	123
rect	281	123	282	124
rect	281	125	282	126
rect	281	126	282	127
rect	281	127	282	128
rect	281	128	282	129
rect	281	129	282	130
rect	281	130	282	131
rect	281	131	282	132
rect	281	132	282	133
rect	281	134	282	135
rect	281	135	282	136
rect	281	137	282	138
rect	281	138	282	139
rect	281	140	282	141
rect	281	141	282	142
rect	281	142	282	143
rect	281	143	282	144
rect	281	144	282	145
rect	281	145	282	146
rect	281	146	282	147
rect	281	147	282	148
rect	281	149	282	150
rect	281	150	282	151
rect	281	152	282	153
rect	281	153	282	154
rect	281	154	282	155
rect	281	155	282	156
rect	281	156	282	157
rect	281	158	282	159
rect	281	159	282	160
rect	281	161	282	162
rect	281	162	282	163
rect	281	164	282	165
rect	281	165	282	166
rect	281	167	282	168
rect	281	168	282	169
rect	281	170	282	171
rect	281	171	282	172
rect	281	173	282	174
rect	281	174	282	175
rect	281	176	282	177
rect	281	177	282	178
rect	281	179	282	180
rect	281	180	282	181
rect	281	181	282	182
rect	281	182	282	183
rect	281	183	282	184
rect	281	185	282	186
rect	281	186	282	187
rect	281	188	282	189
rect	281	189	282	190
rect	281	190	282	191
rect	281	191	282	192
rect	281	192	282	193
rect	281	193	282	194
rect	281	194	282	195
rect	281	195	282	196
rect	281	197	282	198
rect	281	198	282	199
rect	281	199	282	200
rect	281	200	282	201
rect	281	201	282	202
rect	281	202	282	203
rect	281	203	282	204
rect	281	204	282	205
rect	281	205	282	206
rect	281	206	282	207
rect	281	207	282	208
rect	281	208	282	209
rect	281	209	282	210
rect	281	210	282	211
rect	281	211	282	212
rect	281	212	282	213
rect	281	213	282	214
rect	281	214	282	215
rect	281	215	282	216
rect	281	216	282	217
rect	281	218	282	219
rect	288	0	289	1
rect	288	1	289	2
rect	288	2	289	3
rect	288	3	289	4
rect	288	4	289	5
rect	288	5	289	6
rect	288	6	289	7
rect	288	8	289	9
rect	288	9	289	10
rect	288	11	289	12
rect	288	12	289	13
rect	288	14	289	15
rect	288	15	289	16
rect	288	16	289	17
rect	288	17	289	18
rect	288	18	289	19
rect	288	20	289	21
rect	288	21	289	22
rect	288	23	289	24
rect	288	24	289	25
rect	288	25	289	26
rect	288	26	289	27
rect	288	27	289	28
rect	288	29	289	30
rect	288	30	289	31
rect	288	32	289	33
rect	288	33	289	34
rect	288	34	289	35
rect	288	35	289	36
rect	288	36	289	37
rect	288	38	289	39
rect	288	39	289	40
rect	288	41	289	42
rect	288	42	289	43
rect	288	43	289	44
rect	288	44	289	45
rect	288	45	289	46
rect	288	47	289	48
rect	288	48	289	49
rect	288	50	289	51
rect	288	51	289	52
rect	288	52	289	53
rect	288	53	289	54
rect	288	54	289	55
rect	288	56	289	57
rect	288	57	289	58
rect	288	58	289	59
rect	288	59	289	60
rect	288	60	289	61
rect	288	61	289	62
rect	288	62	289	63
rect	288	63	289	64
rect	288	65	289	66
rect	288	66	289	67
rect	288	67	289	68
rect	288	68	289	69
rect	288	69	289	70
rect	288	70	289	71
rect	288	71	289	72
rect	288	72	289	73
rect	288	73	289	74
rect	288	74	289	75
rect	288	75	289	76
rect	288	76	289	77
rect	288	77	289	78
rect	288	78	289	79
rect	288	79	289	80
rect	288	80	289	81
rect	288	81	289	82
rect	288	83	289	84
rect	288	84	289	85
rect	288	86	289	87
rect	288	87	289	88
rect	288	88	289	89
rect	288	89	289	90
rect	288	90	289	91
rect	288	91	289	92
rect	288	92	289	93
rect	288	93	289	94
rect	288	94	289	95
rect	288	95	289	96
rect	288	96	289	97
rect	288	97	289	98
rect	288	98	289	99
rect	288	99	289	100
rect	288	100	289	101
rect	288	101	289	102
rect	288	102	289	103
rect	288	103	289	104
rect	288	104	289	105
rect	288	105	289	106
rect	288	106	289	107
rect	288	107	289	108
rect	288	108	289	109
rect	288	109	289	110
rect	288	110	289	111
rect	288	111	289	112
rect	288	112	289	113
rect	288	113	289	114
rect	288	114	289	115
rect	288	116	289	117
rect	288	117	289	118
rect	288	118	289	119
rect	288	119	289	120
rect	288	120	289	121
rect	288	121	289	122
rect	288	122	289	123
rect	288	123	289	124
rect	288	125	289	126
rect	288	126	289	127
rect	288	127	289	128
rect	288	128	289	129
rect	288	129	289	130
rect	288	130	289	131
rect	288	131	289	132
rect	288	132	289	133
rect	288	133	289	134
rect	288	134	289	135
rect	288	135	289	136
rect	288	137	289	138
rect	288	138	289	139
rect	288	140	289	141
rect	288	141	289	142
rect	288	142	289	143
rect	288	143	289	144
rect	288	144	289	145
rect	288	145	289	146
rect	288	146	289	147
rect	288	147	289	148
rect	288	149	289	150
rect	288	150	289	151
rect	288	152	289	153
rect	288	153	289	154
rect	288	154	289	155
rect	288	155	289	156
rect	288	156	289	157
rect	288	158	289	159
rect	288	159	289	160
rect	288	161	289	162
rect	288	162	289	163
rect	288	163	289	164
rect	288	164	289	165
rect	288	165	289	166
rect	288	167	289	168
rect	288	168	289	169
rect	288	170	289	171
rect	288	171	289	172
rect	288	172	289	173
rect	288	173	289	174
rect	288	174	289	175
rect	288	176	289	177
rect	288	177	289	178
rect	288	179	289	180
rect	288	180	289	181
rect	288	181	289	182
rect	288	182	289	183
rect	288	183	289	184
rect	288	184	289	185
rect	288	185	289	186
rect	288	186	289	187
rect	288	187	289	188
rect	288	188	289	189
rect	288	189	289	190
rect	288	190	289	191
rect	288	191	289	192
rect	288	192	289	193
rect	288	193	289	194
rect	288	194	289	195
rect	288	195	289	196
rect	288	196	289	197
rect	288	197	289	198
rect	288	198	289	199
rect	288	199	289	200
rect	288	200	289	201
rect	288	201	289	202
rect	288	202	289	203
rect	288	203	289	204
rect	288	204	289	205
rect	288	205	289	206
rect	288	206	289	207
rect	288	207	289	208
rect	288	208	289	209
rect	288	209	289	210
rect	288	210	289	211
rect	288	211	289	212
rect	288	212	289	213
rect	288	213	289	214
rect	288	214	289	215
rect	288	215	289	216
rect	288	216	289	217
rect	288	217	289	218
rect	288	218	289	219
rect	290	0	291	1
rect	290	1	291	2
rect	290	2	291	3
rect	290	3	291	4
rect	290	4	291	5
rect	290	5	291	6
rect	290	6	291	7
rect	290	8	291	9
rect	290	9	291	10
rect	290	11	291	12
rect	290	12	291	13
rect	290	14	291	15
rect	290	15	291	16
rect	290	16	291	17
rect	290	17	291	18
rect	290	18	291	19
rect	290	20	291	21
rect	290	21	291	22
rect	290	23	291	24
rect	290	24	291	25
rect	290	25	291	26
rect	290	26	291	27
rect	290	27	291	28
rect	290	29	291	30
rect	290	30	291	31
rect	290	32	291	33
rect	290	33	291	34
rect	290	34	291	35
rect	290	35	291	36
rect	290	36	291	37
rect	290	38	291	39
rect	290	39	291	40
rect	290	41	291	42
rect	290	42	291	43
rect	290	43	291	44
rect	290	44	291	45
rect	290	45	291	46
rect	290	47	291	48
rect	290	48	291	49
rect	290	50	291	51
rect	290	51	291	52
rect	290	52	291	53
rect	290	53	291	54
rect	290	54	291	55
rect	290	56	291	57
rect	290	57	291	58
rect	290	58	291	59
rect	290	59	291	60
rect	290	60	291	61
rect	290	61	291	62
rect	290	62	291	63
rect	290	63	291	64
rect	290	65	291	66
rect	290	66	291	67
rect	290	67	291	68
rect	290	68	291	69
rect	290	69	291	70
rect	290	70	291	71
rect	290	71	291	72
rect	290	72	291	73
rect	290	73	291	74
rect	290	74	291	75
rect	290	75	291	76
rect	290	76	291	77
rect	290	77	291	78
rect	290	78	291	79
rect	290	79	291	80
rect	290	80	291	81
rect	290	81	291	82
rect	290	83	291	84
rect	290	84	291	85
rect	290	86	291	87
rect	290	87	291	88
rect	290	88	291	89
rect	290	89	291	90
rect	290	90	291	91
rect	290	91	291	92
rect	290	92	291	93
rect	290	93	291	94
rect	290	94	291	95
rect	290	95	291	96
rect	290	96	291	97
rect	290	97	291	98
rect	290	98	291	99
rect	290	99	291	100
rect	290	100	291	101
rect	290	101	291	102
rect	290	102	291	103
rect	290	103	291	104
rect	290	104	291	105
rect	290	105	291	106
rect	290	106	291	107
rect	290	107	291	108
rect	290	108	291	109
rect	290	109	291	110
rect	290	110	291	111
rect	290	111	291	112
rect	290	112	291	113
rect	290	113	291	114
rect	290	114	291	115
rect	290	116	291	117
rect	290	117	291	118
rect	290	118	291	119
rect	290	119	291	120
rect	290	120	291	121
rect	290	121	291	122
rect	290	122	291	123
rect	290	123	291	124
rect	290	125	291	126
rect	290	126	291	127
rect	290	127	291	128
rect	290	128	291	129
rect	290	129	291	130
rect	290	130	291	131
rect	290	131	291	132
rect	290	132	291	133
rect	290	133	291	134
rect	290	134	291	135
rect	290	135	291	136
rect	290	137	291	138
rect	290	138	291	139
rect	290	140	291	141
rect	290	141	291	142
rect	290	142	291	143
rect	290	143	291	144
rect	290	144	291	145
rect	290	145	291	146
rect	290	146	291	147
rect	290	147	291	148
rect	290	149	291	150
rect	290	150	291	151
rect	290	152	291	153
rect	290	153	291	154
rect	290	154	291	155
rect	290	155	291	156
rect	290	156	291	157
rect	290	158	291	159
rect	290	159	291	160
rect	290	161	291	162
rect	290	162	291	163
rect	290	163	291	164
rect	290	164	291	165
rect	290	165	291	166
rect	290	167	291	168
rect	290	168	291	169
rect	290	170	291	171
rect	290	171	291	172
rect	290	172	291	173
rect	290	173	291	174
rect	290	174	291	175
rect	290	176	291	177
rect	290	177	291	178
rect	290	179	291	180
rect	290	180	291	181
rect	290	181	291	182
rect	290	182	291	183
rect	290	183	291	184
rect	290	184	291	185
rect	290	185	291	186
rect	290	186	291	187
rect	290	187	291	188
rect	290	188	291	189
rect	290	189	291	190
rect	290	190	291	191
rect	290	191	291	192
rect	290	192	291	193
rect	290	193	291	194
rect	290	194	291	195
rect	291	0	292	1
rect	291	1	292	2
rect	291	2	292	3
rect	291	3	292	4
rect	291	4	292	5
rect	291	5	292	6
rect	291	6	292	7
rect	291	8	292	9
rect	291	9	292	10
rect	291	11	292	12
rect	291	12	292	13
rect	291	14	292	15
rect	291	15	292	16
rect	291	16	292	17
rect	291	17	292	18
rect	291	18	292	19
rect	291	20	292	21
rect	291	21	292	22
rect	291	23	292	24
rect	291	24	292	25
rect	291	25	292	26
rect	291	26	292	27
rect	291	27	292	28
rect	291	29	292	30
rect	291	30	292	31
rect	291	32	292	33
rect	291	33	292	34
rect	291	34	292	35
rect	291	35	292	36
rect	291	36	292	37
rect	291	38	292	39
rect	291	39	292	40
rect	291	41	292	42
rect	291	42	292	43
rect	291	43	292	44
rect	291	44	292	45
rect	291	45	292	46
rect	291	47	292	48
rect	291	48	292	49
rect	291	50	292	51
rect	291	51	292	52
rect	291	52	292	53
rect	291	53	292	54
rect	291	54	292	55
rect	291	56	292	57
rect	291	57	292	58
rect	291	58	292	59
rect	291	59	292	60
rect	291	60	292	61
rect	291	61	292	62
rect	291	62	292	63
rect	291	63	292	64
rect	291	65	292	66
rect	291	66	292	67
rect	291	67	292	68
rect	291	68	292	69
rect	291	69	292	70
rect	291	70	292	71
rect	291	71	292	72
rect	291	72	292	73
rect	291	73	292	74
rect	291	74	292	75
rect	291	75	292	76
rect	291	76	292	77
rect	291	77	292	78
rect	291	78	292	79
rect	291	79	292	80
rect	291	80	292	81
rect	291	81	292	82
rect	291	83	292	84
rect	291	84	292	85
rect	291	86	292	87
rect	291	87	292	88
rect	291	88	292	89
rect	291	89	292	90
rect	291	90	292	91
rect	291	91	292	92
rect	291	92	292	93
rect	291	93	292	94
rect	291	94	292	95
rect	291	95	292	96
rect	291	96	292	97
rect	291	97	292	98
rect	291	98	292	99
rect	291	99	292	100
rect	291	100	292	101
rect	291	101	292	102
rect	291	102	292	103
rect	291	103	292	104
rect	291	104	292	105
rect	291	105	292	106
rect	291	106	292	107
rect	291	107	292	108
rect	291	108	292	109
rect	291	109	292	110
rect	291	110	292	111
rect	291	111	292	112
rect	291	112	292	113
rect	291	113	292	114
rect	291	114	292	115
rect	291	116	292	117
rect	291	117	292	118
rect	291	118	292	119
rect	291	119	292	120
rect	291	120	292	121
rect	291	121	292	122
rect	291	122	292	123
rect	291	123	292	124
rect	291	125	292	126
rect	291	126	292	127
rect	291	127	292	128
rect	291	128	292	129
rect	291	129	292	130
rect	291	130	292	131
rect	291	131	292	132
rect	291	132	292	133
rect	291	133	292	134
rect	291	134	292	135
rect	291	135	292	136
rect	291	137	292	138
rect	291	138	292	139
rect	291	140	292	141
rect	291	141	292	142
rect	291	142	292	143
rect	291	143	292	144
rect	291	144	292	145
rect	291	145	292	146
rect	291	146	292	147
rect	291	147	292	148
rect	291	149	292	150
rect	291	150	292	151
rect	291	152	292	153
rect	291	153	292	154
rect	291	154	292	155
rect	291	155	292	156
rect	291	156	292	157
rect	291	158	292	159
rect	291	159	292	160
rect	291	161	292	162
rect	291	162	292	163
rect	291	163	292	164
rect	291	164	292	165
rect	291	165	292	166
rect	291	167	292	168
rect	291	168	292	169
rect	291	170	292	171
rect	291	171	292	172
rect	291	172	292	173
rect	291	173	292	174
rect	291	174	292	175
rect	291	176	292	177
rect	291	177	292	178
rect	291	179	292	180
rect	291	180	292	181
rect	291	181	292	182
rect	291	182	292	183
rect	291	183	292	184
rect	291	184	292	185
rect	291	185	292	186
rect	291	186	292	187
rect	291	187	292	188
rect	291	188	292	189
rect	291	189	292	190
rect	291	190	292	191
rect	291	191	292	192
rect	291	192	292	193
rect	291	193	292	194
rect	291	194	292	195
rect	292	0	293	1
rect	292	1	293	2
rect	292	2	293	3
rect	292	3	293	4
rect	292	4	293	5
rect	292	5	293	6
rect	292	6	293	7
rect	292	8	293	9
rect	292	9	293	10
rect	292	11	293	12
rect	292	12	293	13
rect	292	14	293	15
rect	292	15	293	16
rect	292	16	293	17
rect	292	17	293	18
rect	292	18	293	19
rect	292	19	293	20
rect	292	20	293	21
rect	292	21	293	22
rect	292	23	293	24
rect	292	24	293	25
rect	292	25	293	26
rect	292	26	293	27
rect	292	27	293	28
rect	292	29	293	30
rect	292	30	293	31
rect	292	32	293	33
rect	292	33	293	34
rect	292	34	293	35
rect	292	35	293	36
rect	292	36	293	37
rect	292	38	293	39
rect	292	39	293	40
rect	292	40	293	41
rect	292	41	293	42
rect	292	42	293	43
rect	292	43	293	44
rect	292	44	293	45
rect	292	45	293	46
rect	292	46	293	47
rect	292	47	293	48
rect	292	48	293	49
rect	292	50	293	51
rect	292	51	293	52
rect	292	52	293	53
rect	292	53	293	54
rect	292	54	293	55
rect	292	55	293	56
rect	292	56	293	57
rect	292	57	293	58
rect	292	58	293	59
rect	292	59	293	60
rect	292	60	293	61
rect	292	61	293	62
rect	292	62	293	63
rect	292	63	293	64
rect	292	65	293	66
rect	292	66	293	67
rect	292	67	293	68
rect	292	68	293	69
rect	292	69	293	70
rect	292	70	293	71
rect	292	71	293	72
rect	292	72	293	73
rect	292	73	293	74
rect	292	74	293	75
rect	292	75	293	76
rect	292	76	293	77
rect	292	77	293	78
rect	292	78	293	79
rect	292	79	293	80
rect	292	80	293	81
rect	292	81	293	82
rect	292	83	293	84
rect	292	84	293	85
rect	292	86	293	87
rect	292	87	293	88
rect	292	88	293	89
rect	292	89	293	90
rect	292	90	293	91
rect	292	91	293	92
rect	292	92	293	93
rect	292	93	293	94
rect	292	94	293	95
rect	292	95	293	96
rect	292	96	293	97
rect	292	97	293	98
rect	292	98	293	99
rect	292	99	293	100
rect	292	100	293	101
rect	292	101	293	102
rect	292	102	293	103
rect	292	103	293	104
rect	292	104	293	105
rect	292	105	293	106
rect	292	106	293	107
rect	292	107	293	108
rect	292	108	293	109
rect	292	109	293	110
rect	292	110	293	111
rect	292	111	293	112
rect	292	112	293	113
rect	292	113	293	114
rect	292	114	293	115
rect	292	116	293	117
rect	292	117	293	118
rect	292	118	293	119
rect	292	119	293	120
rect	292	120	293	121
rect	292	121	293	122
rect	292	122	293	123
rect	292	123	293	124
rect	292	125	293	126
rect	292	126	293	127
rect	292	127	293	128
rect	292	128	293	129
rect	292	129	293	130
rect	292	130	293	131
rect	292	131	293	132
rect	292	132	293	133
rect	292	133	293	134
rect	292	134	293	135
rect	292	135	293	136
rect	292	137	293	138
rect	292	138	293	139
rect	292	140	293	141
rect	292	141	293	142
rect	292	142	293	143
rect	292	143	293	144
rect	292	144	293	145
rect	292	145	293	146
rect	292	146	293	147
rect	292	147	293	148
rect	292	148	293	149
rect	292	149	293	150
rect	292	150	293	151
rect	292	152	293	153
rect	292	153	293	154
rect	292	154	293	155
rect	292	155	293	156
rect	292	156	293	157
rect	292	157	293	158
rect	292	158	293	159
rect	292	159	293	160
rect	292	161	293	162
rect	292	162	293	163
rect	292	163	293	164
rect	292	164	293	165
rect	292	165	293	166
rect	292	167	293	168
rect	292	168	293	169
rect	292	170	293	171
rect	292	171	293	172
rect	292	172	293	173
rect	292	173	293	174
rect	292	174	293	175
rect	292	175	293	176
rect	292	176	293	177
rect	292	177	293	178
rect	292	178	293	179
rect	292	179	293	180
rect	292	180	293	181
rect	292	181	293	182
rect	292	182	293	183
rect	292	183	293	184
rect	292	184	293	185
rect	292	185	293	186
rect	292	186	293	187
rect	292	187	293	188
rect	292	188	293	189
rect	292	189	293	190
rect	292	190	293	191
rect	292	191	293	192
rect	292	192	293	193
rect	292	193	293	194
rect	292	194	293	195
rect	293	0	294	1
rect	293	1	294	2
rect	293	2	294	3
rect	293	3	294	4
rect	293	4	294	5
rect	293	5	294	6
rect	293	6	294	7
rect	293	8	294	9
rect	293	9	294	10
rect	293	11	294	12
rect	293	12	294	13
rect	293	14	294	15
rect	293	15	294	16
rect	293	16	294	17
rect	293	17	294	18
rect	293	18	294	19
rect	293	19	294	20
rect	293	20	294	21
rect	293	21	294	22
rect	293	23	294	24
rect	293	24	294	25
rect	293	25	294	26
rect	293	26	294	27
rect	293	27	294	28
rect	293	29	294	30
rect	293	30	294	31
rect	293	32	294	33
rect	293	33	294	34
rect	293	34	294	35
rect	293	35	294	36
rect	293	36	294	37
rect	293	38	294	39
rect	293	39	294	40
rect	293	40	294	41
rect	293	41	294	42
rect	293	42	294	43
rect	293	43	294	44
rect	293	44	294	45
rect	293	45	294	46
rect	293	46	294	47
rect	293	47	294	48
rect	293	48	294	49
rect	293	50	294	51
rect	293	51	294	52
rect	293	52	294	53
rect	293	53	294	54
rect	293	54	294	55
rect	293	55	294	56
rect	293	56	294	57
rect	293	57	294	58
rect	293	58	294	59
rect	293	59	294	60
rect	293	60	294	61
rect	293	61	294	62
rect	293	62	294	63
rect	293	63	294	64
rect	293	65	294	66
rect	293	66	294	67
rect	293	67	294	68
rect	293	68	294	69
rect	293	69	294	70
rect	293	70	294	71
rect	293	71	294	72
rect	293	72	294	73
rect	293	73	294	74
rect	293	74	294	75
rect	293	75	294	76
rect	293	76	294	77
rect	293	77	294	78
rect	293	78	294	79
rect	293	80	294	81
rect	293	81	294	82
rect	293	83	294	84
rect	293	84	294	85
rect	293	86	294	87
rect	293	87	294	88
rect	293	88	294	89
rect	293	89	294	90
rect	293	90	294	91
rect	293	91	294	92
rect	293	92	294	93
rect	293	93	294	94
rect	293	94	294	95
rect	293	95	294	96
rect	293	96	294	97
rect	293	97	294	98
rect	293	98	294	99
rect	293	99	294	100
rect	293	100	294	101
rect	293	101	294	102
rect	293	102	294	103
rect	293	103	294	104
rect	293	104	294	105
rect	293	105	294	106
rect	293	106	294	107
rect	293	107	294	108
rect	293	108	294	109
rect	293	109	294	110
rect	293	110	294	111
rect	293	111	294	112
rect	293	112	294	113
rect	293	113	294	114
rect	293	114	294	115
rect	293	116	294	117
rect	293	117	294	118
rect	293	118	294	119
rect	293	119	294	120
rect	293	120	294	121
rect	293	121	294	122
rect	293	122	294	123
rect	293	123	294	124
rect	293	125	294	126
rect	293	126	294	127
rect	293	127	294	128
rect	293	128	294	129
rect	293	129	294	130
rect	293	130	294	131
rect	293	131	294	132
rect	293	132	294	133
rect	293	133	294	134
rect	293	134	294	135
rect	293	135	294	136
rect	293	137	294	138
rect	293	138	294	139
rect	293	140	294	141
rect	293	141	294	142
rect	293	142	294	143
rect	293	143	294	144
rect	293	144	294	145
rect	293	145	294	146
rect	293	146	294	147
rect	293	147	294	148
rect	293	148	294	149
rect	293	149	294	150
rect	293	150	294	151
rect	293	152	294	153
rect	293	153	294	154
rect	293	154	294	155
rect	293	155	294	156
rect	293	156	294	157
rect	293	157	294	158
rect	293	158	294	159
rect	293	159	294	160
rect	293	161	294	162
rect	293	162	294	163
rect	293	163	294	164
rect	293	164	294	165
rect	293	165	294	166
rect	293	167	294	168
rect	293	168	294	169
rect	293	170	294	171
rect	293	171	294	172
rect	293	172	294	173
rect	293	173	294	174
rect	293	174	294	175
rect	293	175	294	176
rect	293	176	294	177
rect	293	177	294	178
rect	293	178	294	179
rect	293	179	294	180
rect	293	180	294	181
rect	293	181	294	182
rect	293	182	294	183
rect	293	183	294	184
rect	293	184	294	185
rect	293	185	294	186
rect	293	186	294	187
rect	293	187	294	188
rect	293	188	294	189
rect	293	189	294	190
rect	293	190	294	191
rect	293	191	294	192
rect	293	192	294	193
rect	293	193	294	194
rect	293	194	294	195
rect	294	0	295	1
rect	294	1	295	2
rect	294	2	295	3
rect	294	3	295	4
rect	294	4	295	5
rect	294	5	295	6
rect	294	6	295	7
rect	294	8	295	9
rect	294	9	295	10
rect	294	11	295	12
rect	294	12	295	13
rect	294	14	295	15
rect	294	15	295	16
rect	294	16	295	17
rect	294	17	295	18
rect	294	18	295	19
rect	294	19	295	20
rect	294	20	295	21
rect	294	21	295	22
rect	294	23	295	24
rect	294	24	295	25
rect	294	25	295	26
rect	294	26	295	27
rect	294	27	295	28
rect	294	29	295	30
rect	294	30	295	31
rect	294	32	295	33
rect	294	33	295	34
rect	294	34	295	35
rect	294	35	295	36
rect	294	36	295	37
rect	294	38	295	39
rect	294	39	295	40
rect	294	40	295	41
rect	294	41	295	42
rect	294	42	295	43
rect	294	43	295	44
rect	294	44	295	45
rect	294	45	295	46
rect	294	46	295	47
rect	294	47	295	48
rect	294	48	295	49
rect	294	50	295	51
rect	294	51	295	52
rect	294	52	295	53
rect	294	53	295	54
rect	294	54	295	55
rect	294	55	295	56
rect	294	56	295	57
rect	294	57	295	58
rect	294	58	295	59
rect	294	59	295	60
rect	294	60	295	61
rect	294	61	295	62
rect	294	62	295	63
rect	294	63	295	64
rect	294	65	295	66
rect	294	66	295	67
rect	294	67	295	68
rect	294	68	295	69
rect	294	69	295	70
rect	294	70	295	71
rect	294	71	295	72
rect	294	72	295	73
rect	294	73	295	74
rect	294	74	295	75
rect	294	75	295	76
rect	294	76	295	77
rect	294	77	295	78
rect	294	78	295	79
rect	294	80	295	81
rect	294	81	295	82
rect	294	83	295	84
rect	294	84	295	85
rect	294	86	295	87
rect	294	87	295	88
rect	294	88	295	89
rect	294	89	295	90
rect	294	90	295	91
rect	294	91	295	92
rect	294	92	295	93
rect	294	93	295	94
rect	294	94	295	95
rect	294	95	295	96
rect	294	96	295	97
rect	294	97	295	98
rect	294	98	295	99
rect	294	99	295	100
rect	294	100	295	101
rect	294	101	295	102
rect	294	102	295	103
rect	294	103	295	104
rect	294	104	295	105
rect	294	105	295	106
rect	294	106	295	107
rect	294	107	295	108
rect	294	108	295	109
rect	294	109	295	110
rect	294	110	295	111
rect	294	111	295	112
rect	294	112	295	113
rect	294	113	295	114
rect	294	114	295	115
rect	294	116	295	117
rect	294	117	295	118
rect	294	118	295	119
rect	294	119	295	120
rect	294	120	295	121
rect	294	121	295	122
rect	294	122	295	123
rect	294	123	295	124
rect	294	125	295	126
rect	294	126	295	127
rect	294	127	295	128
rect	294	128	295	129
rect	294	129	295	130
rect	294	130	295	131
rect	294	131	295	132
rect	294	132	295	133
rect	294	133	295	134
rect	294	134	295	135
rect	294	135	295	136
rect	294	137	295	138
rect	294	138	295	139
rect	294	140	295	141
rect	294	141	295	142
rect	294	142	295	143
rect	294	143	295	144
rect	294	144	295	145
rect	294	145	295	146
rect	294	146	295	147
rect	294	147	295	148
rect	294	148	295	149
rect	294	149	295	150
rect	294	150	295	151
rect	294	152	295	153
rect	294	153	295	154
rect	294	154	295	155
rect	294	155	295	156
rect	294	156	295	157
rect	294	157	295	158
rect	294	158	295	159
rect	294	159	295	160
rect	294	161	295	162
rect	294	162	295	163
rect	294	163	295	164
rect	294	164	295	165
rect	294	165	295	166
rect	294	167	295	168
rect	294	168	295	169
rect	294	170	295	171
rect	294	171	295	172
rect	294	172	295	173
rect	294	173	295	174
rect	294	174	295	175
rect	294	175	295	176
rect	294	176	295	177
rect	294	177	295	178
rect	294	178	295	179
rect	294	179	295	180
rect	294	180	295	181
rect	294	181	295	182
rect	294	182	295	183
rect	294	183	295	184
rect	294	184	295	185
rect	294	185	295	186
rect	294	186	295	187
rect	294	187	295	188
rect	294	188	295	189
rect	294	189	295	190
rect	294	190	295	191
rect	294	191	295	192
rect	294	192	295	193
rect	294	193	295	194
rect	294	194	295	195
rect	297	0	298	1
rect	297	1	298	2
rect	297	2	298	3
rect	297	3	298	4
rect	297	4	298	5
rect	297	5	298	6
rect	297	6	298	7
rect	297	8	298	9
rect	297	9	298	10
rect	297	10	298	11
rect	297	11	298	12
rect	297	12	298	13
rect	297	14	298	15
rect	297	15	298	16
rect	297	16	298	17
rect	297	17	298	18
rect	297	18	298	19
rect	297	19	298	20
rect	297	20	298	21
rect	297	21	298	22
rect	297	22	298	23
rect	297	23	298	24
rect	297	24	298	25
rect	297	25	298	26
rect	297	26	298	27
rect	297	27	298	28
rect	297	29	298	30
rect	297	30	298	31
rect	297	32	298	33
rect	297	33	298	34
rect	297	34	298	35
rect	297	35	298	36
rect	297	36	298	37
rect	297	37	298	38
rect	297	38	298	39
rect	297	39	298	40
rect	297	40	298	41
rect	297	41	298	42
rect	297	42	298	43
rect	297	43	298	44
rect	297	44	298	45
rect	297	45	298	46
rect	297	46	298	47
rect	297	47	298	48
rect	297	48	298	49
rect	297	49	298	50
rect	297	50	298	51
rect	297	51	298	52
rect	297	52	298	53
rect	297	53	298	54
rect	297	54	298	55
rect	297	55	298	56
rect	297	56	298	57
rect	297	57	298	58
rect	297	58	298	59
rect	297	59	298	60
rect	297	60	298	61
rect	297	61	298	62
rect	297	62	298	63
rect	297	63	298	64
rect	297	65	298	66
rect	297	66	298	67
rect	297	67	298	68
rect	297	68	298	69
rect	297	69	298	70
rect	297	70	298	71
rect	297	71	298	72
rect	297	72	298	73
rect	297	73	298	74
rect	297	74	298	75
rect	297	75	298	76
rect	297	76	298	77
rect	297	77	298	78
rect	297	78	298	79
rect	297	79	298	80
rect	297	80	298	81
rect	297	81	298	82
rect	297	82	298	83
rect	297	83	298	84
rect	297	84	298	85
rect	297	86	298	87
rect	297	87	298	88
rect	297	88	298	89
rect	297	89	298	90
rect	297	90	298	91
rect	297	91	298	92
rect	297	92	298	93
rect	297	93	298	94
rect	297	94	298	95
rect	297	95	298	96
rect	297	96	298	97
rect	297	97	298	98
rect	297	98	298	99
rect	297	99	298	100
rect	297	100	298	101
rect	297	101	298	102
rect	297	102	298	103
rect	297	103	298	104
rect	297	104	298	105
rect	297	105	298	106
rect	297	106	298	107
rect	297	107	298	108
rect	297	108	298	109
rect	297	109	298	110
rect	297	110	298	111
rect	297	111	298	112
rect	297	112	298	113
rect	297	113	298	114
rect	297	114	298	115
rect	297	116	298	117
rect	297	117	298	118
rect	297	118	298	119
rect	297	119	298	120
rect	297	120	298	121
rect	297	121	298	122
rect	297	122	298	123
rect	297	123	298	124
rect	297	125	298	126
rect	297	126	298	127
rect	297	127	298	128
rect	297	128	298	129
rect	297	129	298	130
rect	297	130	298	131
rect	297	131	298	132
rect	297	132	298	133
rect	297	133	298	134
rect	297	134	298	135
rect	297	135	298	136
rect	297	137	298	138
rect	297	138	298	139
rect	297	140	298	141
rect	297	141	298	142
rect	297	142	298	143
rect	297	143	298	144
rect	297	144	298	145
rect	297	145	298	146
rect	297	146	298	147
rect	297	147	298	148
rect	297	148	298	149
rect	297	149	298	150
rect	297	150	298	151
rect	297	151	298	152
rect	297	152	298	153
rect	297	153	298	154
rect	297	154	298	155
rect	297	155	298	156
rect	297	156	298	157
rect	297	157	298	158
rect	297	158	298	159
rect	297	159	298	160
rect	297	160	298	161
rect	297	161	298	162
rect	297	162	298	163
rect	297	163	298	164
rect	297	164	298	165
rect	297	165	298	166
rect	297	167	298	168
rect	297	168	298	169
rect	297	169	298	170
rect	297	170	298	171
rect	297	171	298	172
rect	297	172	298	173
rect	297	173	298	174
rect	297	174	298	175
rect	297	175	298	176
rect	297	176	298	177
rect	297	177	298	178
rect	297	178	298	179
rect	297	179	298	180
rect	297	180	298	181
rect	297	181	298	182
rect	297	182	298	183
rect	297	183	298	184
rect	297	184	298	185
rect	297	185	298	186
rect	297	186	298	187
rect	297	187	298	188
rect	297	188	298	189
rect	297	189	298	190
rect	297	190	298	191
rect	297	191	298	192
rect	297	192	298	193
rect	297	193	298	194
rect	297	194	298	195
rect	299	0	300	1
rect	299	1	300	2
rect	299	2	300	3
rect	299	3	300	4
rect	299	4	300	5
rect	299	5	300	6
rect	299	6	300	7
rect	299	8	300	9
rect	299	9	300	10
rect	299	10	300	11
rect	299	11	300	12
rect	299	12	300	13
rect	299	14	300	15
rect	299	15	300	16
rect	299	16	300	17
rect	299	17	300	18
rect	299	18	300	19
rect	299	19	300	20
rect	299	20	300	21
rect	299	21	300	22
rect	299	22	300	23
rect	299	23	300	24
rect	299	24	300	25
rect	299	25	300	26
rect	299	26	300	27
rect	299	27	300	28
rect	299	29	300	30
rect	299	30	300	31
rect	299	32	300	33
rect	299	33	300	34
rect	299	34	300	35
rect	299	35	300	36
rect	299	36	300	37
rect	299	37	300	38
rect	299	38	300	39
rect	299	39	300	40
rect	299	40	300	41
rect	299	41	300	42
rect	299	42	300	43
rect	299	43	300	44
rect	299	44	300	45
rect	299	45	300	46
rect	299	46	300	47
rect	299	47	300	48
rect	299	48	300	49
rect	299	49	300	50
rect	299	50	300	51
rect	299	51	300	52
rect	299	52	300	53
rect	299	53	300	54
rect	299	54	300	55
rect	299	55	300	56
rect	299	56	300	57
rect	299	57	300	58
rect	299	58	300	59
rect	299	59	300	60
rect	299	60	300	61
rect	299	61	300	62
rect	299	62	300	63
rect	299	63	300	64
rect	299	65	300	66
rect	299	66	300	67
rect	299	67	300	68
rect	299	68	300	69
rect	299	69	300	70
rect	299	70	300	71
rect	299	71	300	72
rect	299	72	300	73
rect	299	73	300	74
rect	299	74	300	75
rect	299	75	300	76
rect	299	76	300	77
rect	299	77	300	78
rect	299	78	300	79
rect	299	79	300	80
rect	299	80	300	81
rect	299	81	300	82
rect	299	82	300	83
rect	299	83	300	84
rect	299	84	300	85
rect	299	86	300	87
rect	299	87	300	88
rect	299	88	300	89
rect	299	89	300	90
rect	299	90	300	91
rect	299	91	300	92
rect	299	92	300	93
rect	299	93	300	94
rect	299	94	300	95
rect	299	95	300	96
rect	299	96	300	97
rect	299	97	300	98
rect	299	98	300	99
rect	299	99	300	100
rect	299	100	300	101
rect	299	101	300	102
rect	299	102	300	103
rect	299	103	300	104
rect	299	104	300	105
rect	299	105	300	106
rect	299	106	300	107
rect	299	107	300	108
rect	299	108	300	109
rect	299	109	300	110
rect	299	110	300	111
rect	299	111	300	112
rect	299	112	300	113
rect	299	113	300	114
rect	299	114	300	115
rect	299	116	300	117
rect	299	117	300	118
rect	299	118	300	119
rect	299	119	300	120
rect	299	120	300	121
rect	299	121	300	122
rect	299	122	300	123
rect	299	123	300	124
rect	299	125	300	126
rect	299	126	300	127
rect	299	127	300	128
rect	299	128	300	129
rect	299	129	300	130
rect	299	130	300	131
rect	299	131	300	132
rect	299	132	300	133
rect	299	133	300	134
rect	299	134	300	135
rect	299	135	300	136
rect	299	137	300	138
rect	299	138	300	139
rect	299	140	300	141
rect	299	141	300	142
rect	299	142	300	143
rect	299	143	300	144
rect	299	144	300	145
rect	299	145	300	146
rect	299	146	300	147
rect	299	147	300	148
rect	299	148	300	149
rect	299	149	300	150
rect	299	150	300	151
rect	299	151	300	152
rect	299	152	300	153
rect	299	153	300	154
rect	299	154	300	155
rect	299	155	300	156
rect	299	156	300	157
rect	299	157	300	158
rect	299	158	300	159
rect	299	159	300	160
rect	299	160	300	161
rect	299	161	300	162
rect	299	162	300	163
rect	299	163	300	164
rect	299	164	300	165
rect	299	165	300	166
rect	299	167	300	168
rect	300	0	301	1
rect	300	1	301	2
rect	300	2	301	3
rect	300	3	301	4
rect	300	4	301	5
rect	300	5	301	6
rect	300	6	301	7
rect	300	8	301	9
rect	300	9	301	10
rect	300	10	301	11
rect	300	11	301	12
rect	300	12	301	13
rect	300	14	301	15
rect	300	15	301	16
rect	300	16	301	17
rect	300	17	301	18
rect	300	18	301	19
rect	300	19	301	20
rect	300	20	301	21
rect	300	21	301	22
rect	300	22	301	23
rect	300	23	301	24
rect	300	24	301	25
rect	300	25	301	26
rect	300	26	301	27
rect	300	27	301	28
rect	300	29	301	30
rect	300	30	301	31
rect	300	32	301	33
rect	300	33	301	34
rect	300	34	301	35
rect	300	35	301	36
rect	300	36	301	37
rect	300	37	301	38
rect	300	38	301	39
rect	300	39	301	40
rect	300	40	301	41
rect	300	41	301	42
rect	300	42	301	43
rect	300	43	301	44
rect	300	44	301	45
rect	300	45	301	46
rect	300	46	301	47
rect	300	47	301	48
rect	300	48	301	49
rect	300	49	301	50
rect	300	50	301	51
rect	300	51	301	52
rect	300	52	301	53
rect	300	53	301	54
rect	300	54	301	55
rect	300	55	301	56
rect	300	56	301	57
rect	300	57	301	58
rect	300	58	301	59
rect	300	59	301	60
rect	300	60	301	61
rect	300	61	301	62
rect	300	62	301	63
rect	300	63	301	64
rect	300	65	301	66
rect	300	66	301	67
rect	300	67	301	68
rect	300	68	301	69
rect	300	69	301	70
rect	300	70	301	71
rect	300	71	301	72
rect	300	72	301	73
rect	300	73	301	74
rect	300	74	301	75
rect	300	75	301	76
rect	300	76	301	77
rect	300	77	301	78
rect	300	78	301	79
rect	300	79	301	80
rect	300	80	301	81
rect	300	81	301	82
rect	300	82	301	83
rect	300	83	301	84
rect	300	84	301	85
rect	300	86	301	87
rect	300	87	301	88
rect	300	88	301	89
rect	300	89	301	90
rect	300	90	301	91
rect	300	91	301	92
rect	300	92	301	93
rect	300	93	301	94
rect	300	94	301	95
rect	300	95	301	96
rect	300	96	301	97
rect	300	97	301	98
rect	300	98	301	99
rect	300	99	301	100
rect	300	100	301	101
rect	300	101	301	102
rect	300	102	301	103
rect	300	103	301	104
rect	300	104	301	105
rect	300	105	301	106
rect	300	106	301	107
rect	300	107	301	108
rect	300	108	301	109
rect	300	109	301	110
rect	300	110	301	111
rect	300	111	301	112
rect	300	112	301	113
rect	300	113	301	114
rect	300	114	301	115
rect	300	116	301	117
rect	300	117	301	118
rect	300	118	301	119
rect	300	119	301	120
rect	300	120	301	121
rect	300	121	301	122
rect	300	122	301	123
rect	300	123	301	124
rect	300	125	301	126
rect	300	126	301	127
rect	300	127	301	128
rect	300	128	301	129
rect	300	129	301	130
rect	300	130	301	131
rect	300	131	301	132
rect	300	132	301	133
rect	300	133	301	134
rect	300	134	301	135
rect	300	135	301	136
rect	300	137	301	138
rect	300	138	301	139
rect	300	140	301	141
rect	300	141	301	142
rect	300	142	301	143
rect	300	143	301	144
rect	300	144	301	145
rect	300	145	301	146
rect	300	146	301	147
rect	300	147	301	148
rect	300	148	301	149
rect	300	149	301	150
rect	300	150	301	151
rect	300	151	301	152
rect	300	152	301	153
rect	300	153	301	154
rect	300	154	301	155
rect	300	155	301	156
rect	300	156	301	157
rect	300	157	301	158
rect	300	158	301	159
rect	300	159	301	160
rect	300	160	301	161
rect	300	161	301	162
rect	300	162	301	163
rect	300	163	301	164
rect	300	164	301	165
rect	300	165	301	166
rect	300	167	301	168
rect	301	0	302	1
rect	301	1	302	2
rect	301	2	302	3
rect	301	3	302	4
rect	301	4	302	5
rect	301	5	302	6
rect	301	6	302	7
rect	301	8	302	9
rect	301	9	302	10
rect	301	10	302	11
rect	301	11	302	12
rect	301	12	302	13
rect	301	14	302	15
rect	301	15	302	16
rect	301	16	302	17
rect	301	17	302	18
rect	301	18	302	19
rect	301	19	302	20
rect	301	20	302	21
rect	301	21	302	22
rect	301	22	302	23
rect	301	23	302	24
rect	301	24	302	25
rect	301	25	302	26
rect	301	26	302	27
rect	301	27	302	28
rect	301	29	302	30
rect	301	30	302	31
rect	301	32	302	33
rect	301	33	302	34
rect	301	34	302	35
rect	301	35	302	36
rect	301	36	302	37
rect	301	37	302	38
rect	301	38	302	39
rect	301	39	302	40
rect	301	40	302	41
rect	301	41	302	42
rect	301	42	302	43
rect	301	43	302	44
rect	301	44	302	45
rect	301	45	302	46
rect	301	46	302	47
rect	301	47	302	48
rect	301	48	302	49
rect	301	49	302	50
rect	301	50	302	51
rect	301	51	302	52
rect	301	52	302	53
rect	301	53	302	54
rect	301	54	302	55
rect	301	55	302	56
rect	301	56	302	57
rect	301	57	302	58
rect	301	58	302	59
rect	301	59	302	60
rect	301	60	302	61
rect	301	61	302	62
rect	301	62	302	63
rect	301	63	302	64
rect	301	65	302	66
rect	301	66	302	67
rect	301	67	302	68
rect	301	68	302	69
rect	301	69	302	70
rect	301	70	302	71
rect	301	71	302	72
rect	301	72	302	73
rect	301	73	302	74
rect	301	74	302	75
rect	301	75	302	76
rect	301	76	302	77
rect	301	77	302	78
rect	301	78	302	79
rect	301	79	302	80
rect	301	80	302	81
rect	301	81	302	82
rect	301	82	302	83
rect	301	83	302	84
rect	301	84	302	85
rect	301	86	302	87
rect	301	87	302	88
rect	301	88	302	89
rect	301	89	302	90
rect	301	90	302	91
rect	301	91	302	92
rect	301	92	302	93
rect	301	93	302	94
rect	301	94	302	95
rect	301	95	302	96
rect	301	96	302	97
rect	301	97	302	98
rect	301	98	302	99
rect	301	99	302	100
rect	301	100	302	101
rect	301	101	302	102
rect	301	102	302	103
rect	301	103	302	104
rect	301	104	302	105
rect	301	105	302	106
rect	301	106	302	107
rect	301	107	302	108
rect	301	108	302	109
rect	301	109	302	110
rect	301	110	302	111
rect	301	111	302	112
rect	301	112	302	113
rect	301	113	302	114
rect	301	114	302	115
rect	301	116	302	117
rect	301	117	302	118
rect	301	118	302	119
rect	301	119	302	120
rect	301	120	302	121
rect	301	121	302	122
rect	301	122	302	123
rect	301	123	302	124
rect	301	125	302	126
rect	301	126	302	127
rect	301	127	302	128
rect	301	128	302	129
rect	301	129	302	130
rect	301	130	302	131
rect	301	131	302	132
rect	301	132	302	133
rect	301	133	302	134
rect	301	134	302	135
rect	301	135	302	136
rect	301	137	302	138
rect	301	138	302	139
rect	301	140	302	141
rect	301	141	302	142
rect	301	142	302	143
rect	301	143	302	144
rect	301	144	302	145
rect	301	145	302	146
rect	301	146	302	147
rect	301	147	302	148
rect	301	148	302	149
rect	301	149	302	150
rect	301	150	302	151
rect	301	151	302	152
rect	301	152	302	153
rect	301	153	302	154
rect	301	154	302	155
rect	301	155	302	156
rect	301	156	302	157
rect	301	157	302	158
rect	301	158	302	159
rect	301	159	302	160
rect	301	160	302	161
rect	301	161	302	162
rect	301	162	302	163
rect	301	163	302	164
rect	301	164	302	165
rect	301	165	302	166
rect	301	167	302	168
rect	302	0	303	1
rect	302	1	303	2
rect	302	2	303	3
rect	302	3	303	4
rect	302	4	303	5
rect	302	5	303	6
rect	302	6	303	7
rect	302	8	303	9
rect	302	9	303	10
rect	302	10	303	11
rect	302	11	303	12
rect	302	12	303	13
rect	302	14	303	15
rect	302	15	303	16
rect	302	16	303	17
rect	302	17	303	18
rect	302	18	303	19
rect	302	19	303	20
rect	302	20	303	21
rect	302	21	303	22
rect	302	22	303	23
rect	302	23	303	24
rect	302	24	303	25
rect	302	25	303	26
rect	302	26	303	27
rect	302	27	303	28
rect	302	29	303	30
rect	302	30	303	31
rect	302	32	303	33
rect	302	33	303	34
rect	302	34	303	35
rect	302	35	303	36
rect	302	36	303	37
rect	302	37	303	38
rect	302	38	303	39
rect	302	39	303	40
rect	302	40	303	41
rect	302	41	303	42
rect	302	42	303	43
rect	302	43	303	44
rect	302	44	303	45
rect	302	45	303	46
rect	302	46	303	47
rect	302	47	303	48
rect	302	48	303	49
rect	302	49	303	50
rect	302	50	303	51
rect	302	51	303	52
rect	302	52	303	53
rect	302	53	303	54
rect	302	54	303	55
rect	302	55	303	56
rect	302	56	303	57
rect	302	57	303	58
rect	302	58	303	59
rect	302	59	303	60
rect	302	60	303	61
rect	302	61	303	62
rect	302	62	303	63
rect	302	63	303	64
rect	302	65	303	66
rect	302	66	303	67
rect	302	67	303	68
rect	302	68	303	69
rect	302	69	303	70
rect	302	70	303	71
rect	302	71	303	72
rect	302	72	303	73
rect	302	73	303	74
rect	302	74	303	75
rect	302	75	303	76
rect	302	76	303	77
rect	302	77	303	78
rect	302	78	303	79
rect	302	79	303	80
rect	302	80	303	81
rect	302	81	303	82
rect	302	82	303	83
rect	302	83	303	84
rect	302	84	303	85
rect	302	86	303	87
rect	302	87	303	88
rect	302	88	303	89
rect	302	89	303	90
rect	302	90	303	91
rect	302	91	303	92
rect	302	92	303	93
rect	302	93	303	94
rect	302	94	303	95
rect	302	95	303	96
rect	302	96	303	97
rect	302	97	303	98
rect	302	98	303	99
rect	302	99	303	100
rect	302	100	303	101
rect	302	101	303	102
rect	302	102	303	103
rect	302	103	303	104
rect	302	104	303	105
rect	302	105	303	106
rect	302	106	303	107
rect	302	107	303	108
rect	302	108	303	109
rect	302	109	303	110
rect	302	110	303	111
rect	302	111	303	112
rect	302	112	303	113
rect	302	113	303	114
rect	302	114	303	115
rect	302	116	303	117
rect	302	117	303	118
rect	302	118	303	119
rect	302	119	303	120
rect	302	120	303	121
rect	302	121	303	122
rect	302	122	303	123
rect	302	123	303	124
rect	302	125	303	126
rect	302	126	303	127
rect	302	127	303	128
rect	302	128	303	129
rect	302	129	303	130
rect	302	130	303	131
rect	302	131	303	132
rect	302	132	303	133
rect	302	133	303	134
rect	302	134	303	135
rect	302	135	303	136
rect	302	137	303	138
rect	302	138	303	139
rect	302	140	303	141
rect	302	141	303	142
rect	302	142	303	143
rect	302	143	303	144
rect	302	144	303	145
rect	302	145	303	146
rect	302	146	303	147
rect	302	147	303	148
rect	302	148	303	149
rect	302	149	303	150
rect	302	150	303	151
rect	302	151	303	152
rect	302	152	303	153
rect	302	153	303	154
rect	302	154	303	155
rect	302	155	303	156
rect	302	156	303	157
rect	302	157	303	158
rect	302	158	303	159
rect	302	159	303	160
rect	302	160	303	161
rect	302	161	303	162
rect	302	162	303	163
rect	302	163	303	164
rect	302	164	303	165
rect	302	165	303	166
rect	302	167	303	168
rect	303	0	304	1
rect	303	1	304	2
rect	303	2	304	3
rect	303	3	304	4
rect	303	4	304	5
rect	303	5	304	6
rect	303	6	304	7
rect	303	7	304	8
rect	303	8	304	9
rect	303	9	304	10
rect	303	10	304	11
rect	303	11	304	12
rect	303	12	304	13
rect	303	13	304	14
rect	303	14	304	15
rect	303	15	304	16
rect	303	16	304	17
rect	303	17	304	18
rect	303	18	304	19
rect	303	19	304	20
rect	303	20	304	21
rect	303	21	304	22
rect	303	22	304	23
rect	303	23	304	24
rect	303	24	304	25
rect	303	25	304	26
rect	303	26	304	27
rect	303	27	304	28
rect	303	28	304	29
rect	303	29	304	30
rect	303	30	304	31
rect	303	31	304	32
rect	303	32	304	33
rect	303	33	304	34
rect	303	34	304	35
rect	303	35	304	36
rect	303	36	304	37
rect	303	37	304	38
rect	303	38	304	39
rect	303	39	304	40
rect	303	40	304	41
rect	303	41	304	42
rect	303	42	304	43
rect	303	43	304	44
rect	303	44	304	45
rect	303	45	304	46
rect	303	46	304	47
rect	303	47	304	48
rect	303	48	304	49
rect	303	49	304	50
rect	303	50	304	51
rect	303	51	304	52
rect	303	52	304	53
rect	303	53	304	54
rect	303	54	304	55
rect	303	55	304	56
rect	303	56	304	57
rect	303	57	304	58
rect	303	58	304	59
rect	303	59	304	60
rect	303	60	304	61
rect	303	61	304	62
rect	303	62	304	63
rect	303	63	304	64
rect	303	64	304	65
rect	303	65	304	66
rect	303	66	304	67
rect	303	67	304	68
rect	303	68	304	69
rect	303	69	304	70
rect	303	70	304	71
rect	303	71	304	72
rect	303	72	304	73
rect	303	73	304	74
rect	303	74	304	75
rect	303	75	304	76
rect	303	76	304	77
rect	303	77	304	78
rect	303	78	304	79
rect	303	79	304	80
rect	303	80	304	81
rect	303	81	304	82
rect	303	82	304	83
rect	303	83	304	84
rect	303	84	304	85
rect	303	85	304	86
rect	303	86	304	87
rect	303	87	304	88
rect	303	88	304	89
rect	303	89	304	90
rect	303	90	304	91
rect	303	91	304	92
rect	303	92	304	93
rect	303	93	304	94
rect	303	94	304	95
rect	303	95	304	96
rect	303	96	304	97
rect	303	97	304	98
rect	303	98	304	99
rect	303	99	304	100
rect	303	100	304	101
rect	303	101	304	102
rect	303	102	304	103
rect	303	103	304	104
rect	303	104	304	105
rect	303	105	304	106
rect	303	106	304	107
rect	303	107	304	108
rect	303	108	304	109
rect	303	109	304	110
rect	303	110	304	111
rect	303	111	304	112
rect	303	112	304	113
rect	303	113	304	114
rect	303	114	304	115
rect	303	115	304	116
rect	303	116	304	117
rect	303	117	304	118
rect	303	118	304	119
rect	303	119	304	120
rect	303	120	304	121
rect	303	121	304	122
rect	303	122	304	123
rect	303	123	304	124
rect	303	124	304	125
rect	303	125	304	126
rect	303	126	304	127
rect	303	127	304	128
rect	303	128	304	129
rect	303	129	304	130
rect	303	130	304	131
rect	303	131	304	132
rect	303	132	304	133
rect	303	133	304	134
rect	303	134	304	135
rect	303	135	304	136
rect	303	136	304	137
rect	303	137	304	138
rect	303	138	304	139
rect	303	139	304	140
rect	303	140	304	141
rect	303	141	304	142
rect	303	142	304	143
rect	303	143	304	144
rect	303	144	304	145
rect	303	145	304	146
rect	303	146	304	147
rect	303	147	304	148
rect	303	148	304	149
rect	303	149	304	150
rect	303	150	304	151
rect	303	151	304	152
rect	303	152	304	153
rect	303	153	304	154
rect	303	154	304	155
rect	303	155	304	156
rect	303	156	304	157
rect	303	157	304	158
rect	303	158	304	159
rect	303	159	304	160
rect	303	160	304	161
rect	303	161	304	162
rect	303	162	304	163
rect	303	163	304	164
rect	303	164	304	165
rect	303	165	304	166
rect	303	166	304	167
rect	303	167	304	168
rect	308	0	309	1
rect	308	1	309	2
rect	308	2	309	3
rect	308	3	309	4
rect	308	4	309	5
rect	308	5	309	6
rect	308	6	309	7
rect	308	7	309	8
rect	308	8	309	9
rect	308	9	309	10
rect	308	10	309	11
rect	308	11	309	12
rect	308	12	309	13
rect	308	13	309	14
rect	308	14	309	15
rect	308	15	309	16
rect	308	16	309	17
rect	308	17	309	18
rect	308	18	309	19
rect	308	19	309	20
rect	308	20	309	21
rect	308	21	309	22
rect	308	22	309	23
rect	308	23	309	24
rect	308	24	309	25
rect	308	25	309	26
rect	308	26	309	27
rect	308	27	309	28
rect	308	28	309	29
rect	308	29	309	30
rect	308	30	309	31
rect	308	31	309	32
rect	308	32	309	33
rect	308	33	309	34
rect	308	34	309	35
rect	308	35	309	36
rect	308	36	309	37
rect	308	37	309	38
rect	308	38	309	39
rect	308	39	309	40
rect	308	40	309	41
rect	308	41	309	42
rect	308	42	309	43
rect	308	43	309	44
rect	308	44	309	45
rect	308	45	309	46
rect	308	46	309	47
rect	308	47	309	48
rect	308	48	309	49
rect	308	49	309	50
rect	308	50	309	51
rect	308	51	309	52
rect	308	52	309	53
rect	308	53	309	54
rect	308	54	309	55
rect	308	55	309	56
rect	308	56	309	57
rect	308	57	309	58
rect	308	58	309	59
rect	308	59	309	60
rect	308	60	309	61
rect	308	61	309	62
rect	308	62	309	63
rect	308	63	309	64
rect	308	64	309	65
rect	308	65	309	66
rect	308	66	309	67
rect	308	67	309	68
rect	308	68	309	69
rect	308	69	309	70
rect	308	70	309	71
rect	308	71	309	72
rect	308	72	309	73
rect	308	73	309	74
rect	308	74	309	75
rect	308	75	309	76
rect	308	76	309	77
rect	308	77	309	78
rect	308	78	309	79
rect	308	79	309	80
rect	308	80	309	81
rect	308	81	309	82
rect	308	82	309	83
rect	308	83	309	84
rect	308	84	309	85
rect	308	85	309	86
rect	308	86	309	87
rect	308	87	309	88
rect	308	88	309	89
rect	308	89	309	90
rect	308	90	309	91
rect	308	91	309	92
rect	308	92	309	93
rect	308	93	309	94
rect	308	94	309	95
rect	308	95	309	96
rect	308	96	309	97
rect	308	97	309	98
rect	308	98	309	99
rect	308	99	309	100
rect	308	100	309	101
rect	308	101	309	102
rect	308	102	309	103
rect	308	103	309	104
rect	308	104	309	105
rect	308	105	309	106
rect	308	106	309	107
rect	308	107	309	108
rect	308	108	309	109
rect	308	109	309	110
rect	308	110	309	111
rect	308	111	309	112
rect	308	112	309	113
rect	308	113	309	114
rect	308	114	309	115
rect	308	115	309	116
rect	308	116	309	117
rect	308	117	309	118
rect	308	118	309	119
rect	308	119	309	120
rect	308	120	309	121
rect	308	121	309	122
rect	308	122	309	123
rect	308	123	309	124
rect	308	124	309	125
rect	308	125	309	126
rect	308	126	309	127
rect	308	127	309	128
rect	308	128	309	129
rect	308	129	309	130
rect	308	130	309	131
rect	308	131	309	132
rect	308	132	309	133
rect	308	133	309	134
rect	308	134	309	135
rect	308	135	309	136
rect	308	136	309	137
rect	308	137	309	138
rect	308	138	309	139
rect	308	139	309	140
rect	308	140	309	141
rect	308	141	309	142
rect	308	142	309	143
rect	308	143	309	144
rect	308	144	309	145
rect	308	145	309	146
rect	308	146	309	147
rect	308	147	309	148
rect	308	148	309	149
rect	308	149	309	150
rect	308	150	309	151
rect	308	151	309	152
rect	308	152	309	153
rect	308	153	309	154
rect	308	154	309	155
rect	308	155	309	156
rect	308	156	309	157
rect	308	157	309	158
rect	308	158	309	159
rect	308	159	309	160
rect	308	160	309	161
rect	308	161	309	162
rect	308	162	309	163
rect	308	163	309	164
rect	308	164	309	165
rect	308	165	309	166
rect	308	166	309	167
rect	308	167	309	168
<< metal1 >>
rect	0	122	1	123
rect	0	123	1	124
rect	0	124	1	125
rect	0	125	1	126
rect	0	126	1	127
rect	0	127	1	128
rect	0	128	1	129
rect	0	129	1	130
rect	0	130	1	131
rect	0	131	1	132
rect	0	132	1	133
rect	0	133	1	134
rect	0	134	1	135
rect	0	135	1	136
rect	0	136	1	137
rect	0	137	1	138
rect	0	138	1	139
rect	0	139	1	140
rect	0	140	1	141
rect	0	141	1	142
rect	0	142	1	143
rect	0	143	1	144
rect	0	144	1	145
rect	0	145	1	146
rect	0	146	1	147
rect	0	147	1	148
rect	0	148	1	149
rect	0	149	1	150
rect	0	150	1	151
rect	0	151	1	152
rect	0	152	1	153
rect	0	153	1	154
rect	0	154	1	155
rect	0	155	1	156
rect	0	156	1	157
rect	0	157	1	158
rect	0	158	1	159
rect	0	159	1	160
rect	0	160	1	161
rect	0	161	1	162
rect	0	162	1	163
rect	0	163	1	164
rect	0	164	1	165
rect	0	165	1	166
rect	0	166	1	167
rect	0	167	1	168
rect	0	168	1	169
rect	0	169	1	170
rect	0	170	1	171
rect	0	171	1	172
rect	2	53	3	54
rect	2	54	3	55
rect	2	55	3	56
rect	2	56	3	57
rect	2	57	3	58
rect	2	110	3	111
rect	2	111	3	112
rect	2	112	3	113
rect	2	113	3	114
rect	2	114	3	115
rect	2	119	3	120
rect	2	120	3	121
rect	2	122	3	123
rect	2	123	3	124
rect	2	137	3	138
rect	2	138	3	139
rect	2	139	3	140
rect	2	140	3	141
rect	2	141	3	142
rect	2	142	3	143
rect	2	143	3	144
rect	2	144	3	145
rect	4	8	5	9
rect	4	9	5	10
rect	4	10	5	11
rect	4	11	5	12
rect	4	12	5	13
rect	4	13	5	14
rect	4	14	5	15
rect	4	15	5	16
rect	4	16	5	17
rect	4	17	5	18
rect	4	18	5	19
rect	4	19	5	20
rect	4	20	5	21
rect	4	21	5	22
rect	4	22	5	23
rect	4	23	5	24
rect	4	24	5	25
rect	4	25	5	26
rect	4	26	5	27
rect	4	27	5	28
rect	4	28	5	29
rect	4	29	5	30
rect	4	30	5	31
rect	4	31	5	32
rect	4	32	5	33
rect	4	33	5	34
rect	4	34	5	35
rect	4	35	5	36
rect	4	36	5	37
rect	4	37	5	38
rect	4	38	5	39
rect	4	39	5	40
rect	4	40	5	41
rect	4	41	5	42
rect	4	42	5	43
rect	4	43	5	44
rect	4	44	5	45
rect	4	45	5	46
rect	4	46	5	47
rect	4	47	5	48
rect	4	48	5	49
rect	4	49	5	50
rect	4	50	5	51
rect	4	51	5	52
rect	4	53	5	54
rect	4	54	5	55
rect	4	55	5	56
rect	4	56	5	57
rect	4	57	5	58
rect	4	59	5	60
rect	4	60	5	61
rect	4	61	5	62
rect	4	62	5	63
rect	4	63	5	64
rect	4	64	5	65
rect	4	65	5	66
rect	4	66	5	67
rect	4	67	5	68
rect	4	68	5	69
rect	4	69	5	70
rect	4	70	5	71
rect	4	71	5	72
rect	4	72	5	73
rect	4	73	5	74
rect	4	74	5	75
rect	4	75	5	76
rect	4	76	5	77
rect	4	77	5	78
rect	4	78	5	79
rect	4	86	5	87
rect	4	87	5	88
rect	4	88	5	89
rect	4	89	5	90
rect	4	90	5	91
rect	4	107	5	108
rect	4	108	5	109
rect	4	110	5	111
rect	4	111	5	112
rect	4	112	5	113
rect	4	113	5	114
rect	4	114	5	115
rect	4	116	5	117
rect	4	117	5	118
rect	4	119	5	120
rect	4	120	5	121
rect	4	122	5	123
rect	4	123	5	124
rect	4	125	5	126
rect	4	126	5	127
rect	4	127	5	128
rect	4	128	5	129
rect	4	129	5	130
rect	4	130	5	131
rect	4	131	5	132
rect	4	132	5	133
rect	4	133	5	134
rect	4	134	5	135
rect	4	135	5	136
rect	4	137	5	138
rect	4	138	5	139
rect	4	139	5	140
rect	4	140	5	141
rect	4	141	5	142
rect	18	119	19	120
rect	18	120	19	121
rect	18	122	19	123
rect	18	123	19	124
rect	18	125	19	126
rect	18	126	19	127
rect	18	134	19	135
rect	18	135	19	136
rect	18	137	19	138
rect	18	138	19	139
rect	18	164	19	165
rect	18	165	19	166
rect	20	11	21	12
rect	20	12	21	13
rect	20	17	21	18
rect	20	18	21	19
rect	20	20	21	21
rect	20	21	21	22
rect	20	53	21	54
rect	20	54	21	55
rect	20	77	21	78
rect	20	78	21	79
rect	20	80	21	81
rect	20	81	21	82
rect	20	83	21	84
rect	20	84	21	85
rect	20	86	21	87
rect	20	87	21	88
rect	20	89	21	90
rect	20	90	21	91
rect	20	92	21	93
rect	20	93	21	94
rect	20	95	21	96
rect	20	96	21	97
rect	20	98	21	99
rect	20	99	21	100
rect	20	101	21	102
rect	20	102	21	103
rect	20	104	21	105
rect	20	105	21	106
rect	20	107	21	108
rect	20	108	21	109
rect	20	110	21	111
rect	20	111	21	112
rect	20	113	21	114
rect	20	114	21	115
rect	20	116	21	117
rect	20	117	21	118
rect	20	119	21	120
rect	20	120	21	121
rect	20	122	21	123
rect	20	123	21	124
rect	20	125	21	126
rect	20	126	21	127
rect	20	128	21	129
rect	20	129	21	130
rect	20	131	21	132
rect	20	132	21	133
rect	20	134	21	135
rect	20	135	21	136
rect	20	137	21	138
rect	20	138	21	139
rect	20	140	21	141
rect	20	141	21	142
rect	20	143	21	144
rect	20	144	21	145
rect	20	146	21	147
rect	20	147	21	148
rect	20	149	21	150
rect	20	150	21	151
rect	20	152	21	153
rect	20	153	21	154
rect	20	155	21	156
rect	20	156	21	157
rect	20	158	21	159
rect	20	159	21	160
rect	20	161	21	162
rect	20	162	21	163
rect	20	164	21	165
rect	20	165	21	166
rect	20	167	21	168
rect	20	168	21	169
rect	20	170	21	171
rect	20	171	21	172
rect	20	173	21	174
rect	20	174	21	175
rect	20	188	21	189
rect	20	189	21	190
rect	29	113	30	114
rect	29	114	30	115
rect	29	116	30	117
rect	29	117	30	118
rect	29	119	30	120
rect	29	120	30	121
rect	29	122	30	123
rect	29	123	30	124
rect	29	125	30	126
rect	29	126	30	127
rect	29	128	30	129
rect	29	129	30	130
rect	29	131	30	132
rect	29	132	30	133
rect	29	134	30	135
rect	29	135	30	136
rect	29	137	30	138
rect	29	138	30	139
rect	29	140	30	141
rect	29	141	30	142
rect	29	143	30	144
rect	29	144	30	145
rect	29	146	30	147
rect	29	147	30	148
rect	29	149	30	150
rect	29	150	30	151
rect	29	152	30	153
rect	29	153	30	154
rect	29	155	30	156
rect	29	156	30	157
rect	29	158	30	159
rect	29	159	30	160
rect	29	161	30	162
rect	29	162	30	163
rect	29	164	30	165
rect	29	165	30	166
rect	29	167	30	168
rect	29	168	30	169
rect	31	35	32	36
rect	31	36	32	37
rect	31	38	32	39
rect	31	39	32	40
rect	31	41	32	42
rect	31	42	32	43
rect	31	44	32	45
rect	31	45	32	46
rect	31	47	32	48
rect	31	48	32	49
rect	31	50	32	51
rect	31	51	32	52
rect	31	53	32	54
rect	31	54	32	55
rect	31	56	32	57
rect	31	57	32	58
rect	31	59	32	60
rect	31	60	32	61
rect	31	62	32	63
rect	31	63	32	64
rect	31	65	32	66
rect	31	66	32	67
rect	31	68	32	69
rect	31	69	32	70
rect	31	71	32	72
rect	31	72	32	73
rect	31	74	32	75
rect	31	75	32	76
rect	31	77	32	78
rect	31	78	32	79
rect	31	80	32	81
rect	31	81	32	82
rect	31	83	32	84
rect	31	84	32	85
rect	31	86	32	87
rect	31	87	32	88
rect	31	89	32	90
rect	31	90	32	91
rect	31	92	32	93
rect	31	93	32	94
rect	31	95	32	96
rect	31	96	32	97
rect	31	98	32	99
rect	31	99	32	100
rect	31	101	32	102
rect	31	102	32	103
rect	31	104	32	105
rect	31	105	32	106
rect	31	107	32	108
rect	31	108	32	109
rect	31	110	32	111
rect	31	111	32	112
rect	31	113	32	114
rect	31	114	32	115
rect	31	116	32	117
rect	31	117	32	118
rect	31	119	32	120
rect	31	120	32	121
rect	31	122	32	123
rect	31	123	32	124
rect	31	125	32	126
rect	31	126	32	127
rect	31	128	32	129
rect	31	129	32	130
rect	31	131	32	132
rect	31	132	32	133
rect	31	134	32	135
rect	31	135	32	136
rect	31	137	32	138
rect	31	138	32	139
rect	31	140	32	141
rect	31	141	32	142
rect	31	143	32	144
rect	31	144	32	145
rect	31	146	32	147
rect	31	147	32	148
rect	31	149	32	150
rect	31	150	32	151
rect	31	152	32	153
rect	31	153	32	154
rect	31	155	32	156
rect	31	156	32	157
rect	31	158	32	159
rect	31	159	32	160
rect	31	161	32	162
rect	31	162	32	163
rect	31	164	32	165
rect	31	165	32	166
rect	31	167	32	168
rect	31	168	32	169
rect	31	170	32	171
rect	31	171	32	172
rect	31	173	32	174
rect	31	174	32	175
rect	31	176	32	177
rect	31	177	32	178
rect	31	179	32	180
rect	31	180	32	181
rect	31	182	32	183
rect	31	183	32	184
rect	31	185	32	186
rect	31	186	32	187
rect	31	188	32	189
rect	31	189	32	190
rect	31	191	32	192
rect	31	192	32	193
rect	33	29	34	30
rect	33	30	34	31
rect	33	32	34	33
rect	33	33	34	34
rect	33	35	34	36
rect	33	36	34	37
rect	33	38	34	39
rect	33	39	34	40
rect	33	92	34	93
rect	33	93	34	94
rect	33	95	34	96
rect	33	96	34	97
rect	33	104	34	105
rect	33	105	34	106
rect	33	107	34	108
rect	33	108	34	109
rect	33	110	34	111
rect	33	111	34	112
rect	33	113	34	114
rect	33	114	34	115
rect	33	116	34	117
rect	33	117	34	118
rect	33	119	34	120
rect	33	120	34	121
rect	33	122	34	123
rect	33	123	34	124
rect	33	125	34	126
rect	33	126	34	127
rect	33	128	34	129
rect	33	129	34	130
rect	33	131	34	132
rect	33	132	34	133
rect	33	134	34	135
rect	33	135	34	136
rect	33	137	34	138
rect	33	138	34	139
rect	33	140	34	141
rect	33	141	34	142
rect	33	143	34	144
rect	33	144	34	145
rect	33	146	34	147
rect	33	147	34	148
rect	33	149	34	150
rect	33	150	34	151
rect	33	152	34	153
rect	33	153	34	154
rect	33	155	34	156
rect	33	156	34	157
rect	33	158	34	159
rect	33	159	34	160
rect	33	161	34	162
rect	33	162	34	163
rect	33	164	34	165
rect	33	165	34	166
rect	33	167	34	168
rect	33	168	34	169
rect	33	170	34	171
rect	33	171	34	172
rect	33	173	34	174
rect	33	174	34	175
rect	33	176	34	177
rect	33	177	34	178
rect	33	179	34	180
rect	33	180	34	181
rect	33	182	34	183
rect	33	183	34	184
rect	33	185	34	186
rect	33	186	34	187
rect	33	188	34	189
rect	33	189	34	190
rect	33	191	34	192
rect	33	192	34	193
rect	33	194	34	195
rect	33	195	34	196
rect	33	197	34	198
rect	33	198	34	199
rect	33	200	34	201
rect	33	201	34	202
rect	33	203	34	204
rect	33	204	34	205
rect	35	11	36	12
rect	35	12	36	13
rect	35	14	36	15
rect	35	15	36	16
rect	35	17	36	18
rect	35	18	36	19
rect	35	20	36	21
rect	35	21	36	22
rect	35	23	36	24
rect	35	24	36	25
rect	35	26	36	27
rect	35	27	36	28
rect	35	29	36	30
rect	35	30	36	31
rect	35	32	36	33
rect	35	33	36	34
rect	35	35	36	36
rect	35	36	36	37
rect	35	38	36	39
rect	35	39	36	40
rect	35	41	36	42
rect	35	42	36	43
rect	35	44	36	45
rect	35	45	36	46
rect	35	47	36	48
rect	35	48	36	49
rect	35	50	36	51
rect	35	51	36	52
rect	35	53	36	54
rect	35	54	36	55
rect	35	56	36	57
rect	35	57	36	58
rect	35	59	36	60
rect	35	60	36	61
rect	35	62	36	63
rect	35	63	36	64
rect	35	65	36	66
rect	35	66	36	67
rect	35	68	36	69
rect	35	69	36	70
rect	35	71	36	72
rect	35	72	36	73
rect	35	74	36	75
rect	35	75	36	76
rect	35	77	36	78
rect	35	78	36	79
rect	35	80	36	81
rect	35	81	36	82
rect	35	83	36	84
rect	35	84	36	85
rect	35	86	36	87
rect	35	87	36	88
rect	35	89	36	90
rect	35	90	36	91
rect	35	92	36	93
rect	35	93	36	94
rect	35	95	36	96
rect	35	96	36	97
rect	35	98	36	99
rect	35	99	36	100
rect	35	101	36	102
rect	35	102	36	103
rect	35	104	36	105
rect	35	105	36	106
rect	35	107	36	108
rect	35	108	36	109
rect	35	110	36	111
rect	35	111	36	112
rect	35	113	36	114
rect	35	114	36	115
rect	35	116	36	117
rect	35	117	36	118
rect	35	119	36	120
rect	35	120	36	121
rect	35	122	36	123
rect	35	123	36	124
rect	35	125	36	126
rect	35	126	36	127
rect	35	128	36	129
rect	35	129	36	130
rect	35	131	36	132
rect	35	132	36	133
rect	35	134	36	135
rect	35	135	36	136
rect	35	137	36	138
rect	35	138	36	139
rect	35	140	36	141
rect	35	141	36	142
rect	35	143	36	144
rect	35	144	36	145
rect	44	224	45	225
rect	44	225	45	226
rect	44	227	45	228
rect	44	228	45	229
rect	46	11	47	12
rect	46	12	47	13
rect	46	14	47	15
rect	46	15	47	16
rect	46	17	47	18
rect	46	18	47	19
rect	46	86	47	87
rect	46	87	47	88
rect	46	89	47	90
rect	46	90	47	91
rect	46	101	47	102
rect	46	102	47	103
rect	46	104	47	105
rect	46	105	47	106
rect	46	107	47	108
rect	46	108	47	109
rect	46	110	47	111
rect	46	111	47	112
rect	46	131	47	132
rect	46	132	47	133
rect	46	134	47	135
rect	46	135	47	136
rect	46	179	47	180
rect	46	180	47	181
rect	46	185	47	186
rect	46	186	47	187
rect	46	188	47	189
rect	46	189	47	190
rect	46	209	47	210
rect	46	210	47	211
rect	46	212	47	213
rect	46	213	47	214
rect	46	215	47	216
rect	46	216	47	217
rect	46	218	47	219
rect	46	219	47	220
rect	46	221	47	222
rect	46	222	47	223
rect	46	224	47	225
rect	46	225	47	226
rect	46	239	47	240
rect	46	240	47	241
rect	55	116	56	117
rect	55	117	56	118
rect	55	119	56	120
rect	55	120	56	121
rect	55	122	56	123
rect	55	123	56	124
rect	55	293	56	294
rect	55	294	56	295
rect	55	296	56	297
rect	55	297	56	298
rect	57	71	58	72
rect	57	72	58	73
rect	57	74	58	75
rect	57	75	58	76
rect	57	77	58	78
rect	57	78	58	79
rect	57	80	58	81
rect	57	81	58	82
rect	57	83	58	84
rect	57	84	58	85
rect	57	86	58	87
rect	57	87	58	88
rect	57	89	58	90
rect	57	90	58	91
rect	57	92	58	93
rect	57	93	58	94
rect	57	95	58	96
rect	57	96	58	97
rect	57	98	58	99
rect	57	99	58	100
rect	57	101	58	102
rect	57	102	58	103
rect	57	104	58	105
rect	57	105	58	106
rect	57	107	58	108
rect	57	108	58	109
rect	57	110	58	111
rect	57	111	58	112
rect	57	113	58	114
rect	57	114	58	115
rect	57	116	58	117
rect	57	117	58	118
rect	57	119	58	120
rect	57	120	58	121
rect	57	122	58	123
rect	57	123	58	124
rect	57	125	58	126
rect	57	126	58	127
rect	57	128	58	129
rect	57	129	58	130
rect	57	131	58	132
rect	57	132	58	133
rect	57	134	58	135
rect	57	135	58	136
rect	57	137	58	138
rect	57	138	58	139
rect	57	140	58	141
rect	57	141	58	142
rect	57	143	58	144
rect	57	144	58	145
rect	57	146	58	147
rect	57	147	58	148
rect	57	149	58	150
rect	57	150	58	151
rect	57	152	58	153
rect	57	153	58	154
rect	57	155	58	156
rect	57	156	58	157
rect	57	158	58	159
rect	57	159	58	160
rect	57	161	58	162
rect	57	162	58	163
rect	57	164	58	165
rect	57	165	58	166
rect	57	167	58	168
rect	57	168	58	169
rect	57	170	58	171
rect	57	171	58	172
rect	57	173	58	174
rect	57	174	58	175
rect	57	176	58	177
rect	57	177	58	178
rect	57	179	58	180
rect	57	180	58	181
rect	57	182	58	183
rect	57	183	58	184
rect	57	185	58	186
rect	57	186	58	187
rect	57	188	58	189
rect	57	189	58	190
rect	57	191	58	192
rect	57	192	58	193
rect	57	194	58	195
rect	57	195	58	196
rect	57	197	58	198
rect	57	198	58	199
rect	57	200	58	201
rect	57	201	58	202
rect	57	203	58	204
rect	57	204	58	205
rect	57	206	58	207
rect	57	207	58	208
rect	57	209	58	210
rect	57	210	58	211
rect	57	212	58	213
rect	57	213	58	214
rect	57	215	58	216
rect	57	216	58	217
rect	57	218	58	219
rect	57	219	58	220
rect	57	221	58	222
rect	57	222	58	223
rect	57	224	58	225
rect	57	225	58	226
rect	57	227	58	228
rect	57	228	58	229
rect	57	230	58	231
rect	57	231	58	232
rect	57	233	58	234
rect	57	234	58	235
rect	57	236	58	237
rect	57	237	58	238
rect	57	239	58	240
rect	57	240	58	241
rect	57	242	58	243
rect	57	243	58	244
rect	57	245	58	246
rect	57	246	58	247
rect	57	248	58	249
rect	57	249	58	250
rect	57	251	58	252
rect	57	252	58	253
rect	57	254	58	255
rect	57	255	58	256
rect	57	257	58	258
rect	57	258	58	259
rect	57	260	58	261
rect	57	261	58	262
rect	57	263	58	264
rect	57	264	58	265
rect	57	266	58	267
rect	57	267	58	268
rect	57	269	58	270
rect	57	270	58	271
rect	57	272	58	273
rect	57	273	58	274
rect	57	275	58	276
rect	57	276	58	277
rect	57	278	58	279
rect	57	279	58	280
rect	57	281	58	282
rect	57	282	58	283
rect	57	284	58	285
rect	57	285	58	286
rect	57	287	58	288
rect	57	288	58	289
rect	57	290	58	291
rect	57	291	58	292
rect	59	56	60	57
rect	59	57	60	58
rect	59	68	60	69
rect	59	69	60	70
rect	59	71	60	72
rect	59	72	60	73
rect	59	74	60	75
rect	59	75	60	76
rect	59	77	60	78
rect	59	78	60	79
rect	59	80	60	81
rect	59	81	60	82
rect	59	83	60	84
rect	59	84	60	85
rect	59	86	60	87
rect	59	87	60	88
rect	59	89	60	90
rect	59	90	60	91
rect	59	92	60	93
rect	59	93	60	94
rect	59	95	60	96
rect	59	96	60	97
rect	59	98	60	99
rect	59	99	60	100
rect	59	101	60	102
rect	59	102	60	103
rect	59	104	60	105
rect	59	105	60	106
rect	59	107	60	108
rect	59	108	60	109
rect	59	110	60	111
rect	59	111	60	112
rect	59	113	60	114
rect	59	114	60	115
rect	59	116	60	117
rect	59	117	60	118
rect	59	119	60	120
rect	59	120	60	121
rect	59	122	60	123
rect	59	123	60	124
rect	59	125	60	126
rect	59	126	60	127
rect	59	128	60	129
rect	59	129	60	130
rect	59	131	60	132
rect	59	132	60	133
rect	59	134	60	135
rect	59	135	60	136
rect	59	137	60	138
rect	59	138	60	139
rect	59	140	60	141
rect	59	141	60	142
rect	59	143	60	144
rect	59	144	60	145
rect	59	146	60	147
rect	59	147	60	148
rect	59	149	60	150
rect	59	150	60	151
rect	59	152	60	153
rect	59	153	60	154
rect	59	155	60	156
rect	59	156	60	157
rect	59	158	60	159
rect	59	159	60	160
rect	59	161	60	162
rect	59	162	60	163
rect	59	164	60	165
rect	59	165	60	166
rect	59	167	60	168
rect	59	168	60	169
rect	59	170	60	171
rect	59	171	60	172
rect	59	173	60	174
rect	59	174	60	175
rect	59	176	60	177
rect	59	177	60	178
rect	59	179	60	180
rect	59	180	60	181
rect	61	32	62	33
rect	61	33	62	34
rect	61	59	62	60
rect	61	60	62	61
rect	61	62	62	63
rect	61	63	62	64
rect	61	65	62	66
rect	61	66	62	67
rect	61	68	62	69
rect	61	69	62	70
rect	61	71	62	72
rect	61	72	62	73
rect	61	74	62	75
rect	61	75	62	76
rect	61	77	62	78
rect	61	78	62	79
rect	61	80	62	81
rect	61	81	62	82
rect	61	83	62	84
rect	61	84	62	85
rect	61	86	62	87
rect	61	87	62	88
rect	61	89	62	90
rect	61	90	62	91
rect	61	92	62	93
rect	61	93	62	94
rect	61	95	62	96
rect	61	96	62	97
rect	61	98	62	99
rect	61	99	62	100
rect	61	101	62	102
rect	61	102	62	103
rect	61	104	62	105
rect	61	105	62	106
rect	61	107	62	108
rect	61	108	62	109
rect	61	110	62	111
rect	61	111	62	112
rect	61	113	62	114
rect	61	114	62	115
rect	61	116	62	117
rect	61	117	62	118
rect	61	119	62	120
rect	61	120	62	121
rect	61	122	62	123
rect	61	123	62	124
rect	61	125	62	126
rect	61	126	62	127
rect	61	128	62	129
rect	61	129	62	130
rect	61	131	62	132
rect	61	132	62	133
rect	61	134	62	135
rect	61	135	62	136
rect	61	137	62	138
rect	61	138	62	139
rect	61	140	62	141
rect	61	141	62	142
rect	61	143	62	144
rect	61	144	62	145
rect	61	146	62	147
rect	61	147	62	148
rect	61	149	62	150
rect	61	150	62	151
rect	61	152	62	153
rect	61	153	62	154
rect	61	155	62	156
rect	61	156	62	157
rect	61	158	62	159
rect	61	159	62	160
rect	61	161	62	162
rect	61	162	62	163
rect	61	164	62	165
rect	61	165	62	166
rect	63	23	64	24
rect	63	24	64	25
rect	63	26	64	27
rect	63	27	64	28
rect	63	29	64	30
rect	63	30	64	31
rect	63	32	64	33
rect	63	33	64	34
rect	63	35	64	36
rect	63	36	64	37
rect	63	38	64	39
rect	63	39	64	40
rect	63	41	64	42
rect	63	42	64	43
rect	63	44	64	45
rect	63	45	64	46
rect	63	47	64	48
rect	63	48	64	49
rect	63	50	64	51
rect	63	51	64	52
rect	63	53	64	54
rect	63	54	64	55
rect	63	56	64	57
rect	63	57	64	58
rect	63	59	64	60
rect	63	60	64	61
rect	63	62	64	63
rect	63	63	64	64
rect	63	65	64	66
rect	63	66	64	67
rect	63	68	64	69
rect	63	69	64	70
rect	63	71	64	72
rect	63	72	64	73
rect	63	74	64	75
rect	63	75	64	76
rect	63	77	64	78
rect	63	78	64	79
rect	63	80	64	81
rect	63	81	64	82
rect	63	83	64	84
rect	63	84	64	85
rect	63	86	64	87
rect	63	87	64	88
rect	63	89	64	90
rect	63	90	64	91
rect	63	92	64	93
rect	63	93	64	94
rect	63	95	64	96
rect	63	96	64	97
rect	63	98	64	99
rect	63	99	64	100
rect	63	101	64	102
rect	63	102	64	103
rect	63	104	64	105
rect	63	105	64	106
rect	63	107	64	108
rect	63	108	64	109
rect	63	110	64	111
rect	63	111	64	112
rect	63	113	64	114
rect	63	114	64	115
rect	63	116	64	117
rect	63	117	64	118
rect	63	119	64	120
rect	63	120	64	121
rect	63	122	64	123
rect	63	123	64	124
rect	63	125	64	126
rect	63	126	64	127
rect	63	128	64	129
rect	63	129	64	130
rect	63	131	64	132
rect	63	132	64	133
rect	63	134	64	135
rect	63	135	64	136
rect	63	137	64	138
rect	63	138	64	139
rect	63	140	64	141
rect	63	141	64	142
rect	63	143	64	144
rect	63	144	64	145
rect	63	146	64	147
rect	63	147	64	148
rect	63	149	64	150
rect	63	150	64	151
rect	63	152	64	153
rect	63	153	64	154
rect	63	155	64	156
rect	63	156	64	157
rect	63	158	64	159
rect	63	159	64	160
rect	63	161	64	162
rect	63	162	64	163
rect	63	164	64	165
rect	63	165	64	166
rect	63	167	64	168
rect	63	168	64	169
rect	63	170	64	171
rect	63	171	64	172
rect	63	173	64	174
rect	63	174	64	175
rect	63	176	64	177
rect	63	177	64	178
rect	63	179	64	180
rect	63	180	64	181
rect	63	182	64	183
rect	63	183	64	184
rect	63	185	64	186
rect	63	186	64	187
rect	63	188	64	189
rect	63	189	64	190
rect	63	191	64	192
rect	63	192	64	193
rect	63	194	64	195
rect	63	195	64	196
rect	63	197	64	198
rect	63	198	64	199
rect	63	200	64	201
rect	63	201	64	202
rect	63	203	64	204
rect	63	204	64	205
rect	63	206	64	207
rect	63	207	64	208
rect	63	209	64	210
rect	63	210	64	211
rect	63	212	64	213
rect	63	213	64	214
rect	63	215	64	216
rect	63	216	64	217
rect	63	218	64	219
rect	63	219	64	220
rect	63	221	64	222
rect	63	222	64	223
rect	63	224	64	225
rect	63	225	64	226
rect	63	227	64	228
rect	63	228	64	229
rect	63	230	64	231
rect	63	231	64	232
rect	63	233	64	234
rect	63	234	64	235
rect	63	236	64	237
rect	63	237	64	238
rect	63	239	64	240
rect	63	240	64	241
rect	63	242	64	243
rect	63	243	64	244
rect	63	245	64	246
rect	63	246	64	247
rect	63	248	64	249
rect	63	249	64	250
rect	63	251	64	252
rect	63	252	64	253
rect	63	254	64	255
rect	63	255	64	256
rect	63	257	64	258
rect	63	258	64	259
rect	63	260	64	261
rect	63	261	64	262
rect	63	263	64	264
rect	63	264	64	265
rect	72	95	73	96
rect	72	96	73	97
rect	72	140	73	141
rect	72	141	73	142
rect	72	143	73	144
rect	72	144	73	145
rect	72	146	73	147
rect	72	147	73	148
rect	72	149	73	150
rect	72	150	73	151
rect	72	152	73	153
rect	72	153	73	154
rect	72	155	73	156
rect	72	156	73	157
rect	72	158	73	159
rect	72	159	73	160
rect	72	161	73	162
rect	72	162	73	163
rect	72	164	73	165
rect	72	165	73	166
rect	72	167	73	168
rect	72	168	73	169
rect	72	170	73	171
rect	72	171	73	172
rect	72	173	73	174
rect	72	174	73	175
rect	72	176	73	177
rect	72	177	73	178
rect	72	179	73	180
rect	72	180	73	181
rect	72	182	73	183
rect	72	183	73	184
rect	72	185	73	186
rect	72	186	73	187
rect	72	188	73	189
rect	72	189	73	190
rect	72	191	73	192
rect	72	192	73	193
rect	72	194	73	195
rect	72	195	73	196
rect	72	197	73	198
rect	72	198	73	199
rect	72	200	73	201
rect	72	201	73	202
rect	72	203	73	204
rect	72	204	73	205
rect	72	206	73	207
rect	72	207	73	208
rect	72	209	73	210
rect	72	210	73	211
rect	72	212	73	213
rect	72	213	73	214
rect	72	215	73	216
rect	72	216	73	217
rect	72	218	73	219
rect	72	219	73	220
rect	72	221	73	222
rect	72	222	73	223
rect	72	224	73	225
rect	72	225	73	226
rect	72	227	73	228
rect	72	228	73	229
rect	72	230	73	231
rect	72	231	73	232
rect	72	233	73	234
rect	72	234	73	235
rect	72	236	73	237
rect	72	237	73	238
rect	72	239	73	240
rect	72	240	73	241
rect	72	242	73	243
rect	72	243	73	244
rect	72	245	73	246
rect	72	246	73	247
rect	72	248	73	249
rect	72	249	73	250
rect	72	251	73	252
rect	72	252	73	253
rect	72	254	73	255
rect	72	255	73	256
rect	72	257	73	258
rect	72	258	73	259
rect	72	260	73	261
rect	72	261	73	262
rect	72	263	73	264
rect	72	264	73	265
rect	72	266	73	267
rect	72	267	73	268
rect	72	269	73	270
rect	72	270	73	271
rect	72	272	73	273
rect	72	273	73	274
rect	72	275	73	276
rect	72	276	73	277
rect	72	278	73	279
rect	72	279	73	280
rect	72	281	73	282
rect	72	282	73	283
rect	72	284	73	285
rect	72	285	73	286
rect	72	287	73	288
rect	72	288	73	289
rect	72	290	73	291
rect	72	291	73	292
rect	72	293	73	294
rect	72	294	73	295
rect	72	296	73	297
rect	72	297	73	298
rect	72	299	73	300
rect	72	300	73	301
rect	72	302	73	303
rect	72	303	73	304
rect	72	305	73	306
rect	72	306	73	307
rect	74	65	75	66
rect	74	66	75	67
rect	74	68	75	69
rect	74	69	75	70
rect	74	71	75	72
rect	74	72	75	73
rect	74	74	75	75
rect	74	75	75	76
rect	74	77	75	78
rect	74	78	75	79
rect	74	80	75	81
rect	74	81	75	82
rect	74	83	75	84
rect	74	84	75	85
rect	74	86	75	87
rect	74	87	75	88
rect	74	89	75	90
rect	74	90	75	91
rect	74	92	75	93
rect	74	93	75	94
rect	74	95	75	96
rect	74	96	75	97
rect	74	98	75	99
rect	74	99	75	100
rect	74	101	75	102
rect	74	102	75	103
rect	74	104	75	105
rect	74	105	75	106
rect	74	107	75	108
rect	74	108	75	109
rect	74	110	75	111
rect	74	111	75	112
rect	74	113	75	114
rect	74	114	75	115
rect	74	116	75	117
rect	74	117	75	118
rect	74	119	75	120
rect	74	120	75	121
rect	74	122	75	123
rect	74	123	75	124
rect	74	125	75	126
rect	74	126	75	127
rect	74	128	75	129
rect	74	129	75	130
rect	74	131	75	132
rect	74	132	75	133
rect	74	134	75	135
rect	74	135	75	136
rect	74	137	75	138
rect	74	138	75	139
rect	74	140	75	141
rect	74	141	75	142
rect	74	143	75	144
rect	74	144	75	145
rect	74	146	75	147
rect	74	147	75	148
rect	74	149	75	150
rect	74	150	75	151
rect	74	152	75	153
rect	74	153	75	154
rect	74	155	75	156
rect	74	156	75	157
rect	74	158	75	159
rect	74	159	75	160
rect	74	161	75	162
rect	74	162	75	163
rect	74	164	75	165
rect	74	165	75	166
rect	74	167	75	168
rect	74	168	75	169
rect	74	170	75	171
rect	74	171	75	172
rect	74	173	75	174
rect	74	174	75	175
rect	74	176	75	177
rect	74	177	75	178
rect	74	179	75	180
rect	74	180	75	181
rect	74	182	75	183
rect	74	183	75	184
rect	74	185	75	186
rect	74	186	75	187
rect	74	188	75	189
rect	74	189	75	190
rect	74	191	75	192
rect	74	192	75	193
rect	74	194	75	195
rect	74	195	75	196
rect	74	197	75	198
rect	74	198	75	199
rect	74	200	75	201
rect	74	201	75	202
rect	74	203	75	204
rect	74	204	75	205
rect	74	206	75	207
rect	74	207	75	208
rect	74	209	75	210
rect	74	210	75	211
rect	74	212	75	213
rect	74	213	75	214
rect	74	215	75	216
rect	74	216	75	217
rect	74	218	75	219
rect	74	219	75	220
rect	74	221	75	222
rect	74	222	75	223
rect	74	224	75	225
rect	74	225	75	226
rect	74	227	75	228
rect	74	228	75	229
rect	74	230	75	231
rect	74	231	75	232
rect	74	233	75	234
rect	74	234	75	235
rect	74	236	75	237
rect	74	237	75	238
rect	74	239	75	240
rect	74	240	75	241
rect	74	242	75	243
rect	74	243	75	244
rect	74	245	75	246
rect	74	246	75	247
rect	74	248	75	249
rect	74	249	75	250
rect	74	251	75	252
rect	74	252	75	253
rect	74	254	75	255
rect	74	255	75	256
rect	74	257	75	258
rect	74	258	75	259
rect	74	260	75	261
rect	74	261	75	262
rect	74	263	75	264
rect	74	264	75	265
rect	74	266	75	267
rect	74	267	75	268
rect	74	269	75	270
rect	74	270	75	271
rect	74	272	75	273
rect	74	273	75	274
rect	74	275	75	276
rect	74	276	75	277
rect	74	278	75	279
rect	74	279	75	280
rect	74	281	75	282
rect	74	282	75	283
rect	74	284	75	285
rect	74	285	75	286
rect	76	62	77	63
rect	76	63	77	64
rect	76	65	77	66
rect	76	66	77	67
rect	76	68	77	69
rect	76	69	77	70
rect	76	71	77	72
rect	76	72	77	73
rect	76	74	77	75
rect	76	75	77	76
rect	76	77	77	78
rect	76	78	77	79
rect	76	80	77	81
rect	76	81	77	82
rect	76	83	77	84
rect	76	84	77	85
rect	76	86	77	87
rect	76	87	77	88
rect	76	89	77	90
rect	76	90	77	91
rect	76	92	77	93
rect	76	93	77	94
rect	76	95	77	96
rect	76	96	77	97
rect	76	98	77	99
rect	76	99	77	100
rect	76	101	77	102
rect	76	102	77	103
rect	76	104	77	105
rect	76	105	77	106
rect	76	107	77	108
rect	76	108	77	109
rect	76	110	77	111
rect	76	111	77	112
rect	76	113	77	114
rect	76	114	77	115
rect	76	116	77	117
rect	76	117	77	118
rect	76	119	77	120
rect	76	120	77	121
rect	76	122	77	123
rect	76	123	77	124
rect	76	125	77	126
rect	76	126	77	127
rect	76	128	77	129
rect	76	129	77	130
rect	76	131	77	132
rect	76	132	77	133
rect	76	134	77	135
rect	76	135	77	136
rect	76	137	77	138
rect	76	138	77	139
rect	76	140	77	141
rect	76	141	77	142
rect	76	143	77	144
rect	76	144	77	145
rect	76	146	77	147
rect	76	147	77	148
rect	76	149	77	150
rect	76	150	77	151
rect	76	152	77	153
rect	76	153	77	154
rect	76	155	77	156
rect	76	156	77	157
rect	76	158	77	159
rect	76	159	77	160
rect	76	161	77	162
rect	76	162	77	163
rect	76	164	77	165
rect	76	165	77	166
rect	76	167	77	168
rect	76	168	77	169
rect	76	170	77	171
rect	76	171	77	172
rect	76	173	77	174
rect	76	174	77	175
rect	76	176	77	177
rect	76	177	77	178
rect	76	179	77	180
rect	76	180	77	181
rect	76	182	77	183
rect	76	183	77	184
rect	76	185	77	186
rect	76	186	77	187
rect	76	188	77	189
rect	76	189	77	190
rect	76	191	77	192
rect	76	192	77	193
rect	76	194	77	195
rect	76	195	77	196
rect	76	197	77	198
rect	76	198	77	199
rect	76	200	77	201
rect	76	201	77	202
rect	76	203	77	204
rect	76	204	77	205
rect	76	206	77	207
rect	76	207	77	208
rect	76	209	77	210
rect	76	210	77	211
rect	76	212	77	213
rect	76	213	77	214
rect	76	215	77	216
rect	76	216	77	217
rect	76	218	77	219
rect	76	219	77	220
rect	76	221	77	222
rect	76	222	77	223
rect	76	224	77	225
rect	76	225	77	226
rect	76	227	77	228
rect	76	228	77	229
rect	76	230	77	231
rect	76	231	77	232
rect	76	233	77	234
rect	76	234	77	235
rect	76	236	77	237
rect	76	237	77	238
rect	76	239	77	240
rect	76	240	77	241
rect	76	242	77	243
rect	76	243	77	244
rect	76	245	77	246
rect	76	246	77	247
rect	76	248	77	249
rect	76	249	77	250
rect	76	251	77	252
rect	76	252	77	253
rect	76	254	77	255
rect	76	255	77	256
rect	76	257	77	258
rect	76	258	77	259
rect	76	260	77	261
rect	76	261	77	262
rect	76	263	77	264
rect	76	264	77	265
rect	76	266	77	267
rect	76	267	77	268
rect	76	269	77	270
rect	76	270	77	271
rect	76	293	77	294
rect	76	294	77	295
rect	76	296	77	297
rect	76	297	77	298
rect	76	299	77	300
rect	76	300	77	301
rect	76	302	77	303
rect	76	303	77	304
rect	76	305	77	306
rect	76	306	77	307
rect	76	308	77	309
rect	76	309	77	310
rect	78	11	79	12
rect	78	12	79	13
rect	78	32	79	33
rect	78	33	79	34
rect	78	35	79	36
rect	78	36	79	37
rect	78	38	79	39
rect	78	39	79	40
rect	78	41	79	42
rect	78	42	79	43
rect	78	44	79	45
rect	78	45	79	46
rect	78	47	79	48
rect	78	48	79	49
rect	78	50	79	51
rect	78	51	79	52
rect	78	53	79	54
rect	78	54	79	55
rect	78	56	79	57
rect	78	57	79	58
rect	78	59	79	60
rect	78	60	79	61
rect	78	62	79	63
rect	78	63	79	64
rect	78	65	79	66
rect	78	66	79	67
rect	78	68	79	69
rect	78	69	79	70
rect	78	71	79	72
rect	78	72	79	73
rect	78	74	79	75
rect	78	75	79	76
rect	78	77	79	78
rect	78	78	79	79
rect	78	80	79	81
rect	78	81	79	82
rect	78	83	79	84
rect	78	84	79	85
rect	78	86	79	87
rect	78	87	79	88
rect	78	89	79	90
rect	78	90	79	91
rect	78	92	79	93
rect	78	93	79	94
rect	78	95	79	96
rect	78	96	79	97
rect	78	98	79	99
rect	78	99	79	100
rect	78	101	79	102
rect	78	102	79	103
rect	78	104	79	105
rect	78	105	79	106
rect	78	107	79	108
rect	78	108	79	109
rect	78	110	79	111
rect	78	111	79	112
rect	78	113	79	114
rect	78	114	79	115
rect	78	116	79	117
rect	78	117	79	118
rect	78	119	79	120
rect	78	120	79	121
rect	78	122	79	123
rect	78	123	79	124
rect	78	125	79	126
rect	78	126	79	127
rect	78	128	79	129
rect	78	129	79	130
rect	78	131	79	132
rect	78	132	79	133
rect	78	134	79	135
rect	78	135	79	136
rect	78	137	79	138
rect	78	138	79	139
rect	78	140	79	141
rect	78	141	79	142
rect	78	143	79	144
rect	78	144	79	145
rect	78	146	79	147
rect	78	147	79	148
rect	78	149	79	150
rect	78	150	79	151
rect	78	152	79	153
rect	78	153	79	154
rect	78	155	79	156
rect	78	156	79	157
rect	78	158	79	159
rect	78	159	79	160
rect	78	161	79	162
rect	78	162	79	163
rect	78	164	79	165
rect	78	165	79	166
rect	78	167	79	168
rect	78	168	79	169
rect	78	170	79	171
rect	78	171	79	172
rect	78	173	79	174
rect	78	174	79	175
rect	78	176	79	177
rect	78	177	79	178
rect	78	179	79	180
rect	78	180	79	181
rect	78	182	79	183
rect	78	183	79	184
rect	78	185	79	186
rect	78	186	79	187
rect	78	188	79	189
rect	78	189	79	190
rect	78	191	79	192
rect	78	192	79	193
rect	78	194	79	195
rect	78	195	79	196
rect	78	197	79	198
rect	78	198	79	199
rect	78	215	79	216
rect	78	216	79	217
rect	78	272	79	273
rect	78	273	79	274
rect	78	275	79	276
rect	78	276	79	277
rect	78	278	79	279
rect	78	279	79	280
rect	78	281	79	282
rect	78	282	79	283
rect	78	287	79	288
rect	78	288	79	289
rect	78	290	79	291
rect	78	291	79	292
rect	78	299	79	300
rect	78	300	79	301
rect	87	86	88	87
rect	87	87	88	88
rect	87	89	88	90
rect	87	90	88	91
rect	87	92	88	93
rect	87	93	88	94
rect	87	95	88	96
rect	87	96	88	97
rect	87	98	88	99
rect	87	99	88	100
rect	87	113	88	114
rect	87	114	88	115
rect	89	35	90	36
rect	89	36	90	37
rect	89	38	90	39
rect	89	39	90	40
rect	89	41	90	42
rect	89	42	90	43
rect	89	44	90	45
rect	89	45	90	46
rect	89	47	90	48
rect	89	48	90	49
rect	89	50	90	51
rect	89	51	90	52
rect	89	53	90	54
rect	89	54	90	55
rect	89	56	90	57
rect	89	57	90	58
rect	89	59	90	60
rect	89	60	90	61
rect	89	62	90	63
rect	89	63	90	64
rect	89	65	90	66
rect	89	66	90	67
rect	89	68	90	69
rect	89	69	90	70
rect	89	71	90	72
rect	89	72	90	73
rect	89	74	90	75
rect	89	75	90	76
rect	89	77	90	78
rect	89	78	90	79
rect	89	80	90	81
rect	89	81	90	82
rect	89	83	90	84
rect	89	84	90	85
rect	89	86	90	87
rect	89	87	90	88
rect	89	89	90	90
rect	89	90	90	91
rect	89	92	90	93
rect	89	93	90	94
rect	89	95	90	96
rect	89	96	90	97
rect	89	98	90	99
rect	89	99	90	100
rect	89	101	90	102
rect	89	102	90	103
rect	89	104	90	105
rect	89	105	90	106
rect	89	107	90	108
rect	89	108	90	109
rect	89	110	90	111
rect	89	111	90	112
rect	89	113	90	114
rect	89	114	90	115
rect	89	116	90	117
rect	89	117	90	118
rect	89	119	90	120
rect	89	120	90	121
rect	89	122	90	123
rect	89	123	90	124
rect	89	125	90	126
rect	89	126	90	127
rect	89	128	90	129
rect	89	129	90	130
rect	89	131	90	132
rect	89	132	90	133
rect	89	134	90	135
rect	89	135	90	136
rect	89	137	90	138
rect	89	138	90	139
rect	89	140	90	141
rect	89	141	90	142
rect	89	143	90	144
rect	89	144	90	145
rect	89	146	90	147
rect	89	147	90	148
rect	89	149	90	150
rect	89	150	90	151
rect	89	152	90	153
rect	89	153	90	154
rect	89	155	90	156
rect	89	156	90	157
rect	89	158	90	159
rect	89	159	90	160
rect	89	161	90	162
rect	89	162	90	163
rect	89	224	90	225
rect	89	225	90	226
rect	89	227	90	228
rect	89	228	90	229
rect	91	17	92	18
rect	91	18	92	19
rect	91	20	92	21
rect	91	21	92	22
rect	91	23	92	24
rect	91	24	92	25
rect	91	26	92	27
rect	91	27	92	28
rect	91	29	92	30
rect	91	30	92	31
rect	91	32	92	33
rect	91	33	92	34
rect	91	35	92	36
rect	91	36	92	37
rect	91	38	92	39
rect	91	39	92	40
rect	91	41	92	42
rect	91	42	92	43
rect	91	44	92	45
rect	91	45	92	46
rect	91	47	92	48
rect	91	48	92	49
rect	91	50	92	51
rect	91	51	92	52
rect	91	53	92	54
rect	91	54	92	55
rect	91	56	92	57
rect	91	57	92	58
rect	91	59	92	60
rect	91	60	92	61
rect	91	62	92	63
rect	91	63	92	64
rect	91	65	92	66
rect	91	66	92	67
rect	91	68	92	69
rect	91	69	92	70
rect	91	71	92	72
rect	91	72	92	73
rect	91	74	92	75
rect	91	75	92	76
rect	91	77	92	78
rect	91	78	92	79
rect	91	80	92	81
rect	91	81	92	82
rect	91	83	92	84
rect	91	84	92	85
rect	91	86	92	87
rect	91	87	92	88
rect	91	89	92	90
rect	91	90	92	91
rect	91	92	92	93
rect	91	93	92	94
rect	91	95	92	96
rect	91	96	92	97
rect	91	98	92	99
rect	91	99	92	100
rect	91	101	92	102
rect	91	102	92	103
rect	91	104	92	105
rect	91	105	92	106
rect	91	107	92	108
rect	91	108	92	109
rect	91	110	92	111
rect	91	111	92	112
rect	91	113	92	114
rect	91	114	92	115
rect	91	116	92	117
rect	91	117	92	118
rect	91	119	92	120
rect	91	120	92	121
rect	91	122	92	123
rect	91	123	92	124
rect	91	125	92	126
rect	91	126	92	127
rect	91	128	92	129
rect	91	129	92	130
rect	91	131	92	132
rect	91	132	92	133
rect	91	134	92	135
rect	91	135	92	136
rect	91	137	92	138
rect	91	138	92	139
rect	91	140	92	141
rect	91	141	92	142
rect	91	143	92	144
rect	91	144	92	145
rect	91	146	92	147
rect	91	147	92	148
rect	91	149	92	150
rect	91	150	92	151
rect	91	152	92	153
rect	91	153	92	154
rect	91	155	92	156
rect	91	156	92	157
rect	91	158	92	159
rect	91	159	92	160
rect	91	161	92	162
rect	91	162	92	163
rect	91	164	92	165
rect	91	165	92	166
rect	91	167	92	168
rect	91	168	92	169
rect	91	170	92	171
rect	91	171	92	172
rect	91	173	92	174
rect	91	174	92	175
rect	91	176	92	177
rect	91	177	92	178
rect	91	179	92	180
rect	91	180	92	181
rect	91	182	92	183
rect	91	183	92	184
rect	91	185	92	186
rect	91	186	92	187
rect	91	188	92	189
rect	91	189	92	190
rect	91	191	92	192
rect	91	192	92	193
rect	91	194	92	195
rect	91	195	92	196
rect	91	197	92	198
rect	91	198	92	199
rect	91	200	92	201
rect	91	201	92	202
rect	91	203	92	204
rect	91	204	92	205
rect	91	206	92	207
rect	91	207	92	208
rect	91	209	92	210
rect	91	210	92	211
rect	91	212	92	213
rect	91	213	92	214
rect	91	215	92	216
rect	91	216	92	217
rect	91	218	92	219
rect	91	219	92	220
rect	91	221	92	222
rect	91	222	92	223
rect	91	224	92	225
rect	91	225	92	226
rect	91	227	92	228
rect	91	228	92	229
rect	91	230	92	231
rect	91	231	92	232
rect	91	233	92	234
rect	91	234	92	235
rect	91	236	92	237
rect	91	237	92	238
rect	91	239	92	240
rect	91	240	92	241
rect	91	242	92	243
rect	91	243	92	244
rect	91	245	92	246
rect	91	246	92	247
rect	91	248	92	249
rect	91	249	92	250
rect	91	251	92	252
rect	91	252	92	253
rect	91	254	92	255
rect	91	255	92	256
rect	91	257	92	258
rect	91	258	92	259
rect	91	260	92	261
rect	91	261	92	262
rect	91	263	92	264
rect	91	264	92	265
rect	91	266	92	267
rect	91	267	92	268
rect	91	296	92	297
rect	91	297	92	298
rect	91	299	92	300
rect	91	300	92	301
rect	91	308	92	309
rect	91	309	92	310
rect	91	311	92	312
rect	91	312	92	313
rect	100	134	101	135
rect	100	135	101	136
rect	102	62	103	63
rect	102	63	103	64
rect	102	65	103	66
rect	102	66	103	67
rect	102	68	103	69
rect	102	69	103	70
rect	102	71	103	72
rect	102	72	103	73
rect	102	74	103	75
rect	102	75	103	76
rect	102	77	103	78
rect	102	78	103	79
rect	102	80	103	81
rect	102	81	103	82
rect	102	83	103	84
rect	102	84	103	85
rect	102	86	103	87
rect	102	87	103	88
rect	102	89	103	90
rect	102	90	103	91
rect	102	92	103	93
rect	102	93	103	94
rect	102	95	103	96
rect	102	96	103	97
rect	102	98	103	99
rect	102	99	103	100
rect	102	101	103	102
rect	102	102	103	103
rect	102	104	103	105
rect	102	105	103	106
rect	102	107	103	108
rect	102	108	103	109
rect	102	110	103	111
rect	102	111	103	112
rect	102	113	103	114
rect	102	114	103	115
rect	102	116	103	117
rect	102	117	103	118
rect	102	119	103	120
rect	102	120	103	121
rect	102	122	103	123
rect	102	123	103	124
rect	102	125	103	126
rect	102	126	103	127
rect	102	128	103	129
rect	102	129	103	130
rect	102	131	103	132
rect	102	132	103	133
rect	102	134	103	135
rect	102	135	103	136
rect	102	137	103	138
rect	102	138	103	139
rect	102	140	103	141
rect	102	141	103	142
rect	102	143	103	144
rect	102	144	103	145
rect	102	146	103	147
rect	102	147	103	148
rect	102	149	103	150
rect	102	150	103	151
rect	102	152	103	153
rect	102	153	103	154
rect	102	155	103	156
rect	102	156	103	157
rect	102	158	103	159
rect	102	159	103	160
rect	102	161	103	162
rect	102	162	103	163
rect	102	164	103	165
rect	102	165	103	166
rect	102	167	103	168
rect	102	168	103	169
rect	102	170	103	171
rect	102	171	103	172
rect	102	173	103	174
rect	102	174	103	175
rect	102	176	103	177
rect	102	177	103	178
rect	102	179	103	180
rect	102	180	103	181
rect	102	182	103	183
rect	102	183	103	184
rect	102	185	103	186
rect	102	186	103	187
rect	102	188	103	189
rect	102	189	103	190
rect	102	191	103	192
rect	102	192	103	193
rect	102	194	103	195
rect	102	195	103	196
rect	102	197	103	198
rect	102	198	103	199
rect	102	200	103	201
rect	102	201	103	202
rect	102	203	103	204
rect	102	204	103	205
rect	102	206	103	207
rect	102	207	103	208
rect	102	209	103	210
rect	102	210	103	211
rect	102	212	103	213
rect	102	213	103	214
rect	102	215	103	216
rect	102	216	103	217
rect	102	218	103	219
rect	102	219	103	220
rect	102	221	103	222
rect	102	222	103	223
rect	102	224	103	225
rect	102	225	103	226
rect	102	227	103	228
rect	102	228	103	229
rect	102	230	103	231
rect	102	231	103	232
rect	102	233	103	234
rect	102	234	103	235
rect	102	236	103	237
rect	102	237	103	238
rect	102	239	103	240
rect	102	240	103	241
rect	102	242	103	243
rect	102	243	103	244
rect	102	245	103	246
rect	102	246	103	247
rect	102	248	103	249
rect	102	249	103	250
rect	102	251	103	252
rect	102	252	103	253
rect	102	254	103	255
rect	102	255	103	256
rect	104	17	105	18
rect	104	18	105	19
rect	104	23	105	24
rect	104	24	105	25
rect	104	26	105	27
rect	104	27	105	28
rect	104	29	105	30
rect	104	30	105	31
rect	104	32	105	33
rect	104	33	105	34
rect	104	35	105	36
rect	104	36	105	37
rect	104	38	105	39
rect	104	39	105	40
rect	104	41	105	42
rect	104	42	105	43
rect	104	44	105	45
rect	104	45	105	46
rect	104	47	105	48
rect	104	48	105	49
rect	104	50	105	51
rect	104	51	105	52
rect	104	53	105	54
rect	104	54	105	55
rect	104	56	105	57
rect	104	57	105	58
rect	104	59	105	60
rect	104	60	105	61
rect	104	62	105	63
rect	104	63	105	64
rect	104	65	105	66
rect	104	66	105	67
rect	104	68	105	69
rect	104	69	105	70
rect	104	71	105	72
rect	104	72	105	73
rect	104	74	105	75
rect	104	75	105	76
rect	104	77	105	78
rect	104	78	105	79
rect	104	80	105	81
rect	104	81	105	82
rect	104	83	105	84
rect	104	84	105	85
rect	104	86	105	87
rect	104	87	105	88
rect	104	89	105	90
rect	104	90	105	91
rect	104	92	105	93
rect	104	93	105	94
rect	104	95	105	96
rect	104	96	105	97
rect	104	98	105	99
rect	104	99	105	100
rect	104	101	105	102
rect	104	102	105	103
rect	104	104	105	105
rect	104	105	105	106
rect	104	107	105	108
rect	104	108	105	109
rect	104	110	105	111
rect	104	111	105	112
rect	104	113	105	114
rect	104	114	105	115
rect	104	116	105	117
rect	104	117	105	118
rect	104	119	105	120
rect	104	120	105	121
rect	104	122	105	123
rect	104	123	105	124
rect	104	125	105	126
rect	104	126	105	127
rect	104	128	105	129
rect	104	129	105	130
rect	104	131	105	132
rect	104	132	105	133
rect	104	134	105	135
rect	104	135	105	136
rect	104	137	105	138
rect	104	138	105	139
rect	104	140	105	141
rect	104	141	105	142
rect	104	143	105	144
rect	104	144	105	145
rect	104	146	105	147
rect	104	147	105	148
rect	104	149	105	150
rect	104	150	105	151
rect	104	152	105	153
rect	104	153	105	154
rect	104	155	105	156
rect	104	156	105	157
rect	104	158	105	159
rect	104	159	105	160
rect	104	161	105	162
rect	104	162	105	163
rect	104	164	105	165
rect	104	165	105	166
rect	104	167	105	168
rect	104	168	105	169
rect	104	170	105	171
rect	104	171	105	172
rect	104	173	105	174
rect	104	174	105	175
rect	104	176	105	177
rect	104	177	105	178
rect	104	179	105	180
rect	104	180	105	181
rect	104	182	105	183
rect	104	183	105	184
rect	104	185	105	186
rect	104	186	105	187
rect	104	188	105	189
rect	104	189	105	190
rect	104	191	105	192
rect	104	192	105	193
rect	104	194	105	195
rect	104	195	105	196
rect	104	197	105	198
rect	104	198	105	199
rect	104	200	105	201
rect	104	201	105	202
rect	104	203	105	204
rect	104	204	105	205
rect	104	206	105	207
rect	104	207	105	208
rect	104	209	105	210
rect	104	210	105	211
rect	104	212	105	213
rect	104	213	105	214
rect	104	215	105	216
rect	104	216	105	217
rect	104	218	105	219
rect	104	219	105	220
rect	104	221	105	222
rect	104	222	105	223
rect	104	224	105	225
rect	104	225	105	226
rect	104	227	105	228
rect	104	228	105	229
rect	104	230	105	231
rect	104	231	105	232
rect	104	233	105	234
rect	104	234	105	235
rect	104	236	105	237
rect	104	237	105	238
rect	104	239	105	240
rect	104	240	105	241
rect	104	242	105	243
rect	104	243	105	244
rect	104	245	105	246
rect	104	246	105	247
rect	104	248	105	249
rect	104	249	105	250
rect	104	251	105	252
rect	104	252	105	253
rect	104	254	105	255
rect	104	255	105	256
rect	104	257	105	258
rect	104	258	105	259
rect	104	260	105	261
rect	104	261	105	262
rect	104	263	105	264
rect	104	264	105	265
rect	106	11	107	12
rect	106	12	107	13
rect	106	14	107	15
rect	106	15	107	16
rect	106	17	107	18
rect	106	18	107	19
rect	106	20	107	21
rect	106	21	107	22
rect	106	23	107	24
rect	106	24	107	25
rect	106	26	107	27
rect	106	27	107	28
rect	106	29	107	30
rect	106	30	107	31
rect	106	32	107	33
rect	106	33	107	34
rect	106	35	107	36
rect	106	36	107	37
rect	106	38	107	39
rect	106	39	107	40
rect	106	41	107	42
rect	106	42	107	43
rect	106	44	107	45
rect	106	45	107	46
rect	106	47	107	48
rect	106	48	107	49
rect	106	50	107	51
rect	106	51	107	52
rect	106	53	107	54
rect	106	54	107	55
rect	106	56	107	57
rect	106	57	107	58
rect	106	59	107	60
rect	106	60	107	61
rect	106	62	107	63
rect	106	63	107	64
rect	106	65	107	66
rect	106	66	107	67
rect	106	68	107	69
rect	106	69	107	70
rect	106	71	107	72
rect	106	72	107	73
rect	106	74	107	75
rect	106	75	107	76
rect	106	77	107	78
rect	106	78	107	79
rect	106	80	107	81
rect	106	81	107	82
rect	106	83	107	84
rect	106	84	107	85
rect	106	86	107	87
rect	106	87	107	88
rect	106	89	107	90
rect	106	90	107	91
rect	106	92	107	93
rect	106	93	107	94
rect	106	95	107	96
rect	106	96	107	97
rect	106	98	107	99
rect	106	99	107	100
rect	106	101	107	102
rect	106	102	107	103
rect	106	104	107	105
rect	106	105	107	106
rect	106	107	107	108
rect	106	108	107	109
rect	106	110	107	111
rect	106	111	107	112
rect	106	113	107	114
rect	106	114	107	115
rect	106	116	107	117
rect	106	117	107	118
rect	106	119	107	120
rect	106	120	107	121
rect	106	122	107	123
rect	106	123	107	124
rect	106	125	107	126
rect	106	126	107	127
rect	106	128	107	129
rect	106	129	107	130
rect	106	131	107	132
rect	106	132	107	133
rect	106	134	107	135
rect	106	135	107	136
rect	106	137	107	138
rect	106	138	107	139
rect	106	140	107	141
rect	106	141	107	142
rect	106	143	107	144
rect	106	144	107	145
rect	106	146	107	147
rect	106	147	107	148
rect	106	149	107	150
rect	106	150	107	151
rect	106	152	107	153
rect	106	153	107	154
rect	106	155	107	156
rect	106	156	107	157
rect	106	158	107	159
rect	106	159	107	160
rect	106	161	107	162
rect	106	162	107	163
rect	106	164	107	165
rect	106	165	107	166
rect	106	167	107	168
rect	106	168	107	169
rect	106	170	107	171
rect	106	171	107	172
rect	106	173	107	174
rect	106	174	107	175
rect	106	176	107	177
rect	106	177	107	178
rect	106	179	107	180
rect	106	180	107	181
rect	106	182	107	183
rect	106	183	107	184
rect	106	185	107	186
rect	106	186	107	187
rect	106	188	107	189
rect	106	189	107	190
rect	106	191	107	192
rect	106	192	107	193
rect	106	194	107	195
rect	106	195	107	196
rect	106	197	107	198
rect	106	198	107	199
rect	106	200	107	201
rect	106	201	107	202
rect	106	203	107	204
rect	106	204	107	205
rect	106	206	107	207
rect	106	207	107	208
rect	106	209	107	210
rect	106	210	107	211
rect	106	212	107	213
rect	106	213	107	214
rect	106	215	107	216
rect	106	216	107	217
rect	106	218	107	219
rect	106	219	107	220
rect	106	221	107	222
rect	106	222	107	223
rect	106	224	107	225
rect	106	225	107	226
rect	106	227	107	228
rect	106	228	107	229
rect	106	230	107	231
rect	106	231	107	232
rect	106	233	107	234
rect	106	234	107	235
rect	106	236	107	237
rect	106	237	107	238
rect	106	254	107	255
rect	106	255	107	256
rect	106	257	107	258
rect	106	258	107	259
rect	106	287	107	288
rect	106	288	107	289
rect	106	290	107	291
rect	106	291	107	292
rect	115	11	116	12
rect	115	12	116	13
rect	115	14	116	15
rect	115	15	116	16
rect	115	29	116	30
rect	115	30	116	31
rect	115	32	116	33
rect	115	33	116	34
rect	115	35	116	36
rect	115	36	116	37
rect	115	38	116	39
rect	115	39	116	40
rect	115	41	116	42
rect	115	42	116	43
rect	115	44	116	45
rect	115	45	116	46
rect	115	47	116	48
rect	115	48	116	49
rect	115	50	116	51
rect	115	51	116	52
rect	115	53	116	54
rect	115	54	116	55
rect	115	56	116	57
rect	115	57	116	58
rect	115	59	116	60
rect	115	60	116	61
rect	115	62	116	63
rect	115	63	116	64
rect	115	65	116	66
rect	115	66	116	67
rect	115	68	116	69
rect	115	69	116	70
rect	115	71	116	72
rect	115	72	116	73
rect	115	74	116	75
rect	115	75	116	76
rect	115	77	116	78
rect	115	78	116	79
rect	115	80	116	81
rect	115	81	116	82
rect	115	83	116	84
rect	115	84	116	85
rect	115	86	116	87
rect	115	87	116	88
rect	115	89	116	90
rect	115	90	116	91
rect	115	92	116	93
rect	115	93	116	94
rect	115	95	116	96
rect	115	96	116	97
rect	115	98	116	99
rect	115	99	116	100
rect	115	101	116	102
rect	115	102	116	103
rect	115	104	116	105
rect	115	105	116	106
rect	115	107	116	108
rect	115	108	116	109
rect	115	110	116	111
rect	115	111	116	112
rect	115	113	116	114
rect	115	114	116	115
rect	115	116	116	117
rect	115	117	116	118
rect	115	119	116	120
rect	115	120	116	121
rect	115	122	116	123
rect	115	123	116	124
rect	115	125	116	126
rect	115	126	116	127
rect	115	128	116	129
rect	115	129	116	130
rect	115	131	116	132
rect	115	132	116	133
rect	115	134	116	135
rect	115	135	116	136
rect	115	137	116	138
rect	115	138	116	139
rect	115	140	116	141
rect	115	141	116	142
rect	115	143	116	144
rect	115	144	116	145
rect	115	146	116	147
rect	115	147	116	148
rect	115	149	116	150
rect	115	150	116	151
rect	115	152	116	153
rect	115	153	116	154
rect	115	155	116	156
rect	115	156	116	157
rect	115	158	116	159
rect	115	159	116	160
rect	115	161	116	162
rect	115	162	116	163
rect	115	164	116	165
rect	115	165	116	166
rect	115	167	116	168
rect	115	168	116	169
rect	115	170	116	171
rect	115	171	116	172
rect	115	173	116	174
rect	115	174	116	175
rect	115	176	116	177
rect	115	177	116	178
rect	115	179	116	180
rect	115	180	116	181
rect	115	182	116	183
rect	115	183	116	184
rect	115	185	116	186
rect	115	186	116	187
rect	115	188	116	189
rect	115	189	116	190
rect	115	191	116	192
rect	115	192	116	193
rect	115	194	116	195
rect	115	195	116	196
rect	115	197	116	198
rect	115	198	116	199
rect	115	200	116	201
rect	115	201	116	202
rect	115	203	116	204
rect	115	204	116	205
rect	115	206	116	207
rect	115	207	116	208
rect	115	209	116	210
rect	115	210	116	211
rect	117	5	118	6
rect	117	6	118	7
rect	117	11	118	12
rect	117	12	118	13
rect	117	14	118	15
rect	117	15	118	16
rect	117	17	118	18
rect	117	18	118	19
rect	117	20	118	21
rect	117	21	118	22
rect	117	23	118	24
rect	117	24	118	25
rect	117	26	118	27
rect	117	27	118	28
rect	117	29	118	30
rect	117	30	118	31
rect	117	32	118	33
rect	117	33	118	34
rect	117	35	118	36
rect	117	36	118	37
rect	117	38	118	39
rect	117	39	118	40
rect	117	41	118	42
rect	117	42	118	43
rect	117	44	118	45
rect	117	45	118	46
rect	117	47	118	48
rect	117	48	118	49
rect	117	50	118	51
rect	117	51	118	52
rect	117	53	118	54
rect	117	54	118	55
rect	117	56	118	57
rect	117	57	118	58
rect	117	59	118	60
rect	117	60	118	61
rect	117	62	118	63
rect	117	63	118	64
rect	117	65	118	66
rect	117	66	118	67
rect	117	68	118	69
rect	117	69	118	70
rect	117	71	118	72
rect	117	72	118	73
rect	117	74	118	75
rect	117	75	118	76
rect	117	77	118	78
rect	117	78	118	79
rect	117	80	118	81
rect	117	81	118	82
rect	117	83	118	84
rect	117	84	118	85
rect	117	86	118	87
rect	117	87	118	88
rect	117	89	118	90
rect	117	90	118	91
rect	117	92	118	93
rect	117	93	118	94
rect	117	95	118	96
rect	117	96	118	97
rect	117	98	118	99
rect	117	99	118	100
rect	117	101	118	102
rect	117	102	118	103
rect	117	104	118	105
rect	117	105	118	106
rect	117	107	118	108
rect	117	108	118	109
rect	117	203	118	204
rect	117	204	118	205
rect	117	206	118	207
rect	117	207	118	208
rect	117	209	118	210
rect	117	210	118	211
rect	117	212	118	213
rect	117	213	118	214
rect	117	257	118	258
rect	117	258	118	259
rect	117	260	118	261
rect	117	261	118	262
rect	117	284	118	285
rect	117	285	118	286
rect	117	287	118	288
rect	117	288	118	289
rect	126	134	127	135
rect	126	135	127	136
rect	126	137	127	138
rect	126	138	127	139
rect	126	140	127	141
rect	126	141	127	142
rect	126	143	127	144
rect	126	144	127	145
rect	126	146	127	147
rect	126	147	127	148
rect	126	224	127	225
rect	126	225	127	226
rect	126	311	127	312
rect	126	312	127	313
rect	126	314	127	315
rect	126	315	127	316
rect	126	323	127	324
rect	126	324	127	325
rect	126	326	127	327
rect	126	327	127	328
rect	126	329	127	330
rect	126	330	127	331
rect	126	332	127	333
rect	126	333	127	334
rect	126	335	127	336
rect	126	336	127	337
rect	126	338	127	339
rect	126	339	127	340
rect	126	341	127	342
rect	126	342	127	343
rect	126	344	127	345
rect	126	345	127	346
rect	126	347	127	348
rect	126	348	127	349
rect	128	2	129	3
rect	128	3	129	4
rect	128	5	129	6
rect	128	6	129	7
rect	128	8	129	9
rect	128	9	129	10
rect	128	29	129	30
rect	128	30	129	31
rect	128	32	129	33
rect	128	33	129	34
rect	128	35	129	36
rect	128	36	129	37
rect	128	62	129	63
rect	128	63	129	64
rect	128	113	129	114
rect	128	114	129	115
rect	128	116	129	117
rect	128	117	129	118
rect	128	119	129	120
rect	128	120	129	121
rect	128	122	129	123
rect	128	123	129	124
rect	128	125	129	126
rect	128	126	129	127
rect	128	128	129	129
rect	128	129	129	130
rect	128	131	129	132
rect	128	132	129	133
rect	128	134	129	135
rect	128	135	129	136
rect	128	137	129	138
rect	128	138	129	139
rect	128	140	129	141
rect	128	141	129	142
rect	128	143	129	144
rect	128	144	129	145
rect	128	146	129	147
rect	128	147	129	148
rect	128	149	129	150
rect	128	150	129	151
rect	128	152	129	153
rect	128	153	129	154
rect	128	155	129	156
rect	128	156	129	157
rect	128	158	129	159
rect	128	159	129	160
rect	128	161	129	162
rect	128	162	129	163
rect	128	164	129	165
rect	128	165	129	166
rect	128	167	129	168
rect	128	168	129	169
rect	128	170	129	171
rect	128	171	129	172
rect	128	173	129	174
rect	128	174	129	175
rect	128	176	129	177
rect	128	177	129	178
rect	128	179	129	180
rect	128	180	129	181
rect	128	182	129	183
rect	128	183	129	184
rect	128	185	129	186
rect	128	186	129	187
rect	128	188	129	189
rect	128	189	129	190
rect	128	191	129	192
rect	128	192	129	193
rect	128	194	129	195
rect	128	195	129	196
rect	128	197	129	198
rect	128	198	129	199
rect	128	200	129	201
rect	128	201	129	202
rect	128	203	129	204
rect	128	204	129	205
rect	128	206	129	207
rect	128	207	129	208
rect	128	209	129	210
rect	128	210	129	211
rect	128	212	129	213
rect	128	213	129	214
rect	128	215	129	216
rect	128	216	129	217
rect	128	218	129	219
rect	128	219	129	220
rect	128	221	129	222
rect	128	222	129	223
rect	128	224	129	225
rect	128	225	129	226
rect	128	227	129	228
rect	128	228	129	229
rect	128	230	129	231
rect	128	231	129	232
rect	128	233	129	234
rect	128	234	129	235
rect	128	236	129	237
rect	128	237	129	238
rect	128	239	129	240
rect	128	240	129	241
rect	128	242	129	243
rect	128	243	129	244
rect	128	245	129	246
rect	128	246	129	247
rect	128	248	129	249
rect	128	249	129	250
rect	128	251	129	252
rect	128	252	129	253
rect	128	254	129	255
rect	128	255	129	256
rect	128	257	129	258
rect	128	258	129	259
rect	128	260	129	261
rect	128	261	129	262
rect	128	263	129	264
rect	128	264	129	265
rect	128	266	129	267
rect	128	267	129	268
rect	128	269	129	270
rect	128	270	129	271
rect	128	272	129	273
rect	128	273	129	274
rect	128	275	129	276
rect	128	276	129	277
rect	128	278	129	279
rect	128	279	129	280
rect	128	281	129	282
rect	128	282	129	283
rect	128	284	129	285
rect	128	285	129	286
rect	128	287	129	288
rect	128	288	129	289
rect	128	290	129	291
rect	128	291	129	292
rect	128	293	129	294
rect	128	294	129	295
rect	128	296	129	297
rect	128	297	129	298
rect	128	299	129	300
rect	128	300	129	301
rect	128	302	129	303
rect	128	303	129	304
rect	128	305	129	306
rect	128	306	129	307
rect	128	308	129	309
rect	128	309	129	310
rect	128	311	129	312
rect	128	312	129	313
rect	128	314	129	315
rect	128	315	129	316
rect	128	317	129	318
rect	128	318	129	319
rect	128	320	129	321
rect	128	321	129	322
rect	128	323	129	324
rect	128	324	129	325
rect	128	326	129	327
rect	128	327	129	328
rect	128	329	129	330
rect	128	330	129	331
rect	128	332	129	333
rect	128	333	129	334
rect	137	68	138	69
rect	137	69	138	70
rect	137	71	138	72
rect	137	72	138	73
rect	137	74	138	75
rect	137	75	138	76
rect	137	77	138	78
rect	137	78	138	79
rect	137	80	138	81
rect	137	81	138	82
rect	137	83	138	84
rect	137	84	138	85
rect	137	86	138	87
rect	137	87	138	88
rect	137	128	138	129
rect	137	129	138	130
rect	137	131	138	132
rect	137	132	138	133
rect	137	134	138	135
rect	137	135	138	136
rect	137	137	138	138
rect	137	138	138	139
rect	137	140	138	141
rect	137	141	138	142
rect	137	143	138	144
rect	137	144	138	145
rect	137	146	138	147
rect	137	147	138	148
rect	137	149	138	150
rect	137	150	138	151
rect	137	152	138	153
rect	137	153	138	154
rect	137	155	138	156
rect	137	156	138	157
rect	137	158	138	159
rect	137	159	138	160
rect	137	161	138	162
rect	137	162	138	163
rect	137	164	138	165
rect	137	165	138	166
rect	137	167	138	168
rect	137	168	138	169
rect	137	170	138	171
rect	137	171	138	172
rect	137	173	138	174
rect	137	174	138	175
rect	137	176	138	177
rect	137	177	138	178
rect	137	179	138	180
rect	137	180	138	181
rect	137	248	138	249
rect	137	249	138	250
rect	137	251	138	252
rect	137	252	138	253
rect	139	62	140	63
rect	139	63	140	64
rect	139	65	140	66
rect	139	66	140	67
rect	139	68	140	69
rect	139	69	140	70
rect	139	71	140	72
rect	139	72	140	73
rect	139	74	140	75
rect	139	75	140	76
rect	139	77	140	78
rect	139	78	140	79
rect	139	80	140	81
rect	139	81	140	82
rect	139	83	140	84
rect	139	84	140	85
rect	139	86	140	87
rect	139	87	140	88
rect	139	89	140	90
rect	139	90	140	91
rect	139	92	140	93
rect	139	93	140	94
rect	139	95	140	96
rect	139	96	140	97
rect	139	98	140	99
rect	139	99	140	100
rect	139	101	140	102
rect	139	102	140	103
rect	139	104	140	105
rect	139	105	140	106
rect	139	107	140	108
rect	139	108	140	109
rect	139	110	140	111
rect	139	111	140	112
rect	139	113	140	114
rect	139	114	140	115
rect	139	116	140	117
rect	139	117	140	118
rect	139	119	140	120
rect	139	120	140	121
rect	139	122	140	123
rect	139	123	140	124
rect	139	125	140	126
rect	139	126	140	127
rect	139	128	140	129
rect	139	129	140	130
rect	139	131	140	132
rect	139	132	140	133
rect	139	134	140	135
rect	139	135	140	136
rect	139	137	140	138
rect	139	138	140	139
rect	139	140	140	141
rect	139	141	140	142
rect	139	143	140	144
rect	139	144	140	145
rect	139	146	140	147
rect	139	147	140	148
rect	139	149	140	150
rect	139	150	140	151
rect	139	152	140	153
rect	139	153	140	154
rect	139	155	140	156
rect	139	156	140	157
rect	139	158	140	159
rect	139	159	140	160
rect	139	161	140	162
rect	139	162	140	163
rect	139	164	140	165
rect	139	165	140	166
rect	139	167	140	168
rect	139	168	140	169
rect	139	170	140	171
rect	139	171	140	172
rect	139	173	140	174
rect	139	174	140	175
rect	139	176	140	177
rect	139	177	140	178
rect	139	179	140	180
rect	139	180	140	181
rect	139	182	140	183
rect	139	183	140	184
rect	139	185	140	186
rect	139	186	140	187
rect	139	188	140	189
rect	139	189	140	190
rect	139	191	140	192
rect	139	192	140	193
rect	139	194	140	195
rect	139	195	140	196
rect	139	197	140	198
rect	139	198	140	199
rect	139	200	140	201
rect	139	201	140	202
rect	139	203	140	204
rect	139	204	140	205
rect	139	206	140	207
rect	139	207	140	208
rect	139	209	140	210
rect	139	210	140	211
rect	139	212	140	213
rect	139	213	140	214
rect	139	215	140	216
rect	139	216	140	217
rect	139	218	140	219
rect	139	219	140	220
rect	139	221	140	222
rect	139	222	140	223
rect	139	224	140	225
rect	139	225	140	226
rect	139	227	140	228
rect	139	228	140	229
rect	139	230	140	231
rect	139	231	140	232
rect	139	233	140	234
rect	139	234	140	235
rect	139	236	140	237
rect	139	237	140	238
rect	139	239	140	240
rect	139	240	140	241
rect	139	242	140	243
rect	139	243	140	244
rect	139	245	140	246
rect	139	246	140	247
rect	139	248	140	249
rect	139	249	140	250
rect	139	251	140	252
rect	139	252	140	253
rect	139	254	140	255
rect	139	255	140	256
rect	139	257	140	258
rect	139	258	140	259
rect	139	260	140	261
rect	139	261	140	262
rect	139	263	140	264
rect	139	264	140	265
rect	139	266	140	267
rect	139	267	140	268
rect	139	269	140	270
rect	139	270	140	271
rect	139	272	140	273
rect	139	273	140	274
rect	139	275	140	276
rect	139	276	140	277
rect	139	278	140	279
rect	139	279	140	280
rect	139	281	140	282
rect	139	282	140	283
rect	139	284	140	285
rect	139	285	140	286
rect	139	308	140	309
rect	139	309	140	310
rect	139	311	140	312
rect	139	312	140	313
rect	141	50	142	51
rect	141	51	142	52
rect	141	53	142	54
rect	141	54	142	55
rect	141	56	142	57
rect	141	57	142	58
rect	141	59	142	60
rect	141	60	142	61
rect	141	62	142	63
rect	141	63	142	64
rect	141	65	142	66
rect	141	66	142	67
rect	141	68	142	69
rect	141	69	142	70
rect	141	71	142	72
rect	141	72	142	73
rect	141	74	142	75
rect	141	75	142	76
rect	141	77	142	78
rect	141	78	142	79
rect	141	80	142	81
rect	141	81	142	82
rect	141	83	142	84
rect	141	84	142	85
rect	141	86	142	87
rect	141	87	142	88
rect	141	89	142	90
rect	141	90	142	91
rect	141	92	142	93
rect	141	93	142	94
rect	141	95	142	96
rect	141	96	142	97
rect	141	98	142	99
rect	141	99	142	100
rect	141	101	142	102
rect	141	102	142	103
rect	141	104	142	105
rect	141	105	142	106
rect	141	107	142	108
rect	141	108	142	109
rect	141	110	142	111
rect	141	111	142	112
rect	141	113	142	114
rect	141	114	142	115
rect	141	116	142	117
rect	141	117	142	118
rect	141	119	142	120
rect	141	120	142	121
rect	141	122	142	123
rect	141	123	142	124
rect	141	125	142	126
rect	141	126	142	127
rect	141	128	142	129
rect	141	129	142	130
rect	141	131	142	132
rect	141	132	142	133
rect	141	134	142	135
rect	141	135	142	136
rect	141	137	142	138
rect	141	138	142	139
rect	141	140	142	141
rect	141	141	142	142
rect	141	143	142	144
rect	141	144	142	145
rect	141	146	142	147
rect	141	147	142	148
rect	141	149	142	150
rect	141	150	142	151
rect	141	152	142	153
rect	141	153	142	154
rect	141	155	142	156
rect	141	156	142	157
rect	141	158	142	159
rect	141	159	142	160
rect	141	161	142	162
rect	141	162	142	163
rect	141	164	142	165
rect	141	165	142	166
rect	141	167	142	168
rect	141	168	142	169
rect	141	170	142	171
rect	141	171	142	172
rect	141	173	142	174
rect	141	174	142	175
rect	141	176	142	177
rect	141	177	142	178
rect	141	179	142	180
rect	141	180	142	181
rect	141	182	142	183
rect	141	183	142	184
rect	141	185	142	186
rect	141	186	142	187
rect	141	188	142	189
rect	141	189	142	190
rect	141	191	142	192
rect	141	192	142	193
rect	141	194	142	195
rect	141	195	142	196
rect	141	197	142	198
rect	141	198	142	199
rect	141	200	142	201
rect	141	201	142	202
rect	141	203	142	204
rect	141	204	142	205
rect	141	206	142	207
rect	141	207	142	208
rect	141	209	142	210
rect	141	210	142	211
rect	141	212	142	213
rect	141	213	142	214
rect	141	215	142	216
rect	141	216	142	217
rect	141	218	142	219
rect	141	219	142	220
rect	141	221	142	222
rect	141	222	142	223
rect	141	224	142	225
rect	141	225	142	226
rect	141	227	142	228
rect	141	228	142	229
rect	141	230	142	231
rect	141	231	142	232
rect	141	233	142	234
rect	141	234	142	235
rect	141	236	142	237
rect	141	237	142	238
rect	141	239	142	240
rect	141	240	142	241
rect	141	242	142	243
rect	141	243	142	244
rect	141	245	142	246
rect	141	246	142	247
rect	141	248	142	249
rect	141	249	142	250
rect	141	251	142	252
rect	141	252	142	253
rect	141	254	142	255
rect	141	255	142	256
rect	141	257	142	258
rect	141	258	142	259
rect	141	260	142	261
rect	141	261	142	262
rect	141	263	142	264
rect	141	264	142	265
rect	141	266	142	267
rect	141	267	142	268
rect	141	269	142	270
rect	141	270	142	271
rect	141	272	142	273
rect	141	273	142	274
rect	141	275	142	276
rect	141	276	142	277
rect	141	278	142	279
rect	141	279	142	280
rect	141	281	142	282
rect	141	282	142	283
rect	141	284	142	285
rect	141	285	142	286
rect	141	287	142	288
rect	141	288	142	289
rect	141	290	142	291
rect	141	291	142	292
rect	141	293	142	294
rect	141	294	142	295
rect	141	302	142	303
rect	141	303	142	304
rect	141	305	142	306
rect	141	306	142	307
rect	141	308	142	309
rect	141	309	142	310
rect	150	176	151	177
rect	150	177	151	178
rect	150	179	151	180
rect	150	180	151	181
rect	150	182	151	183
rect	150	183	151	184
rect	150	185	151	186
rect	150	186	151	187
rect	150	188	151	189
rect	150	189	151	190
rect	152	140	153	141
rect	152	141	153	142
rect	152	143	153	144
rect	152	144	153	145
rect	152	146	153	147
rect	152	147	153	148
rect	152	149	153	150
rect	152	150	153	151
rect	152	152	153	153
rect	152	153	153	154
rect	152	155	153	156
rect	152	156	153	157
rect	152	158	153	159
rect	152	159	153	160
rect	152	161	153	162
rect	152	162	153	163
rect	152	164	153	165
rect	152	165	153	166
rect	152	167	153	168
rect	152	168	153	169
rect	152	170	153	171
rect	152	171	153	172
rect	152	173	153	174
rect	152	174	153	175
rect	152	176	153	177
rect	152	177	153	178
rect	152	179	153	180
rect	152	180	153	181
rect	152	182	153	183
rect	152	183	153	184
rect	152	185	153	186
rect	152	186	153	187
rect	154	116	155	117
rect	154	117	155	118
rect	154	134	155	135
rect	154	135	155	136
rect	154	137	155	138
rect	154	138	155	139
rect	154	140	155	141
rect	154	141	155	142
rect	154	143	155	144
rect	154	144	155	145
rect	154	146	155	147
rect	154	147	155	148
rect	154	149	155	150
rect	154	150	155	151
rect	154	152	155	153
rect	154	153	155	154
rect	154	155	155	156
rect	154	156	155	157
rect	154	158	155	159
rect	154	159	155	160
rect	154	161	155	162
rect	154	162	155	163
rect	154	164	155	165
rect	154	165	155	166
rect	154	167	155	168
rect	154	168	155	169
rect	154	170	155	171
rect	154	171	155	172
rect	154	173	155	174
rect	154	174	155	175
rect	154	176	155	177
rect	154	177	155	178
rect	154	179	155	180
rect	154	180	155	181
rect	154	182	155	183
rect	154	183	155	184
rect	154	185	155	186
rect	154	186	155	187
rect	154	188	155	189
rect	154	189	155	190
rect	154	191	155	192
rect	154	192	155	193
rect	154	194	155	195
rect	154	195	155	196
rect	154	197	155	198
rect	154	198	155	199
rect	154	200	155	201
rect	154	201	155	202
rect	154	203	155	204
rect	154	204	155	205
rect	154	206	155	207
rect	154	207	155	208
rect	154	209	155	210
rect	154	210	155	211
rect	154	212	155	213
rect	154	213	155	214
rect	154	215	155	216
rect	154	216	155	217
rect	154	218	155	219
rect	154	219	155	220
rect	154	221	155	222
rect	154	222	155	223
rect	154	224	155	225
rect	154	225	155	226
rect	154	227	155	228
rect	154	228	155	229
rect	154	230	155	231
rect	154	231	155	232
rect	154	233	155	234
rect	154	234	155	235
rect	154	236	155	237
rect	154	237	155	238
rect	154	239	155	240
rect	154	240	155	241
rect	154	242	155	243
rect	154	243	155	244
rect	154	245	155	246
rect	154	246	155	247
rect	154	248	155	249
rect	154	249	155	250
rect	154	251	155	252
rect	154	252	155	253
rect	154	254	155	255
rect	154	255	155	256
rect	154	257	155	258
rect	154	258	155	259
rect	154	260	155	261
rect	154	261	155	262
rect	154	263	155	264
rect	154	264	155	265
rect	154	266	155	267
rect	154	267	155	268
rect	154	269	155	270
rect	154	270	155	271
rect	154	272	155	273
rect	154	273	155	274
rect	154	275	155	276
rect	154	276	155	277
rect	154	278	155	279
rect	154	279	155	280
rect	154	281	155	282
rect	154	282	155	283
rect	154	284	155	285
rect	154	285	155	286
rect	154	287	155	288
rect	154	288	155	289
rect	154	290	155	291
rect	154	291	155	292
rect	154	293	155	294
rect	154	294	155	295
rect	154	296	155	297
rect	154	297	155	298
rect	154	299	155	300
rect	154	300	155	301
rect	154	302	155	303
rect	154	303	155	304
rect	154	304	155	305
rect	154	305	155	306
rect	154	306	155	307
rect	154	308	155	309
rect	154	309	155	310
rect	154	311	155	312
rect	154	312	155	313
rect	154	314	155	315
rect	154	315	155	316
rect	154	317	155	318
rect	154	318	155	319
rect	154	320	155	321
rect	154	321	155	322
rect	154	323	155	324
rect	154	324	155	325
rect	154	326	155	327
rect	154	327	155	328
rect	154	329	155	330
rect	154	330	155	331
rect	154	332	155	333
rect	154	333	155	334
rect	154	335	155	336
rect	154	336	155	337
rect	154	337	155	338
rect	154	338	155	339
rect	154	339	155	340
rect	154	341	155	342
rect	154	342	155	343
rect	154	344	155	345
rect	154	345	155	346
rect	156	89	157	90
rect	156	90	157	91
rect	156	92	157	93
rect	156	93	157	94
rect	156	95	157	96
rect	156	96	157	97
rect	156	98	157	99
rect	156	99	157	100
rect	156	101	157	102
rect	156	102	157	103
rect	156	104	157	105
rect	156	105	157	106
rect	156	107	157	108
rect	156	108	157	109
rect	156	110	157	111
rect	156	111	157	112
rect	156	113	157	114
rect	156	114	157	115
rect	156	116	157	117
rect	156	117	157	118
rect	156	119	157	120
rect	156	120	157	121
rect	156	122	157	123
rect	156	123	157	124
rect	156	125	157	126
rect	156	126	157	127
rect	156	128	157	129
rect	156	129	157	130
rect	156	131	157	132
rect	156	132	157	133
rect	156	134	157	135
rect	156	135	157	136
rect	156	137	157	138
rect	156	138	157	139
rect	156	140	157	141
rect	156	141	157	142
rect	156	143	157	144
rect	156	144	157	145
rect	156	146	157	147
rect	156	147	157	148
rect	156	149	157	150
rect	156	150	157	151
rect	156	152	157	153
rect	156	153	157	154
rect	156	155	157	156
rect	156	156	157	157
rect	156	158	157	159
rect	156	159	157	160
rect	156	161	157	162
rect	156	162	157	163
rect	156	164	157	165
rect	156	165	157	166
rect	156	167	157	168
rect	156	168	157	169
rect	156	170	157	171
rect	156	171	157	172
rect	156	173	157	174
rect	156	174	157	175
rect	156	176	157	177
rect	156	177	157	178
rect	156	179	157	180
rect	156	180	157	181
rect	156	182	157	183
rect	156	183	157	184
rect	156	185	157	186
rect	156	186	157	187
rect	156	188	157	189
rect	156	189	157	190
rect	156	191	157	192
rect	156	192	157	193
rect	156	194	157	195
rect	156	195	157	196
rect	156	197	157	198
rect	156	198	157	199
rect	156	200	157	201
rect	156	201	157	202
rect	156	203	157	204
rect	156	204	157	205
rect	156	206	157	207
rect	156	207	157	208
rect	156	209	157	210
rect	156	210	157	211
rect	156	212	157	213
rect	156	213	157	214
rect	156	215	157	216
rect	156	216	157	217
rect	156	218	157	219
rect	156	219	157	220
rect	156	221	157	222
rect	156	222	157	223
rect	156	224	157	225
rect	156	225	157	226
rect	156	227	157	228
rect	156	228	157	229
rect	156	230	157	231
rect	156	231	157	232
rect	156	233	157	234
rect	156	234	157	235
rect	156	236	157	237
rect	156	237	157	238
rect	156	239	157	240
rect	156	240	157	241
rect	156	242	157	243
rect	156	243	157	244
rect	156	245	157	246
rect	156	246	157	247
rect	156	248	157	249
rect	156	249	157	250
rect	156	251	157	252
rect	156	252	157	253
rect	156	254	157	255
rect	156	255	157	256
rect	156	257	157	258
rect	156	258	157	259
rect	156	260	157	261
rect	156	261	157	262
rect	156	263	157	264
rect	156	264	157	265
rect	156	266	157	267
rect	156	267	157	268
rect	156	269	157	270
rect	156	270	157	271
rect	156	272	157	273
rect	156	273	157	274
rect	156	275	157	276
rect	156	276	157	277
rect	156	278	157	279
rect	156	279	157	280
rect	156	281	157	282
rect	156	282	157	283
rect	156	284	157	285
rect	156	285	157	286
rect	156	287	157	288
rect	156	288	157	289
rect	156	290	157	291
rect	156	291	157	292
rect	156	293	157	294
rect	156	294	157	295
rect	156	332	157	333
rect	156	333	157	334
rect	156	335	157	336
rect	156	336	157	337
rect	156	341	157	342
rect	156	342	157	343
rect	156	344	157	345
rect	156	345	157	346
rect	156	347	157	348
rect	156	348	157	349
rect	156	350	157	351
rect	156	351	157	352
rect	156	353	157	354
rect	156	354	157	355
rect	156	356	157	357
rect	156	357	157	358
rect	156	359	157	360
rect	156	360	157	361
rect	156	362	157	363
rect	156	363	157	364
rect	156	365	157	366
rect	156	366	157	367
rect	156	368	157	369
rect	156	369	157	370
rect	158	11	159	12
rect	158	12	159	13
rect	158	14	159	15
rect	158	15	159	16
rect	158	83	159	84
rect	158	84	159	85
rect	158	86	159	87
rect	158	87	159	88
rect	158	89	159	90
rect	158	90	159	91
rect	158	92	159	93
rect	158	93	159	94
rect	158	95	159	96
rect	158	96	159	97
rect	158	98	159	99
rect	158	99	159	100
rect	158	101	159	102
rect	158	102	159	103
rect	158	104	159	105
rect	158	105	159	106
rect	158	107	159	108
rect	158	108	159	109
rect	158	110	159	111
rect	158	111	159	112
rect	158	113	159	114
rect	158	114	159	115
rect	158	116	159	117
rect	158	117	159	118
rect	158	119	159	120
rect	158	120	159	121
rect	158	122	159	123
rect	158	123	159	124
rect	158	125	159	126
rect	158	126	159	127
rect	158	128	159	129
rect	158	129	159	130
rect	158	131	159	132
rect	158	132	159	133
rect	158	134	159	135
rect	158	135	159	136
rect	158	137	159	138
rect	158	138	159	139
rect	158	140	159	141
rect	158	141	159	142
rect	158	143	159	144
rect	158	144	159	145
rect	158	146	159	147
rect	158	147	159	148
rect	158	149	159	150
rect	158	150	159	151
rect	158	152	159	153
rect	158	153	159	154
rect	158	155	159	156
rect	158	156	159	157
rect	158	158	159	159
rect	158	159	159	160
rect	158	161	159	162
rect	158	162	159	163
rect	158	164	159	165
rect	158	165	159	166
rect	158	167	159	168
rect	158	168	159	169
rect	158	170	159	171
rect	158	171	159	172
rect	158	173	159	174
rect	158	174	159	175
rect	158	176	159	177
rect	158	177	159	178
rect	158	179	159	180
rect	158	180	159	181
rect	158	182	159	183
rect	158	183	159	184
rect	158	185	159	186
rect	158	186	159	187
rect	158	188	159	189
rect	158	189	159	190
rect	158	191	159	192
rect	158	192	159	193
rect	158	194	159	195
rect	158	195	159	196
rect	158	197	159	198
rect	158	198	159	199
rect	158	200	159	201
rect	158	201	159	202
rect	158	203	159	204
rect	158	204	159	205
rect	158	206	159	207
rect	158	207	159	208
rect	158	209	159	210
rect	158	210	159	211
rect	158	212	159	213
rect	158	213	159	214
rect	158	215	159	216
rect	158	216	159	217
rect	158	218	159	219
rect	158	219	159	220
rect	158	221	159	222
rect	158	222	159	223
rect	158	224	159	225
rect	158	225	159	226
rect	158	227	159	228
rect	158	228	159	229
rect	158	230	159	231
rect	158	231	159	232
rect	158	233	159	234
rect	158	234	159	235
rect	158	236	159	237
rect	158	237	159	238
rect	158	239	159	240
rect	158	240	159	241
rect	158	242	159	243
rect	158	243	159	244
rect	158	245	159	246
rect	158	246	159	247
rect	158	248	159	249
rect	158	249	159	250
rect	158	251	159	252
rect	158	252	159	253
rect	158	254	159	255
rect	158	255	159	256
rect	158	257	159	258
rect	158	258	159	259
rect	158	260	159	261
rect	158	261	159	262
rect	158	263	159	264
rect	158	264	159	265
rect	158	266	159	267
rect	158	267	159	268
rect	158	269	159	270
rect	158	270	159	271
rect	158	272	159	273
rect	158	273	159	274
rect	158	275	159	276
rect	158	276	159	277
rect	158	278	159	279
rect	158	279	159	280
rect	158	320	159	321
rect	158	321	159	322
rect	158	323	159	324
rect	158	324	159	325
rect	158	326	159	327
rect	158	327	159	328
rect	158	329	159	330
rect	158	330	159	331
rect	158	332	159	333
rect	158	333	159	334
rect	158	335	159	336
rect	158	336	159	337
rect	158	338	159	339
rect	158	339	159	340
rect	158	341	159	342
rect	158	342	159	343
rect	158	344	159	345
rect	158	345	159	346
rect	158	347	159	348
rect	158	348	159	349
rect	167	47	168	48
rect	167	48	168	49
rect	167	50	168	51
rect	167	51	168	52
rect	167	53	168	54
rect	167	54	168	55
rect	167	56	168	57
rect	167	57	168	58
rect	167	59	168	60
rect	167	60	168	61
rect	167	62	168	63
rect	167	63	168	64
rect	167	65	168	66
rect	167	66	168	67
rect	167	68	168	69
rect	167	69	168	70
rect	167	71	168	72
rect	167	72	168	73
rect	167	74	168	75
rect	167	75	168	76
rect	167	77	168	78
rect	167	78	168	79
rect	167	80	168	81
rect	167	81	168	82
rect	167	83	168	84
rect	167	84	168	85
rect	167	86	168	87
rect	167	87	168	88
rect	167	89	168	90
rect	167	90	168	91
rect	167	92	168	93
rect	167	93	168	94
rect	167	95	168	96
rect	167	96	168	97
rect	167	98	168	99
rect	167	99	168	100
rect	167	101	168	102
rect	167	102	168	103
rect	167	104	168	105
rect	167	105	168	106
rect	167	107	168	108
rect	167	108	168	109
rect	167	110	168	111
rect	167	111	168	112
rect	167	113	168	114
rect	167	114	168	115
rect	167	116	168	117
rect	167	117	168	118
rect	167	119	168	120
rect	167	120	168	121
rect	167	122	168	123
rect	167	123	168	124
rect	167	125	168	126
rect	167	126	168	127
rect	167	128	168	129
rect	167	129	168	130
rect	167	131	168	132
rect	167	132	168	133
rect	167	134	168	135
rect	167	135	168	136
rect	167	137	168	138
rect	167	138	168	139
rect	167	140	168	141
rect	167	141	168	142
rect	167	143	168	144
rect	167	144	168	145
rect	167	146	168	147
rect	167	147	168	148
rect	167	149	168	150
rect	167	150	168	151
rect	167	152	168	153
rect	167	153	168	154
rect	167	155	168	156
rect	167	156	168	157
rect	167	158	168	159
rect	167	159	168	160
rect	167	161	168	162
rect	167	162	168	163
rect	167	164	168	165
rect	167	165	168	166
rect	167	167	168	168
rect	167	168	168	169
rect	167	170	168	171
rect	167	171	168	172
rect	167	173	168	174
rect	167	174	168	175
rect	167	176	168	177
rect	167	177	168	178
rect	167	179	168	180
rect	167	180	168	181
rect	167	182	168	183
rect	167	183	168	184
rect	167	185	168	186
rect	167	186	168	187
rect	167	188	168	189
rect	167	189	168	190
rect	167	191	168	192
rect	167	192	168	193
rect	167	194	168	195
rect	167	195	168	196
rect	167	197	168	198
rect	167	198	168	199
rect	167	200	168	201
rect	167	201	168	202
rect	167	203	168	204
rect	167	204	168	205
rect	167	206	168	207
rect	167	207	168	208
rect	167	209	168	210
rect	167	210	168	211
rect	167	212	168	213
rect	167	213	168	214
rect	167	215	168	216
rect	167	216	168	217
rect	167	218	168	219
rect	167	219	168	220
rect	167	221	168	222
rect	167	222	168	223
rect	167	224	168	225
rect	167	225	168	226
rect	167	227	168	228
rect	167	228	168	229
rect	167	230	168	231
rect	167	231	168	232
rect	167	233	168	234
rect	167	234	168	235
rect	167	236	168	237
rect	167	237	168	238
rect	167	239	168	240
rect	167	240	168	241
rect	167	242	168	243
rect	167	243	168	244
rect	167	245	168	246
rect	167	246	168	247
rect	167	248	168	249
rect	167	249	168	250
rect	167	251	168	252
rect	167	252	168	253
rect	167	254	168	255
rect	167	255	168	256
rect	167	257	168	258
rect	167	258	168	259
rect	167	260	168	261
rect	167	261	168	262
rect	167	263	168	264
rect	167	264	168	265
rect	167	266	168	267
rect	167	267	168	268
rect	167	269	168	270
rect	167	270	168	271
rect	167	272	168	273
rect	167	273	168	274
rect	167	275	168	276
rect	167	276	168	277
rect	167	278	168	279
rect	167	279	168	280
rect	167	281	168	282
rect	167	282	168	283
rect	167	284	168	285
rect	167	285	168	286
rect	167	287	168	288
rect	167	288	168	289
rect	167	290	168	291
rect	167	291	168	292
rect	167	293	168	294
rect	167	294	168	295
rect	167	296	168	297
rect	167	297	168	298
rect	167	299	168	300
rect	167	300	168	301
rect	167	302	168	303
rect	167	303	168	304
rect	167	304	168	305
rect	167	305	168	306
rect	167	306	168	307
rect	167	308	168	309
rect	167	309	168	310
rect	167	311	168	312
rect	167	312	168	313
rect	167	314	168	315
rect	167	315	168	316
rect	167	317	168	318
rect	167	318	168	319
rect	167	320	168	321
rect	167	321	168	322
rect	167	323	168	324
rect	167	324	168	325
rect	167	326	168	327
rect	167	327	168	328
rect	167	328	168	329
rect	167	329	168	330
rect	167	330	168	331
rect	167	332	168	333
rect	167	333	168	334
rect	167	335	168	336
rect	167	336	168	337
rect	167	337	168	338
rect	167	338	168	339
rect	167	339	168	340
rect	167	340	168	341
rect	167	341	168	342
rect	167	342	168	343
rect	167	343	168	344
rect	167	344	168	345
rect	167	345	168	346
rect	167	347	168	348
rect	167	348	168	349
rect	167	350	168	351
rect	167	351	168	352
rect	167	353	168	354
rect	167	354	168	355
rect	167	356	168	357
rect	167	357	168	358
rect	169	44	170	45
rect	169	45	170	46
rect	169	47	170	48
rect	169	48	170	49
rect	169	50	170	51
rect	169	51	170	52
rect	169	53	170	54
rect	169	54	170	55
rect	169	56	170	57
rect	169	57	170	58
rect	169	59	170	60
rect	169	60	170	61
rect	169	62	170	63
rect	169	63	170	64
rect	169	65	170	66
rect	169	66	170	67
rect	169	68	170	69
rect	169	69	170	70
rect	169	71	170	72
rect	169	72	170	73
rect	169	74	170	75
rect	169	75	170	76
rect	169	77	170	78
rect	169	78	170	79
rect	169	80	170	81
rect	169	81	170	82
rect	169	83	170	84
rect	169	84	170	85
rect	169	86	170	87
rect	169	87	170	88
rect	169	89	170	90
rect	169	90	170	91
rect	169	92	170	93
rect	169	93	170	94
rect	169	95	170	96
rect	169	96	170	97
rect	169	98	170	99
rect	169	99	170	100
rect	169	101	170	102
rect	169	102	170	103
rect	169	104	170	105
rect	169	105	170	106
rect	169	107	170	108
rect	169	108	170	109
rect	169	110	170	111
rect	169	111	170	112
rect	169	113	170	114
rect	169	114	170	115
rect	169	116	170	117
rect	169	117	170	118
rect	169	119	170	120
rect	169	120	170	121
rect	169	122	170	123
rect	169	123	170	124
rect	169	125	170	126
rect	169	126	170	127
rect	169	128	170	129
rect	169	129	170	130
rect	169	131	170	132
rect	169	132	170	133
rect	169	134	170	135
rect	169	135	170	136
rect	169	137	170	138
rect	169	138	170	139
rect	169	140	170	141
rect	169	141	170	142
rect	169	143	170	144
rect	169	144	170	145
rect	169	146	170	147
rect	169	147	170	148
rect	169	149	170	150
rect	169	150	170	151
rect	169	152	170	153
rect	169	153	170	154
rect	169	155	170	156
rect	169	156	170	157
rect	169	158	170	159
rect	169	159	170	160
rect	169	161	170	162
rect	169	162	170	163
rect	169	164	170	165
rect	169	165	170	166
rect	169	167	170	168
rect	169	168	170	169
rect	169	170	170	171
rect	169	171	170	172
rect	169	173	170	174
rect	169	174	170	175
rect	169	176	170	177
rect	169	177	170	178
rect	169	179	170	180
rect	169	180	170	181
rect	169	182	170	183
rect	169	183	170	184
rect	169	185	170	186
rect	169	186	170	187
rect	169	188	170	189
rect	169	189	170	190
rect	169	191	170	192
rect	169	192	170	193
rect	169	194	170	195
rect	169	195	170	196
rect	169	197	170	198
rect	169	198	170	199
rect	169	200	170	201
rect	169	201	170	202
rect	169	203	170	204
rect	169	204	170	205
rect	169	206	170	207
rect	169	207	170	208
rect	169	209	170	210
rect	169	210	170	211
rect	169	212	170	213
rect	169	213	170	214
rect	169	215	170	216
rect	169	216	170	217
rect	169	218	170	219
rect	169	219	170	220
rect	169	221	170	222
rect	169	222	170	223
rect	169	224	170	225
rect	169	225	170	226
rect	169	227	170	228
rect	169	228	170	229
rect	171	5	172	6
rect	171	6	172	7
rect	171	8	172	9
rect	171	9	172	10
rect	171	11	172	12
rect	171	12	172	13
rect	171	14	172	15
rect	171	15	172	16
rect	171	17	172	18
rect	171	18	172	19
rect	171	20	172	21
rect	171	21	172	22
rect	171	23	172	24
rect	171	24	172	25
rect	171	26	172	27
rect	171	27	172	28
rect	171	29	172	30
rect	171	30	172	31
rect	171	32	172	33
rect	171	33	172	34
rect	171	35	172	36
rect	171	36	172	37
rect	171	38	172	39
rect	171	39	172	40
rect	171	41	172	42
rect	171	42	172	43
rect	171	44	172	45
rect	171	45	172	46
rect	171	47	172	48
rect	171	48	172	49
rect	171	50	172	51
rect	171	51	172	52
rect	171	53	172	54
rect	171	54	172	55
rect	171	56	172	57
rect	171	57	172	58
rect	171	59	172	60
rect	171	60	172	61
rect	171	62	172	63
rect	171	63	172	64
rect	171	65	172	66
rect	171	66	172	67
rect	171	68	172	69
rect	171	69	172	70
rect	171	71	172	72
rect	171	72	172	73
rect	171	74	172	75
rect	171	75	172	76
rect	171	86	172	87
rect	171	87	172	88
rect	171	149	172	150
rect	171	150	172	151
rect	171	152	172	153
rect	171	153	172	154
rect	171	155	172	156
rect	171	156	172	157
rect	171	158	172	159
rect	171	159	172	160
rect	171	161	172	162
rect	171	162	172	163
rect	171	164	172	165
rect	171	165	172	166
rect	171	167	172	168
rect	171	168	172	169
rect	171	314	172	315
rect	171	315	172	316
rect	171	317	172	318
rect	171	318	172	319
rect	180	92	181	93
rect	180	93	181	94
rect	180	95	181	96
rect	180	96	181	97
rect	180	98	181	99
rect	180	99	181	100
rect	180	101	181	102
rect	180	102	181	103
rect	180	104	181	105
rect	180	105	181	106
rect	180	107	181	108
rect	180	108	181	109
rect	180	110	181	111
rect	180	111	181	112
rect	180	113	181	114
rect	180	114	181	115
rect	180	116	181	117
rect	180	117	181	118
rect	180	119	181	120
rect	180	120	181	121
rect	180	122	181	123
rect	180	123	181	124
rect	180	125	181	126
rect	180	126	181	127
rect	180	128	181	129
rect	180	129	181	130
rect	180	131	181	132
rect	180	132	181	133
rect	180	134	181	135
rect	180	135	181	136
rect	180	137	181	138
rect	180	138	181	139
rect	180	140	181	141
rect	180	141	181	142
rect	180	143	181	144
rect	180	144	181	145
rect	180	146	181	147
rect	180	147	181	148
rect	180	149	181	150
rect	180	150	181	151
rect	180	152	181	153
rect	180	153	181	154
rect	180	155	181	156
rect	180	156	181	157
rect	180	158	181	159
rect	180	159	181	160
rect	180	161	181	162
rect	180	162	181	163
rect	180	164	181	165
rect	180	165	181	166
rect	180	167	181	168
rect	180	168	181	169
rect	180	170	181	171
rect	180	171	181	172
rect	180	173	181	174
rect	180	174	181	175
rect	180	176	181	177
rect	180	177	181	178
rect	180	179	181	180
rect	180	180	181	181
rect	180	182	181	183
rect	180	183	181	184
rect	180	185	181	186
rect	180	186	181	187
rect	180	188	181	189
rect	180	189	181	190
rect	180	191	181	192
rect	180	192	181	193
rect	180	194	181	195
rect	180	195	181	196
rect	180	197	181	198
rect	180	198	181	199
rect	180	200	181	201
rect	180	201	181	202
rect	180	203	181	204
rect	180	204	181	205
rect	180	206	181	207
rect	180	207	181	208
rect	180	209	181	210
rect	180	210	181	211
rect	180	212	181	213
rect	180	213	181	214
rect	180	215	181	216
rect	180	216	181	217
rect	180	218	181	219
rect	180	219	181	220
rect	180	221	181	222
rect	180	222	181	223
rect	180	224	181	225
rect	180	225	181	226
rect	180	227	181	228
rect	180	228	181	229
rect	180	230	181	231
rect	180	231	181	232
rect	180	233	181	234
rect	180	234	181	235
rect	180	236	181	237
rect	180	237	181	238
rect	180	239	181	240
rect	180	240	181	241
rect	180	242	181	243
rect	180	243	181	244
rect	180	245	181	246
rect	180	246	181	247
rect	180	248	181	249
rect	180	249	181	250
rect	180	251	181	252
rect	180	252	181	253
rect	180	254	181	255
rect	180	255	181	256
rect	180	257	181	258
rect	180	258	181	259
rect	180	260	181	261
rect	180	261	181	262
rect	180	263	181	264
rect	180	264	181	265
rect	180	266	181	267
rect	180	267	181	268
rect	180	269	181	270
rect	180	270	181	271
rect	180	272	181	273
rect	180	273	181	274
rect	180	275	181	276
rect	180	276	181	277
rect	180	278	181	279
rect	180	279	181	280
rect	180	281	181	282
rect	180	282	181	283
rect	180	284	181	285
rect	180	285	181	286
rect	180	287	181	288
rect	180	288	181	289
rect	180	290	181	291
rect	180	291	181	292
rect	180	293	181	294
rect	180	294	181	295
rect	180	296	181	297
rect	180	297	181	298
rect	180	299	181	300
rect	180	300	181	301
rect	180	302	181	303
rect	180	303	181	304
rect	180	304	181	305
rect	180	305	181	306
rect	180	306	181	307
rect	182	77	183	78
rect	182	78	183	79
rect	182	80	183	81
rect	182	81	183	82
rect	182	83	183	84
rect	182	84	183	85
rect	182	86	183	87
rect	182	87	183	88
rect	182	89	183	90
rect	182	90	183	91
rect	182	92	183	93
rect	182	93	183	94
rect	182	95	183	96
rect	182	96	183	97
rect	182	98	183	99
rect	182	99	183	100
rect	182	101	183	102
rect	182	102	183	103
rect	182	104	183	105
rect	182	105	183	106
rect	182	107	183	108
rect	182	108	183	109
rect	182	110	183	111
rect	182	111	183	112
rect	182	113	183	114
rect	182	114	183	115
rect	182	116	183	117
rect	182	117	183	118
rect	182	119	183	120
rect	182	120	183	121
rect	182	122	183	123
rect	182	123	183	124
rect	182	125	183	126
rect	182	126	183	127
rect	182	128	183	129
rect	182	129	183	130
rect	182	131	183	132
rect	182	132	183	133
rect	182	134	183	135
rect	182	135	183	136
rect	182	137	183	138
rect	182	138	183	139
rect	182	140	183	141
rect	182	141	183	142
rect	182	143	183	144
rect	182	144	183	145
rect	182	146	183	147
rect	182	147	183	148
rect	182	149	183	150
rect	182	150	183	151
rect	182	152	183	153
rect	182	153	183	154
rect	182	155	183	156
rect	182	156	183	157
rect	182	158	183	159
rect	182	159	183	160
rect	182	161	183	162
rect	182	162	183	163
rect	182	164	183	165
rect	182	165	183	166
rect	182	167	183	168
rect	182	168	183	169
rect	182	170	183	171
rect	182	171	183	172
rect	182	173	183	174
rect	182	174	183	175
rect	182	176	183	177
rect	182	177	183	178
rect	182	179	183	180
rect	182	180	183	181
rect	182	182	183	183
rect	182	183	183	184
rect	182	185	183	186
rect	182	186	183	187
rect	182	188	183	189
rect	182	189	183	190
rect	182	191	183	192
rect	182	192	183	193
rect	182	194	183	195
rect	182	195	183	196
rect	182	197	183	198
rect	182	198	183	199
rect	182	200	183	201
rect	182	201	183	202
rect	182	203	183	204
rect	182	204	183	205
rect	182	206	183	207
rect	182	207	183	208
rect	182	209	183	210
rect	182	210	183	211
rect	182	212	183	213
rect	182	213	183	214
rect	182	215	183	216
rect	182	216	183	217
rect	182	218	183	219
rect	182	219	183	220
rect	182	221	183	222
rect	182	222	183	223
rect	182	224	183	225
rect	182	225	183	226
rect	182	227	183	228
rect	182	228	183	229
rect	182	230	183	231
rect	182	231	183	232
rect	182	233	183	234
rect	182	234	183	235
rect	182	236	183	237
rect	182	237	183	238
rect	182	239	183	240
rect	182	240	183	241
rect	182	242	183	243
rect	182	243	183	244
rect	182	245	183	246
rect	182	246	183	247
rect	182	248	183	249
rect	182	249	183	250
rect	182	251	183	252
rect	182	252	183	253
rect	182	254	183	255
rect	182	255	183	256
rect	182	257	183	258
rect	182	258	183	259
rect	182	260	183	261
rect	182	261	183	262
rect	182	263	183	264
rect	182	264	183	265
rect	184	74	185	75
rect	184	75	185	76
rect	184	77	185	78
rect	184	78	185	79
rect	184	83	185	84
rect	184	84	185	85
rect	184	86	185	87
rect	184	87	185	88
rect	184	89	185	90
rect	184	90	185	91
rect	184	92	185	93
rect	184	93	185	94
rect	184	95	185	96
rect	184	96	185	97
rect	184	98	185	99
rect	184	99	185	100
rect	184	101	185	102
rect	184	102	185	103
rect	184	104	185	105
rect	184	105	185	106
rect	184	107	185	108
rect	184	108	185	109
rect	184	110	185	111
rect	184	111	185	112
rect	184	113	185	114
rect	184	114	185	115
rect	184	116	185	117
rect	184	117	185	118
rect	184	119	185	120
rect	184	120	185	121
rect	184	122	185	123
rect	184	123	185	124
rect	184	125	185	126
rect	184	126	185	127
rect	184	128	185	129
rect	184	129	185	130
rect	184	131	185	132
rect	184	132	185	133
rect	184	134	185	135
rect	184	135	185	136
rect	184	137	185	138
rect	184	138	185	139
rect	184	140	185	141
rect	184	141	185	142
rect	184	143	185	144
rect	184	144	185	145
rect	184	146	185	147
rect	184	147	185	148
rect	184	149	185	150
rect	184	150	185	151
rect	184	152	185	153
rect	184	153	185	154
rect	184	155	185	156
rect	184	156	185	157
rect	184	158	185	159
rect	184	159	185	160
rect	184	161	185	162
rect	184	162	185	163
rect	184	164	185	165
rect	184	165	185	166
rect	184	167	185	168
rect	184	168	185	169
rect	184	170	185	171
rect	184	171	185	172
rect	184	173	185	174
rect	184	174	185	175
rect	184	176	185	177
rect	184	177	185	178
rect	184	179	185	180
rect	184	180	185	181
rect	184	182	185	183
rect	184	183	185	184
rect	184	185	185	186
rect	184	186	185	187
rect	184	188	185	189
rect	184	189	185	190
rect	184	191	185	192
rect	184	192	185	193
rect	184	194	185	195
rect	184	195	185	196
rect	184	197	185	198
rect	184	198	185	199
rect	184	200	185	201
rect	184	201	185	202
rect	184	203	185	204
rect	184	204	185	205
rect	186	38	187	39
rect	186	39	187	40
rect	186	41	187	42
rect	186	42	187	43
rect	186	44	187	45
rect	186	45	187	46
rect	186	47	187	48
rect	186	48	187	49
rect	186	50	187	51
rect	186	51	187	52
rect	186	53	187	54
rect	186	54	187	55
rect	186	56	187	57
rect	186	57	187	58
rect	186	59	187	60
rect	186	60	187	61
rect	186	62	187	63
rect	186	63	187	64
rect	186	65	187	66
rect	186	66	187	67
rect	186	68	187	69
rect	186	69	187	70
rect	186	71	187	72
rect	186	72	187	73
rect	186	74	187	75
rect	186	75	187	76
rect	186	77	187	78
rect	186	78	187	79
rect	186	80	187	81
rect	186	81	187	82
rect	186	83	187	84
rect	186	84	187	85
rect	186	86	187	87
rect	186	87	187	88
rect	186	89	187	90
rect	186	90	187	91
rect	186	92	187	93
rect	186	93	187	94
rect	186	95	187	96
rect	186	96	187	97
rect	186	98	187	99
rect	186	99	187	100
rect	186	101	187	102
rect	186	102	187	103
rect	186	104	187	105
rect	186	105	187	106
rect	186	107	187	108
rect	186	108	187	109
rect	186	110	187	111
rect	186	111	187	112
rect	186	113	187	114
rect	186	114	187	115
rect	186	116	187	117
rect	186	117	187	118
rect	186	119	187	120
rect	186	120	187	121
rect	186	122	187	123
rect	186	123	187	124
rect	186	125	187	126
rect	186	126	187	127
rect	186	128	187	129
rect	186	129	187	130
rect	186	185	187	186
rect	186	186	187	187
rect	186	278	187	279
rect	186	279	187	280
rect	186	281	187	282
rect	186	282	187	283
rect	186	284	187	285
rect	186	285	187	286
rect	188	20	189	21
rect	188	21	189	22
rect	188	23	189	24
rect	188	24	189	25
rect	188	26	189	27
rect	188	27	189	28
rect	188	35	189	36
rect	188	36	189	37
rect	188	38	189	39
rect	188	39	189	40
rect	188	41	189	42
rect	188	42	189	43
rect	188	44	189	45
rect	188	45	189	46
rect	188	47	189	48
rect	188	48	189	49
rect	188	50	189	51
rect	188	51	189	52
rect	188	53	189	54
rect	188	54	189	55
rect	188	56	189	57
rect	188	57	189	58
rect	188	59	189	60
rect	188	60	189	61
rect	188	62	189	63
rect	188	63	189	64
rect	188	65	189	66
rect	188	66	189	67
rect	188	68	189	69
rect	188	69	189	70
rect	188	71	189	72
rect	188	72	189	73
rect	188	74	189	75
rect	188	75	189	76
rect	188	77	189	78
rect	188	78	189	79
rect	188	80	189	81
rect	188	81	189	82
rect	188	83	189	84
rect	188	84	189	85
rect	188	86	189	87
rect	188	87	189	88
rect	188	89	189	90
rect	188	90	189	91
rect	188	92	189	93
rect	188	93	189	94
rect	188	95	189	96
rect	188	96	189	97
rect	188	98	189	99
rect	188	99	189	100
rect	188	101	189	102
rect	188	102	189	103
rect	188	104	189	105
rect	188	105	189	106
rect	188	107	189	108
rect	188	108	189	109
rect	188	110	189	111
rect	188	111	189	112
rect	188	113	189	114
rect	188	114	189	115
rect	188	116	189	117
rect	188	117	189	118
rect	188	119	189	120
rect	188	120	189	121
rect	188	122	189	123
rect	188	123	189	124
rect	188	125	189	126
rect	188	126	189	127
rect	188	128	189	129
rect	188	129	189	130
rect	188	131	189	132
rect	188	132	189	133
rect	188	134	189	135
rect	188	135	189	136
rect	188	137	189	138
rect	188	138	189	139
rect	188	140	189	141
rect	188	141	189	142
rect	188	143	189	144
rect	188	144	189	145
rect	188	146	189	147
rect	188	147	189	148
rect	188	149	189	150
rect	188	150	189	151
rect	188	152	189	153
rect	188	153	189	154
rect	188	155	189	156
rect	188	156	189	157
rect	188	158	189	159
rect	188	159	189	160
rect	188	161	189	162
rect	188	162	189	163
rect	188	164	189	165
rect	188	165	189	166
rect	188	167	189	168
rect	188	168	189	169
rect	188	170	189	171
rect	188	171	189	172
rect	188	173	189	174
rect	188	174	189	175
rect	188	176	189	177
rect	188	177	189	178
rect	188	179	189	180
rect	188	180	189	181
rect	188	182	189	183
rect	188	183	189	184
rect	188	185	189	186
rect	188	186	189	187
rect	188	188	189	189
rect	188	189	189	190
rect	188	191	189	192
rect	188	192	189	193
rect	188	194	189	195
rect	188	195	189	196
rect	188	197	189	198
rect	188	198	189	199
rect	188	200	189	201
rect	188	201	189	202
rect	188	203	189	204
rect	188	204	189	205
rect	188	206	189	207
rect	188	207	189	208
rect	188	209	189	210
rect	188	210	189	211
rect	188	212	189	213
rect	188	213	189	214
rect	188	215	189	216
rect	188	216	189	217
rect	188	218	189	219
rect	188	219	189	220
rect	188	221	189	222
rect	188	222	189	223
rect	188	224	189	225
rect	188	225	189	226
rect	188	227	189	228
rect	188	228	189	229
rect	188	230	189	231
rect	188	231	189	232
rect	188	236	189	237
rect	188	237	189	238
rect	188	239	189	240
rect	188	240	189	241
rect	188	272	189	273
rect	188	273	189	274
rect	188	275	189	276
rect	188	276	189	277
rect	188	278	189	279
rect	188	279	189	280
rect	188	311	189	312
rect	188	312	189	313
rect	188	314	189	315
rect	188	315	189	316
rect	188	317	189	318
rect	188	318	189	319
rect	188	356	189	357
rect	188	357	189	358
rect	190	5	191	6
rect	190	6	191	7
rect	190	8	191	9
rect	190	9	191	10
rect	190	11	191	12
rect	190	12	191	13
rect	190	14	191	15
rect	190	15	191	16
rect	190	17	191	18
rect	190	18	191	19
rect	190	20	191	21
rect	190	21	191	22
rect	190	23	191	24
rect	190	24	191	25
rect	190	26	191	27
rect	190	27	191	28
rect	190	29	191	30
rect	190	30	191	31
rect	190	32	191	33
rect	190	33	191	34
rect	190	35	191	36
rect	190	36	191	37
rect	190	38	191	39
rect	190	39	191	40
rect	190	41	191	42
rect	190	42	191	43
rect	190	44	191	45
rect	190	45	191	46
rect	190	47	191	48
rect	190	48	191	49
rect	190	50	191	51
rect	190	51	191	52
rect	190	53	191	54
rect	190	54	191	55
rect	190	56	191	57
rect	190	57	191	58
rect	190	59	191	60
rect	190	60	191	61
rect	190	62	191	63
rect	190	63	191	64
rect	190	65	191	66
rect	190	66	191	67
rect	190	68	191	69
rect	190	69	191	70
rect	190	71	191	72
rect	190	72	191	73
rect	190	74	191	75
rect	190	75	191	76
rect	190	77	191	78
rect	190	78	191	79
rect	190	80	191	81
rect	190	81	191	82
rect	190	83	191	84
rect	190	84	191	85
rect	190	86	191	87
rect	190	87	191	88
rect	190	89	191	90
rect	190	90	191	91
rect	190	92	191	93
rect	190	93	191	94
rect	190	95	191	96
rect	190	96	191	97
rect	190	98	191	99
rect	190	99	191	100
rect	190	101	191	102
rect	190	102	191	103
rect	190	104	191	105
rect	190	105	191	106
rect	190	107	191	108
rect	190	108	191	109
rect	190	110	191	111
rect	190	111	191	112
rect	190	113	191	114
rect	190	114	191	115
rect	190	116	191	117
rect	190	117	191	118
rect	190	119	191	120
rect	190	120	191	121
rect	190	122	191	123
rect	190	123	191	124
rect	190	125	191	126
rect	190	126	191	127
rect	190	128	191	129
rect	190	129	191	130
rect	190	131	191	132
rect	190	132	191	133
rect	190	134	191	135
rect	190	135	191	136
rect	190	137	191	138
rect	190	138	191	139
rect	190	140	191	141
rect	190	141	191	142
rect	190	143	191	144
rect	190	144	191	145
rect	190	146	191	147
rect	190	147	191	148
rect	190	149	191	150
rect	190	150	191	151
rect	190	152	191	153
rect	190	153	191	154
rect	190	155	191	156
rect	190	156	191	157
rect	190	158	191	159
rect	190	159	191	160
rect	190	161	191	162
rect	190	162	191	163
rect	190	164	191	165
rect	190	165	191	166
rect	190	167	191	168
rect	190	168	191	169
rect	190	170	191	171
rect	190	171	191	172
rect	190	173	191	174
rect	190	174	191	175
rect	190	176	191	177
rect	190	177	191	178
rect	190	179	191	180
rect	190	180	191	181
rect	190	182	191	183
rect	190	183	191	184
rect	190	185	191	186
rect	190	186	191	187
rect	190	188	191	189
rect	190	189	191	190
rect	190	191	191	192
rect	190	192	191	193
rect	190	194	191	195
rect	190	195	191	196
rect	190	197	191	198
rect	190	198	191	199
rect	190	200	191	201
rect	190	201	191	202
rect	190	203	191	204
rect	190	204	191	205
rect	190	206	191	207
rect	190	207	191	208
rect	190	209	191	210
rect	190	210	191	211
rect	190	212	191	213
rect	190	213	191	214
rect	190	215	191	216
rect	190	216	191	217
rect	190	218	191	219
rect	190	219	191	220
rect	190	221	191	222
rect	190	222	191	223
rect	190	224	191	225
rect	190	225	191	226
rect	190	227	191	228
rect	190	228	191	229
rect	190	230	191	231
rect	190	231	191	232
rect	190	233	191	234
rect	190	234	191	235
rect	190	236	191	237
rect	190	237	191	238
rect	190	239	191	240
rect	190	240	191	241
rect	190	242	191	243
rect	190	243	191	244
rect	190	245	191	246
rect	190	246	191	247
rect	190	248	191	249
rect	190	249	191	250
rect	190	251	191	252
rect	190	252	191	253
rect	190	254	191	255
rect	190	255	191	256
rect	190	257	191	258
rect	190	258	191	259
rect	190	260	191	261
rect	190	261	191	262
rect	190	263	191	264
rect	190	264	191	265
rect	190	266	191	267
rect	190	267	191	268
rect	190	269	191	270
rect	190	270	191	271
rect	190	272	191	273
rect	190	273	191	274
rect	190	275	191	276
rect	190	276	191	277
rect	190	278	191	279
rect	190	279	191	280
rect	190	281	191	282
rect	190	282	191	283
rect	190	284	191	285
rect	190	285	191	286
rect	190	287	191	288
rect	190	288	191	289
rect	190	290	191	291
rect	190	291	191	292
rect	190	293	191	294
rect	190	294	191	295
rect	190	296	191	297
rect	190	297	191	298
rect	190	299	191	300
rect	190	300	191	301
rect	190	302	191	303
rect	190	303	191	304
rect	190	304	191	305
rect	190	305	191	306
rect	190	306	191	307
rect	190	308	191	309
rect	190	309	191	310
rect	190	311	191	312
rect	190	312	191	313
rect	190	314	191	315
rect	190	315	191	316
rect	190	317	191	318
rect	190	318	191	319
rect	190	319	191	320
rect	190	320	191	321
rect	190	321	191	322
rect	190	323	191	324
rect	190	324	191	325
rect	190	326	191	327
rect	190	327	191	328
rect	190	328	191	329
rect	190	329	191	330
rect	190	330	191	331
rect	190	332	191	333
rect	190	333	191	334
rect	190	335	191	336
rect	190	336	191	337
rect	190	337	191	338
rect	190	338	191	339
rect	190	339	191	340
rect	190	340	191	341
rect	190	341	191	342
rect	190	342	191	343
rect	190	343	191	344
rect	190	344	191	345
rect	190	345	191	346
rect	190	347	191	348
rect	190	348	191	349
rect	190	350	191	351
rect	190	351	191	352
rect	190	352	191	353
rect	190	353	191	354
rect	190	354	191	355
rect	190	356	191	357
rect	190	357	191	358
rect	190	359	191	360
rect	190	360	191	361
rect	190	361	191	362
rect	190	362	191	363
rect	190	363	191	364
rect	190	365	191	366
rect	190	366	191	367
rect	199	296	200	297
rect	199	297	200	298
rect	199	299	200	300
rect	199	300	200	301
rect	199	302	200	303
rect	199	303	200	304
rect	201	254	202	255
rect	201	255	202	256
rect	201	257	202	258
rect	201	258	202	259
rect	201	260	202	261
rect	201	261	202	262
rect	201	262	202	263
rect	201	263	202	264
rect	201	264	202	265
rect	201	266	202	267
rect	201	267	202	268
rect	201	269	202	270
rect	201	270	202	271
rect	201	272	202	273
rect	201	273	202	274
rect	201	275	202	276
rect	201	276	202	277
rect	201	278	202	279
rect	201	279	202	280
rect	201	281	202	282
rect	201	282	202	283
rect	201	284	202	285
rect	201	285	202	286
rect	201	287	202	288
rect	201	288	202	289
rect	201	290	202	291
rect	201	291	202	292
rect	201	293	202	294
rect	201	294	202	295
rect	201	296	202	297
rect	201	297	202	298
rect	201	299	202	300
rect	201	300	202	301
rect	201	302	202	303
rect	201	303	202	304
rect	201	305	202	306
rect	201	306	202	307
rect	201	308	202	309
rect	201	309	202	310
rect	201	311	202	312
rect	201	312	202	313
rect	201	314	202	315
rect	201	315	202	316
rect	201	317	202	318
rect	201	318	202	319
rect	201	319	202	320
rect	201	320	202	321
rect	201	321	202	322
rect	201	322	202	323
rect	201	323	202	324
rect	201	324	202	325
rect	201	325	202	326
rect	201	326	202	327
rect	201	327	202	328
rect	201	328	202	329
rect	201	329	202	330
rect	201	330	202	331
rect	201	332	202	333
rect	201	333	202	334
rect	201	335	202	336
rect	201	336	202	337
rect	201	337	202	338
rect	201	338	202	339
rect	201	339	202	340
rect	201	340	202	341
rect	201	341	202	342
rect	201	342	202	343
rect	203	101	204	102
rect	203	102	204	103
rect	203	104	204	105
rect	203	105	204	106
rect	203	107	204	108
rect	203	108	204	109
rect	203	110	204	111
rect	203	111	204	112
rect	203	116	204	117
rect	203	117	204	118
rect	203	119	204	120
rect	203	120	204	121
rect	203	152	204	153
rect	203	153	204	154
rect	203	191	204	192
rect	203	192	204	193
rect	203	194	204	195
rect	203	195	204	196
rect	203	197	204	198
rect	203	198	204	199
rect	203	200	204	201
rect	203	201	204	202
rect	203	203	204	204
rect	203	204	204	205
rect	203	206	204	207
rect	203	207	204	208
rect	203	209	204	210
rect	203	210	204	211
rect	203	224	204	225
rect	203	225	204	226
rect	203	227	204	228
rect	203	228	204	229
rect	203	230	204	231
rect	203	231	204	232
rect	203	233	204	234
rect	203	234	204	235
rect	203	236	204	237
rect	203	237	204	238
rect	203	239	204	240
rect	203	240	204	241
rect	203	242	204	243
rect	203	243	204	244
rect	203	245	204	246
rect	203	246	204	247
rect	203	248	204	249
rect	203	249	204	250
rect	203	251	204	252
rect	203	252	204	253
rect	203	254	204	255
rect	203	255	204	256
rect	203	257	204	258
rect	203	258	204	259
rect	203	260	204	261
rect	203	261	204	262
rect	203	262	204	263
rect	203	263	204	264
rect	203	264	204	265
rect	203	266	204	267
rect	203	267	204	268
rect	203	269	204	270
rect	203	270	204	271
rect	203	272	204	273
rect	203	273	204	274
rect	203	275	204	276
rect	203	276	204	277
rect	203	278	204	279
rect	203	279	204	280
rect	203	281	204	282
rect	203	282	204	283
rect	203	284	204	285
rect	203	285	204	286
rect	203	287	204	288
rect	203	288	204	289
rect	203	290	204	291
rect	203	291	204	292
rect	203	293	204	294
rect	203	294	204	295
rect	203	296	204	297
rect	203	297	204	298
rect	203	299	204	300
rect	203	300	204	301
rect	203	302	204	303
rect	203	303	204	304
rect	203	305	204	306
rect	203	306	204	307
rect	203	308	204	309
rect	203	309	204	310
rect	203	311	204	312
rect	203	312	204	313
rect	203	314	204	315
rect	203	315	204	316
rect	203	317	204	318
rect	203	318	204	319
rect	203	319	204	320
rect	203	320	204	321
rect	203	321	204	322
rect	203	322	204	323
rect	203	323	204	324
rect	203	324	204	325
rect	203	325	204	326
rect	203	326	204	327
rect	203	327	204	328
rect	203	328	204	329
rect	203	329	204	330
rect	203	330	204	331
rect	203	332	204	333
rect	203	333	204	334
rect	203	335	204	336
rect	203	336	204	337
rect	203	337	204	338
rect	203	338	204	339
rect	203	339	204	340
rect	203	340	204	341
rect	203	341	204	342
rect	203	342	204	343
rect	203	344	204	345
rect	203	345	204	346
rect	205	38	206	39
rect	205	39	206	40
rect	205	41	206	42
rect	205	42	206	43
rect	205	44	206	45
rect	205	45	206	46
rect	205	47	206	48
rect	205	48	206	49
rect	205	50	206	51
rect	205	51	206	52
rect	205	53	206	54
rect	205	54	206	55
rect	205	56	206	57
rect	205	57	206	58
rect	205	59	206	60
rect	205	60	206	61
rect	205	62	206	63
rect	205	63	206	64
rect	205	65	206	66
rect	205	66	206	67
rect	205	68	206	69
rect	205	69	206	70
rect	205	71	206	72
rect	205	72	206	73
rect	205	74	206	75
rect	205	75	206	76
rect	205	77	206	78
rect	205	78	206	79
rect	205	80	206	81
rect	205	81	206	82
rect	205	83	206	84
rect	205	84	206	85
rect	205	86	206	87
rect	205	87	206	88
rect	205	89	206	90
rect	205	90	206	91
rect	205	92	206	93
rect	205	93	206	94
rect	205	95	206	96
rect	205	96	206	97
rect	205	98	206	99
rect	205	99	206	100
rect	205	101	206	102
rect	205	102	206	103
rect	205	104	206	105
rect	205	105	206	106
rect	205	107	206	108
rect	205	108	206	109
rect	205	110	206	111
rect	205	111	206	112
rect	205	113	206	114
rect	205	114	206	115
rect	205	116	206	117
rect	205	117	206	118
rect	205	119	206	120
rect	205	120	206	121
rect	205	122	206	123
rect	205	123	206	124
rect	205	125	206	126
rect	205	126	206	127
rect	205	128	206	129
rect	205	129	206	130
rect	205	131	206	132
rect	205	132	206	133
rect	205	134	206	135
rect	205	135	206	136
rect	205	137	206	138
rect	205	138	206	139
rect	205	140	206	141
rect	205	141	206	142
rect	205	143	206	144
rect	205	144	206	145
rect	205	146	206	147
rect	205	147	206	148
rect	205	149	206	150
rect	205	150	206	151
rect	205	152	206	153
rect	205	153	206	154
rect	205	155	206	156
rect	205	156	206	157
rect	205	158	206	159
rect	205	159	206	160
rect	205	161	206	162
rect	205	162	206	163
rect	205	164	206	165
rect	205	165	206	166
rect	205	167	206	168
rect	205	168	206	169
rect	205	170	206	171
rect	205	171	206	172
rect	205	173	206	174
rect	205	174	206	175
rect	205	176	206	177
rect	205	177	206	178
rect	205	179	206	180
rect	205	180	206	181
rect	205	182	206	183
rect	205	183	206	184
rect	205	185	206	186
rect	205	186	206	187
rect	205	188	206	189
rect	205	189	206	190
rect	205	191	206	192
rect	205	192	206	193
rect	205	194	206	195
rect	205	195	206	196
rect	205	197	206	198
rect	205	198	206	199
rect	205	200	206	201
rect	205	201	206	202
rect	205	203	206	204
rect	205	204	206	205
rect	205	206	206	207
rect	205	207	206	208
rect	205	209	206	210
rect	205	210	206	211
rect	205	212	206	213
rect	205	213	206	214
rect	205	215	206	216
rect	205	216	206	217
rect	205	218	206	219
rect	205	219	206	220
rect	205	221	206	222
rect	205	222	206	223
rect	205	224	206	225
rect	205	225	206	226
rect	205	227	206	228
rect	205	228	206	229
rect	205	230	206	231
rect	205	231	206	232
rect	205	233	206	234
rect	205	234	206	235
rect	205	236	206	237
rect	205	237	206	238
rect	205	239	206	240
rect	205	240	206	241
rect	205	242	206	243
rect	205	243	206	244
rect	205	245	206	246
rect	205	246	206	247
rect	205	248	206	249
rect	205	249	206	250
rect	205	251	206	252
rect	205	252	206	253
rect	205	254	206	255
rect	205	255	206	256
rect	205	257	206	258
rect	205	258	206	259
rect	205	260	206	261
rect	205	261	206	262
rect	205	262	206	263
rect	205	263	206	264
rect	205	264	206	265
rect	205	266	206	267
rect	205	267	206	268
rect	205	269	206	270
rect	205	270	206	271
rect	205	272	206	273
rect	205	273	206	274
rect	205	275	206	276
rect	205	276	206	277
rect	205	278	206	279
rect	205	279	206	280
rect	205	281	206	282
rect	205	282	206	283
rect	205	284	206	285
rect	205	285	206	286
rect	205	287	206	288
rect	205	288	206	289
rect	205	289	206	290
rect	205	290	206	291
rect	205	291	206	292
rect	205	293	206	294
rect	205	294	206	295
rect	205	296	206	297
rect	205	297	206	298
rect	205	299	206	300
rect	205	300	206	301
rect	205	302	206	303
rect	205	303	206	304
rect	205	304	206	305
rect	205	305	206	306
rect	205	306	206	307
rect	207	5	208	6
rect	207	6	208	7
rect	207	17	208	18
rect	207	18	208	19
rect	207	20	208	21
rect	207	21	208	22
rect	207	23	208	24
rect	207	24	208	25
rect	207	26	208	27
rect	207	27	208	28
rect	207	29	208	30
rect	207	30	208	31
rect	207	32	208	33
rect	207	33	208	34
rect	207	35	208	36
rect	207	36	208	37
rect	207	38	208	39
rect	207	39	208	40
rect	207	41	208	42
rect	207	42	208	43
rect	207	44	208	45
rect	207	45	208	46
rect	207	47	208	48
rect	207	48	208	49
rect	207	50	208	51
rect	207	51	208	52
rect	207	53	208	54
rect	207	54	208	55
rect	207	56	208	57
rect	207	57	208	58
rect	207	59	208	60
rect	207	60	208	61
rect	207	62	208	63
rect	207	63	208	64
rect	207	65	208	66
rect	207	66	208	67
rect	207	68	208	69
rect	207	69	208	70
rect	207	71	208	72
rect	207	72	208	73
rect	207	74	208	75
rect	207	75	208	76
rect	207	77	208	78
rect	207	78	208	79
rect	207	80	208	81
rect	207	81	208	82
rect	207	83	208	84
rect	207	84	208	85
rect	207	86	208	87
rect	207	87	208	88
rect	207	89	208	90
rect	207	90	208	91
rect	207	92	208	93
rect	207	93	208	94
rect	207	95	208	96
rect	207	96	208	97
rect	207	98	208	99
rect	207	99	208	100
rect	207	101	208	102
rect	207	102	208	103
rect	207	104	208	105
rect	207	105	208	106
rect	207	107	208	108
rect	207	108	208	109
rect	207	110	208	111
rect	207	111	208	112
rect	207	113	208	114
rect	207	114	208	115
rect	207	116	208	117
rect	207	117	208	118
rect	207	119	208	120
rect	207	120	208	121
rect	207	122	208	123
rect	207	123	208	124
rect	207	125	208	126
rect	207	126	208	127
rect	207	128	208	129
rect	207	129	208	130
rect	207	131	208	132
rect	207	132	208	133
rect	207	134	208	135
rect	207	135	208	136
rect	207	137	208	138
rect	207	138	208	139
rect	207	140	208	141
rect	207	141	208	142
rect	207	143	208	144
rect	207	144	208	145
rect	207	146	208	147
rect	207	147	208	148
rect	207	149	208	150
rect	207	150	208	151
rect	207	152	208	153
rect	207	153	208	154
rect	207	155	208	156
rect	207	156	208	157
rect	207	158	208	159
rect	207	159	208	160
rect	207	161	208	162
rect	207	162	208	163
rect	207	164	208	165
rect	207	165	208	166
rect	207	167	208	168
rect	207	168	208	169
rect	207	170	208	171
rect	207	171	208	172
rect	207	173	208	174
rect	207	174	208	175
rect	207	176	208	177
rect	207	177	208	178
rect	207	179	208	180
rect	207	180	208	181
rect	207	182	208	183
rect	207	183	208	184
rect	207	185	208	186
rect	207	186	208	187
rect	207	188	208	189
rect	207	189	208	190
rect	207	191	208	192
rect	207	192	208	193
rect	207	194	208	195
rect	207	195	208	196
rect	207	197	208	198
rect	207	198	208	199
rect	207	200	208	201
rect	207	201	208	202
rect	207	203	208	204
rect	207	204	208	205
rect	207	206	208	207
rect	207	207	208	208
rect	207	209	208	210
rect	207	210	208	211
rect	207	212	208	213
rect	207	213	208	214
rect	207	215	208	216
rect	207	216	208	217
rect	207	218	208	219
rect	207	219	208	220
rect	207	221	208	222
rect	207	222	208	223
rect	207	224	208	225
rect	207	225	208	226
rect	207	227	208	228
rect	207	228	208	229
rect	207	230	208	231
rect	207	231	208	232
rect	207	233	208	234
rect	207	234	208	235
rect	207	236	208	237
rect	207	237	208	238
rect	207	239	208	240
rect	207	240	208	241
rect	207	242	208	243
rect	207	243	208	244
rect	207	245	208	246
rect	207	246	208	247
rect	207	248	208	249
rect	207	249	208	250
rect	207	251	208	252
rect	207	252	208	253
rect	207	254	208	255
rect	207	255	208	256
rect	207	257	208	258
rect	207	258	208	259
rect	207	260	208	261
rect	207	261	208	262
rect	207	262	208	263
rect	207	263	208	264
rect	207	264	208	265
rect	207	266	208	267
rect	207	267	208	268
rect	207	269	208	270
rect	207	270	208	271
rect	207	272	208	273
rect	207	273	208	274
rect	207	275	208	276
rect	207	276	208	277
rect	207	278	208	279
rect	207	279	208	280
rect	207	281	208	282
rect	207	282	208	283
rect	207	284	208	285
rect	207	285	208	286
rect	207	287	208	288
rect	207	288	208	289
rect	207	289	208	290
rect	207	290	208	291
rect	207	291	208	292
rect	207	293	208	294
rect	207	294	208	295
rect	207	296	208	297
rect	207	297	208	298
rect	207	299	208	300
rect	207	300	208	301
rect	207	302	208	303
rect	207	303	208	304
rect	207	304	208	305
rect	207	305	208	306
rect	207	306	208	307
rect	207	308	208	309
rect	207	309	208	310
rect	207	311	208	312
rect	207	312	208	313
rect	216	5	217	6
rect	216	6	217	7
rect	216	8	217	9
rect	216	9	217	10
rect	216	11	217	12
rect	216	12	217	13
rect	216	14	217	15
rect	216	15	217	16
rect	216	17	217	18
rect	216	18	217	19
rect	216	20	217	21
rect	216	21	217	22
rect	216	23	217	24
rect	216	24	217	25
rect	216	26	217	27
rect	216	27	217	28
rect	216	29	217	30
rect	216	30	217	31
rect	216	32	217	33
rect	216	33	217	34
rect	216	35	217	36
rect	216	36	217	37
rect	216	38	217	39
rect	216	39	217	40
rect	216	41	217	42
rect	216	42	217	43
rect	216	44	217	45
rect	216	45	217	46
rect	216	47	217	48
rect	216	48	217	49
rect	216	50	217	51
rect	216	51	217	52
rect	216	53	217	54
rect	216	54	217	55
rect	216	56	217	57
rect	216	57	217	58
rect	216	59	217	60
rect	216	60	217	61
rect	216	62	217	63
rect	216	63	217	64
rect	216	65	217	66
rect	216	66	217	67
rect	216	68	217	69
rect	216	69	217	70
rect	216	71	217	72
rect	216	72	217	73
rect	216	74	217	75
rect	216	75	217	76
rect	216	77	217	78
rect	216	78	217	79
rect	216	80	217	81
rect	216	81	217	82
rect	216	83	217	84
rect	216	84	217	85
rect	216	86	217	87
rect	216	87	217	88
rect	216	89	217	90
rect	216	90	217	91
rect	216	92	217	93
rect	216	93	217	94
rect	216	95	217	96
rect	216	96	217	97
rect	216	98	217	99
rect	216	99	217	100
rect	216	101	217	102
rect	216	102	217	103
rect	216	104	217	105
rect	216	105	217	106
rect	216	107	217	108
rect	216	108	217	109
rect	216	110	217	111
rect	216	111	217	112
rect	216	113	217	114
rect	216	114	217	115
rect	216	116	217	117
rect	216	117	217	118
rect	216	119	217	120
rect	216	120	217	121
rect	216	122	217	123
rect	216	123	217	124
rect	216	125	217	126
rect	216	126	217	127
rect	216	128	217	129
rect	216	129	217	130
rect	216	131	217	132
rect	216	132	217	133
rect	216	134	217	135
rect	216	135	217	136
rect	216	137	217	138
rect	216	138	217	139
rect	216	140	217	141
rect	216	141	217	142
rect	216	143	217	144
rect	216	144	217	145
rect	216	146	217	147
rect	216	147	217	148
rect	216	149	217	150
rect	216	150	217	151
rect	216	152	217	153
rect	216	153	217	154
rect	216	155	217	156
rect	216	156	217	157
rect	216	158	217	159
rect	216	159	217	160
rect	216	161	217	162
rect	216	162	217	163
rect	216	164	217	165
rect	216	165	217	166
rect	216	167	217	168
rect	216	168	217	169
rect	216	170	217	171
rect	216	171	217	172
rect	216	173	217	174
rect	216	174	217	175
rect	216	176	217	177
rect	216	177	217	178
rect	216	179	217	180
rect	216	180	217	181
rect	216	182	217	183
rect	216	183	217	184
rect	216	185	217	186
rect	216	186	217	187
rect	216	188	217	189
rect	216	189	217	190
rect	216	191	217	192
rect	216	192	217	193
rect	216	194	217	195
rect	216	195	217	196
rect	216	197	217	198
rect	216	198	217	199
rect	216	200	217	201
rect	216	201	217	202
rect	216	203	217	204
rect	216	204	217	205
rect	216	206	217	207
rect	216	207	217	208
rect	218	2	219	3
rect	218	3	219	4
rect	218	5	219	6
rect	218	6	219	7
rect	218	14	219	15
rect	218	15	219	16
rect	218	17	219	18
rect	218	18	219	19
rect	218	74	219	75
rect	218	75	219	76
rect	218	77	219	78
rect	218	78	219	79
rect	218	80	219	81
rect	218	81	219	82
rect	218	83	219	84
rect	218	84	219	85
rect	218	86	219	87
rect	218	87	219	88
rect	218	89	219	90
rect	218	90	219	91
rect	218	92	219	93
rect	218	93	219	94
rect	218	95	219	96
rect	218	96	219	97
rect	218	98	219	99
rect	218	99	219	100
rect	218	101	219	102
rect	218	102	219	103
rect	218	104	219	105
rect	218	105	219	106
rect	218	131	219	132
rect	218	132	219	133
rect	218	134	219	135
rect	218	135	219	136
rect	218	137	219	138
rect	218	138	219	139
rect	218	146	219	147
rect	218	147	219	148
rect	218	149	219	150
rect	218	150	219	151
rect	218	176	219	177
rect	218	177	219	178
rect	218	179	219	180
rect	218	180	219	181
rect	218	239	219	240
rect	218	240	219	241
rect	218	242	219	243
rect	218	243	219	244
rect	218	245	219	246
rect	218	246	219	247
rect	218	257	219	258
rect	218	258	219	259
rect	218	260	219	261
rect	218	261	219	262
rect	218	262	219	263
rect	218	263	219	264
rect	218	264	219	265
rect	218	278	219	279
rect	218	279	219	280
rect	218	280	219	281
rect	218	281	219	282
rect	218	282	219	283
rect	227	200	228	201
rect	227	201	228	202
rect	227	203	228	204
rect	227	204	228	205
rect	227	206	228	207
rect	227	207	228	208
rect	229	203	230	204
rect	229	204	230	205
rect	229	206	230	207
rect	229	207	230	208
rect	231	140	232	141
rect	231	141	232	142
rect	231	143	232	144
rect	231	144	232	145
rect	231	146	232	147
rect	231	147	232	148
rect	231	149	232	150
rect	231	150	232	151
rect	231	152	232	153
rect	231	153	232	154
rect	231	155	232	156
rect	231	156	232	157
rect	231	158	232	159
rect	231	159	232	160
rect	231	161	232	162
rect	231	162	232	163
rect	231	164	232	165
rect	231	165	232	166
rect	231	167	232	168
rect	231	168	232	169
rect	231	170	232	171
rect	231	171	232	172
rect	231	173	232	174
rect	231	174	232	175
rect	231	176	232	177
rect	231	177	232	178
rect	231	179	232	180
rect	231	180	232	181
rect	231	182	232	183
rect	231	183	232	184
rect	231	185	232	186
rect	231	186	232	187
rect	231	188	232	189
rect	231	189	232	190
rect	231	191	232	192
rect	231	192	232	193
rect	231	194	232	195
rect	231	195	232	196
rect	231	197	232	198
rect	231	198	232	199
rect	231	200	232	201
rect	231	201	232	202
rect	231	203	232	204
rect	231	204	232	205
rect	231	206	232	207
rect	231	207	232	208
rect	231	209	232	210
rect	231	210	232	211
rect	231	212	232	213
rect	231	213	232	214
rect	231	215	232	216
rect	231	216	232	217
rect	231	218	232	219
rect	231	219	232	220
rect	231	221	232	222
rect	231	222	232	223
rect	231	224	232	225
rect	231	225	232	226
rect	231	227	232	228
rect	231	228	232	229
rect	231	230	232	231
rect	231	231	232	232
rect	231	233	232	234
rect	231	234	232	235
rect	231	236	232	237
rect	231	237	232	238
rect	231	239	232	240
rect	231	240	232	241
rect	231	242	232	243
rect	231	243	232	244
rect	231	245	232	246
rect	231	246	232	247
rect	231	248	232	249
rect	231	249	232	250
rect	231	251	232	252
rect	231	252	232	253
rect	233	8	234	9
rect	233	9	234	10
rect	233	11	234	12
rect	233	12	234	13
rect	233	26	234	27
rect	233	27	234	28
rect	233	32	234	33
rect	233	33	234	34
rect	233	35	234	36
rect	233	36	234	37
rect	233	38	234	39
rect	233	39	234	40
rect	233	41	234	42
rect	233	42	234	43
rect	233	44	234	45
rect	233	45	234	46
rect	233	47	234	48
rect	233	48	234	49
rect	233	50	234	51
rect	233	51	234	52
rect	233	53	234	54
rect	233	54	234	55
rect	233	71	234	72
rect	233	72	234	73
rect	233	74	234	75
rect	233	75	234	76
rect	233	77	234	78
rect	233	78	234	79
rect	233	80	234	81
rect	233	81	234	82
rect	233	83	234	84
rect	233	84	234	85
rect	233	86	234	87
rect	233	87	234	88
rect	233	89	234	90
rect	233	90	234	91
rect	233	92	234	93
rect	233	93	234	94
rect	233	95	234	96
rect	233	96	234	97
rect	233	98	234	99
rect	233	99	234	100
rect	233	101	234	102
rect	233	102	234	103
rect	233	104	234	105
rect	233	105	234	106
rect	233	107	234	108
rect	233	108	234	109
rect	233	110	234	111
rect	233	111	234	112
rect	233	113	234	114
rect	233	114	234	115
rect	233	116	234	117
rect	233	117	234	118
rect	233	119	234	120
rect	233	120	234	121
rect	233	122	234	123
rect	233	123	234	124
rect	233	125	234	126
rect	233	126	234	127
rect	233	128	234	129
rect	233	129	234	130
rect	233	130	234	131
rect	233	131	234	132
rect	233	132	234	133
rect	233	134	234	135
rect	233	135	234	136
rect	233	137	234	138
rect	233	138	234	139
rect	233	140	234	141
rect	233	141	234	142
rect	233	143	234	144
rect	233	144	234	145
rect	233	146	234	147
rect	233	147	234	148
rect	233	149	234	150
rect	233	150	234	151
rect	233	152	234	153
rect	233	153	234	154
rect	233	155	234	156
rect	233	156	234	157
rect	233	158	234	159
rect	233	159	234	160
rect	233	161	234	162
rect	233	162	234	163
rect	233	164	234	165
rect	233	165	234	166
rect	233	167	234	168
rect	233	168	234	169
rect	233	170	234	171
rect	233	171	234	172
rect	233	173	234	174
rect	233	174	234	175
rect	233	176	234	177
rect	233	177	234	178
rect	233	179	234	180
rect	233	180	234	181
rect	233	182	234	183
rect	233	183	234	184
rect	233	185	234	186
rect	233	186	234	187
rect	233	188	234	189
rect	233	189	234	190
rect	233	191	234	192
rect	233	192	234	193
rect	233	194	234	195
rect	233	195	234	196
rect	233	197	234	198
rect	233	198	234	199
rect	233	200	234	201
rect	233	201	234	202
rect	233	203	234	204
rect	233	204	234	205
rect	233	206	234	207
rect	233	207	234	208
rect	233	209	234	210
rect	233	210	234	211
rect	233	212	234	213
rect	233	213	234	214
rect	233	215	234	216
rect	233	216	234	217
rect	233	218	234	219
rect	233	219	234	220
rect	233	221	234	222
rect	233	222	234	223
rect	233	224	234	225
rect	233	225	234	226
rect	233	227	234	228
rect	233	228	234	229
rect	233	230	234	231
rect	233	231	234	232
rect	233	233	234	234
rect	233	234	234	235
rect	233	236	234	237
rect	233	237	234	238
rect	233	239	234	240
rect	233	240	234	241
rect	242	155	243	156
rect	242	156	243	157
rect	242	158	243	159
rect	242	159	243	160
rect	242	161	243	162
rect	242	162	243	163
rect	242	164	243	165
rect	242	165	243	166
rect	242	167	243	168
rect	242	168	243	169
rect	242	170	243	171
rect	242	171	243	172
rect	242	197	243	198
rect	242	198	243	199
rect	242	200	243	201
rect	242	201	243	202
rect	242	203	243	204
rect	242	204	243	205
rect	242	206	243	207
rect	242	207	243	208
rect	242	209	243	210
rect	242	210	243	211
rect	242	212	243	213
rect	242	213	243	214
rect	242	215	243	216
rect	242	216	243	217
rect	242	218	243	219
rect	242	219	243	220
rect	242	221	243	222
rect	242	222	243	223
rect	242	224	243	225
rect	242	225	243	226
rect	242	227	243	228
rect	242	228	243	229
rect	242	230	243	231
rect	242	231	243	232
rect	242	233	243	234
rect	242	234	243	235
rect	242	236	243	237
rect	242	237	243	238
rect	242	239	243	240
rect	242	240	243	241
rect	242	241	243	242
rect	242	242	243	243
rect	242	243	243	244
rect	244	23	245	24
rect	244	24	245	25
rect	244	32	245	33
rect	244	33	245	34
rect	244	35	245	36
rect	244	36	245	37
rect	244	119	245	120
rect	244	120	245	121
rect	244	152	245	153
rect	244	153	245	154
rect	244	155	245	156
rect	244	156	245	157
rect	244	158	245	159
rect	244	159	245	160
rect	244	161	245	162
rect	244	162	245	163
rect	244	164	245	165
rect	244	165	245	166
rect	244	167	245	168
rect	244	168	245	169
rect	244	197	245	198
rect	244	198	245	199
rect	244	200	245	201
rect	244	201	245	202
rect	244	203	245	204
rect	244	204	245	205
rect	244	206	245	207
rect	244	207	245	208
rect	244	209	245	210
rect	244	210	245	211
rect	244	242	245	243
rect	244	243	245	244
rect	244	245	245	246
rect	244	246	245	247
rect	244	248	245	249
rect	244	249	245	250
rect	253	8	254	9
rect	253	9	254	10
rect	253	11	254	12
rect	253	12	254	13
rect	253	23	254	24
rect	253	24	254	25
rect	253	26	254	27
rect	253	27	254	28
rect	253	62	254	63
rect	253	63	254	64
rect	253	152	254	153
rect	253	153	254	154
rect	253	215	254	216
rect	253	216	254	217
rect	253	218	254	219
rect	253	219	254	220
rect	253	221	254	222
rect	253	222	254	223
rect	253	236	254	237
rect	253	237	254	238
rect	253	251	254	252
rect	253	252	254	253
rect	253	253	254	254
rect	253	254	254	255
rect	253	255	254	256
rect	262	35	263	36
rect	262	36	263	37
rect	262	38	263	39
rect	262	39	263	40
rect	262	98	263	99
rect	262	99	263	100
rect	262	101	263	102
rect	262	102	263	103
rect	262	104	263	105
rect	262	105	263	106
rect	262	137	263	138
rect	262	138	263	139
rect	262	140	263	141
rect	262	141	263	142
rect	262	200	263	201
rect	262	201	263	202
rect	262	203	263	204
rect	262	204	263	205
rect	262	221	263	222
rect	262	222	263	223
rect	262	224	263	225
rect	262	225	263	226
rect	271	188	272	189
rect	271	189	272	190
rect	271	190	272	191
rect	271	191	272	192
rect	271	192	272	193
rect	273	8	274	9
rect	273	9	274	10
rect	273	11	274	12
rect	273	12	274	13
rect	273	47	274	48
rect	273	48	274	49
rect	273	50	274	51
rect	273	51	274	52
rect	273	176	274	177
rect	273	177	274	178
rect	273	179	274	180
rect	273	180	274	181
rect	273	182	274	183
rect	273	183	274	184
rect	273	185	274	186
rect	273	186	274	187
rect	273	188	274	189
rect	273	189	274	190
rect	273	212	274	213
rect	273	213	274	214
rect	273	214	274	215
rect	273	215	274	216
rect	273	216	274	217
rect	282	164	283	165
rect	282	165	283	166
rect	282	167	283	168
rect	282	168	283	169
rect	282	170	283	171
rect	282	171	283	172
rect	282	173	283	174
rect	282	174	283	175
rect	282	176	283	177
rect	282	177	283	178
rect	284	86	285	87
rect	284	87	285	88
rect	284	110	285	111
rect	284	111	285	112
rect	284	112	285	113
rect	284	113	285	114
rect	284	114	285	115
rect	284	158	285	159
rect	284	159	285	160
rect	284	161	285	162
rect	284	162	285	163
rect	284	164	285	165
rect	284	165	285	166
rect	284	167	285	168
rect	284	168	285	169
rect	284	170	285	171
rect	284	171	285	172
rect	284	173	285	174
rect	284	174	285	175
rect	284	176	285	177
rect	284	177	285	178
rect	284	179	285	180
rect	284	180	285	181
rect	284	181	285	182
rect	284	182	285	183
rect	284	183	285	184
rect	284	185	285	186
rect	284	186	285	187
rect	284	188	285	189
rect	284	189	285	190
rect	284	190	285	191
rect	284	191	285	192
rect	284	192	285	193
rect	284	193	285	194
rect	284	194	285	195
rect	284	195	285	196
rect	286	53	287	54
rect	286	54	287	55
rect	286	56	287	57
rect	286	57	287	58
rect	286	58	287	59
rect	286	59	287	60
rect	286	60	287	61
rect	286	62	287	63
rect	286	63	287	64
rect	286	65	287	66
rect	286	66	287	67
rect	286	67	287	68
rect	286	68	287	69
rect	286	69	287	70
rect	286	70	287	71
rect	286	71	287	72
rect	286	72	287	73
rect	286	73	287	74
rect	286	74	287	75
rect	286	75	287	76
rect	286	76	287	77
rect	286	77	287	78
rect	286	78	287	79
rect	286	80	287	81
rect	286	81	287	82
rect	286	83	287	84
rect	286	84	287	85
rect	286	86	287	87
rect	286	87	287	88
rect	286	89	287	90
rect	286	90	287	91
rect	286	91	287	92
rect	286	92	287	93
rect	286	93	287	94
rect	286	94	287	95
rect	286	95	287	96
rect	286	96	287	97
rect	286	97	287	98
rect	286	98	287	99
rect	286	99	287	100
rect	286	100	287	101
rect	286	101	287	102
rect	286	102	287	103
rect	286	103	287	104
rect	286	104	287	105
rect	286	105	287	106
rect	286	106	287	107
rect	286	107	287	108
rect	286	108	287	109
rect	286	110	287	111
rect	286	111	287	112
rect	286	112	287	113
rect	286	113	287	114
rect	286	114	287	115
rect	286	116	287	117
rect	286	117	287	118
rect	286	119	287	120
rect	286	120	287	121
rect	286	121	287	122
rect	286	122	287	123
rect	286	123	287	124
rect	286	125	287	126
rect	286	126	287	127
rect	286	127	287	128
rect	286	128	287	129
rect	286	129	287	130
rect	286	130	287	131
rect	286	131	287	132
rect	286	132	287	133
rect	286	134	287	135
rect	286	135	287	136
rect	286	137	287	138
rect	286	138	287	139
rect	286	140	287	141
rect	286	141	287	142
rect	286	142	287	143
rect	286	143	287	144
rect	286	144	287	145
rect	286	145	287	146
rect	286	146	287	147
rect	286	147	287	148
rect	286	149	287	150
rect	286	150	287	151
rect	286	152	287	153
rect	286	153	287	154
rect	286	154	287	155
rect	286	155	287	156
rect	286	156	287	157
rect	286	158	287	159
rect	286	159	287	160
rect	286	161	287	162
rect	286	162	287	163
rect	286	164	287	165
rect	286	165	287	166
rect	286	167	287	168
rect	286	168	287	169
rect	286	170	287	171
rect	286	171	287	172
rect	286	173	287	174
rect	286	174	287	175
rect	286	176	287	177
rect	286	177	287	178
rect	286	179	287	180
rect	286	180	287	181
rect	286	181	287	182
rect	286	182	287	183
rect	286	183	287	184
rect	286	185	287	186
rect	286	186	287	187
rect	286	188	287	189
rect	286	189	287	190
rect	286	190	287	191
rect	286	191	287	192
rect	286	192	287	193
rect	286	193	287	194
rect	286	194	287	195
rect	286	195	287	196
rect	286	197	287	198
rect	286	198	287	199
rect	286	199	287	200
rect	286	200	287	201
rect	286	201	287	202
rect	286	202	287	203
rect	286	203	287	204
rect	286	204	287	205
rect	286	205	287	206
rect	286	206	287	207
rect	286	207	287	208
rect	286	208	287	209
rect	286	209	287	210
rect	286	210	287	211
rect	286	211	287	212
rect	286	212	287	213
rect	286	213	287	214
rect	286	214	287	215
rect	286	215	287	216
rect	286	216	287	217
rect	295	5	296	6
rect	295	6	296	7
rect	295	14	296	15
rect	295	15	296	16
rect	295	16	296	17
rect	295	17	296	18
rect	295	18	296	19
rect	295	44	296	45
rect	295	45	296	46
rect	295	80	296	81
rect	295	81	296	82
rect	295	149	296	150
rect	295	150	296	151
rect	295	152	296	153
rect	295	153	296	154
rect	304	89	305	90
rect	304	90	305	91
rect	304	91	305	92
rect	304	92	305	93
rect	304	93	305	94
rect	304	94	305	95
rect	304	95	305	96
rect	304	96	305	97
rect	304	97	305	98
rect	304	98	305	99
rect	304	99	305	100
rect	304	100	305	101
rect	304	101	305	102
rect	304	102	305	103
rect	304	103	305	104
rect	304	104	305	105
rect	304	105	305	106
rect	304	106	305	107
rect	304	107	305	108
rect	304	108	305	109
rect	304	109	305	110
rect	304	110	305	111
rect	304	111	305	112
rect	304	112	305	113
rect	304	113	305	114
rect	304	114	305	115
rect	304	125	305	126
rect	304	126	305	127
rect	304	127	305	128
rect	304	128	305	129
rect	304	129	305	130
rect	304	140	305	141
rect	304	141	305	142
rect	306	5	307	6
rect	306	6	307	7
rect	306	26	307	27
rect	306	27	307	28
rect	306	83	307	84
rect	306	84	307	85
rect	306	85	307	86
rect	306	86	307	87
rect	306	87	307	88
rect	306	89	307	90
rect	306	90	307	91
rect	306	91	307	92
rect	306	92	307	93
rect	306	93	307	94
rect	306	94	307	95
rect	306	95	307	96
rect	306	96	307	97
rect	306	97	307	98
rect	306	98	307	99
rect	306	99	307	100
rect	306	100	307	101
rect	306	101	307	102
rect	306	102	307	103
rect	306	103	307	104
rect	306	104	307	105
rect	306	105	307	106
rect	306	106	307	107
rect	306	107	307	108
rect	306	108	307	109
rect	306	109	307	110
rect	306	110	307	111
rect	306	111	307	112
rect	306	112	307	113
rect	306	113	307	114
rect	306	114	307	115
rect	306	116	307	117
rect	306	117	307	118
rect	306	118	307	119
rect	306	119	307	120
rect	306	120	307	121
rect	306	121	307	122
rect	306	122	307	123
rect	306	123	307	124
rect	306	125	307	126
rect	306	126	307	127
rect	306	127	307	128
rect	306	128	307	129
rect	306	129	307	130
rect	306	131	307	132
rect	306	132	307	133
rect	306	133	307	134
rect	306	134	307	135
rect	306	135	307	136
rect	306	136	307	137
rect	306	137	307	138
rect	306	138	307	139
rect	306	140	307	141
rect	306	141	307	142
rect	306	143	307	144
rect	306	144	307	145
rect	306	145	307	146
rect	306	146	307	147
rect	306	147	307	148
rect	306	148	307	149
rect	306	149	307	150
rect	306	150	307	151
rect	306	151	307	152
rect	306	152	307	153
rect	306	153	307	154
rect	306	154	307	155
rect	306	155	307	156
rect	306	156	307	157
rect	306	157	307	158
rect	306	158	307	159
rect	306	159	307	160
rect	306	160	307	161
rect	306	161	307	162
rect	306	162	307	163
rect	306	163	307	164
rect	306	164	307	165
rect	306	165	307	166
<< metal2 >>
rect	1	121	2	122
rect	1	172	2	173
rect	2	121	3	122
rect	2	172	3	173
rect	3	52	4	53
rect	3	58	4	59
rect	3	109	4	110
rect	3	115	4	116
rect	3	118	4	119
rect	3	121	4	122
rect	3	124	4	125
rect	3	136	4	137
rect	3	145	4	146
rect	3	172	4	173
rect	4	52	5	53
rect	4	58	5	59
rect	4	109	5	110
rect	4	115	5	116
rect	4	118	5	119
rect	4	121	5	122
rect	4	124	5	125
rect	4	136	5	137
rect	4	145	5	146
rect	4	172	5	173
rect	5	7	6	8
rect	5	52	6	53
rect	5	58	6	59
rect	5	79	6	80
rect	5	85	6	86
rect	5	91	6	92
rect	5	106	6	107
rect	5	109	6	110
rect	5	115	6	116
rect	5	118	6	119
rect	5	121	6	122
rect	5	124	6	125
rect	5	136	6	137
rect	5	142	6	143
rect	5	145	6	146
rect	5	172	6	173
rect	6	94	7	95
rect	6	115	7	116
rect	6	163	7	164
rect	6	367	7	368
rect	7	1	8	2
rect	7	4	8	5
rect	7	7	8	8
rect	7	10	8	11
rect	7	13	8	14
rect	7	16	8	17
rect	7	19	8	20
rect	7	22	8	23
rect	7	25	8	26
rect	7	28	8	29
rect	7	31	8	32
rect	7	34	8	35
rect	7	37	8	38
rect	7	40	8	41
rect	7	43	8	44
rect	7	46	8	47
rect	7	49	8	50
rect	7	52	8	53
rect	7	55	8	56
rect	7	58	8	59
rect	7	61	8	62
rect	7	64	8	65
rect	7	67	8	68
rect	7	70	8	71
rect	7	73	8	74
rect	7	76	8	77
rect	7	79	8	80
rect	7	82	8	83
rect	7	85	8	86
rect	7	88	8	89
rect	7	91	8	92
rect	7	94	8	95
rect	7	97	8	98
rect	7	100	8	101
rect	7	103	8	104
rect	7	106	8	107
rect	7	109	8	110
rect	7	112	8	113
rect	7	115	8	116
rect	7	118	8	119
rect	7	121	8	122
rect	7	124	8	125
rect	7	127	8	128
rect	7	130	8	131
rect	7	133	8	134
rect	7	136	8	137
rect	7	139	8	140
rect	7	142	8	143
rect	7	145	8	146
rect	7	148	8	149
rect	7	151	8	152
rect	7	154	8	155
rect	7	157	8	158
rect	7	160	8	161
rect	7	163	8	164
rect	7	166	8	167
rect	7	169	8	170
rect	7	172	8	173
rect	7	175	8	176
rect	7	178	8	179
rect	7	181	8	182
rect	7	184	8	185
rect	7	187	8	188
rect	7	190	8	191
rect	7	193	8	194
rect	7	196	8	197
rect	7	199	8	200
rect	7	202	8	203
rect	7	205	8	206
rect	7	208	8	209
rect	7	211	8	212
rect	7	214	8	215
rect	7	217	8	218
rect	7	220	8	221
rect	7	223	8	224
rect	7	226	8	227
rect	7	229	8	230
rect	7	232	8	233
rect	7	235	8	236
rect	7	238	8	239
rect	7	241	8	242
rect	7	244	8	245
rect	7	247	8	248
rect	7	250	8	251
rect	7	253	8	254
rect	7	256	8	257
rect	7	259	8	260
rect	7	262	8	263
rect	7	265	8	266
rect	7	268	8	269
rect	7	271	8	272
rect	7	274	8	275
rect	7	277	8	278
rect	7	280	8	281
rect	7	283	8	284
rect	7	286	8	287
rect	7	289	8	290
rect	7	292	8	293
rect	7	295	8	296
rect	7	298	8	299
rect	7	301	8	302
rect	7	304	8	305
rect	7	307	8	308
rect	7	310	8	311
rect	7	313	8	314
rect	7	316	8	317
rect	7	319	8	320
rect	7	322	8	323
rect	7	325	8	326
rect	7	328	8	329
rect	7	331	8	332
rect	7	334	8	335
rect	7	337	8	338
rect	7	340	8	341
rect	7	343	8	344
rect	7	346	8	347
rect	7	349	8	350
rect	7	352	8	353
rect	7	355	8	356
rect	7	358	8	359
rect	7	361	8	362
rect	7	364	8	365
rect	7	367	8	368
rect	7	373	8	374
rect	7	376	8	377
rect	7	379	8	380
rect	7	385	8	386
rect	8	1	9	2
rect	8	4	9	5
rect	8	7	9	8
rect	8	10	9	11
rect	8	13	9	14
rect	8	16	9	17
rect	8	19	9	20
rect	8	22	9	23
rect	8	25	9	26
rect	8	28	9	29
rect	8	31	9	32
rect	8	34	9	35
rect	8	37	9	38
rect	8	40	9	41
rect	8	43	9	44
rect	8	46	9	47
rect	8	49	9	50
rect	8	52	9	53
rect	8	55	9	56
rect	8	58	9	59
rect	8	61	9	62
rect	8	64	9	65
rect	8	67	9	68
rect	8	70	9	71
rect	8	73	9	74
rect	8	76	9	77
rect	8	79	9	80
rect	8	82	9	83
rect	8	85	9	86
rect	8	88	9	89
rect	8	91	9	92
rect	8	94	9	95
rect	8	97	9	98
rect	8	100	9	101
rect	8	103	9	104
rect	8	106	9	107
rect	8	109	9	110
rect	8	112	9	113
rect	8	115	9	116
rect	8	118	9	119
rect	8	121	9	122
rect	8	124	9	125
rect	8	127	9	128
rect	8	130	9	131
rect	8	133	9	134
rect	8	136	9	137
rect	8	139	9	140
rect	8	142	9	143
rect	8	145	9	146
rect	8	148	9	149
rect	8	151	9	152
rect	8	154	9	155
rect	8	157	9	158
rect	8	160	9	161
rect	8	163	9	164
rect	8	166	9	167
rect	8	169	9	170
rect	8	172	9	173
rect	8	175	9	176
rect	8	178	9	179
rect	8	181	9	182
rect	8	184	9	185
rect	8	187	9	188
rect	8	190	9	191
rect	8	193	9	194
rect	8	196	9	197
rect	8	199	9	200
rect	8	202	9	203
rect	8	205	9	206
rect	8	208	9	209
rect	8	211	9	212
rect	8	214	9	215
rect	8	217	9	218
rect	8	220	9	221
rect	8	223	9	224
rect	8	226	9	227
rect	8	229	9	230
rect	8	232	9	233
rect	8	235	9	236
rect	8	238	9	239
rect	8	241	9	242
rect	8	244	9	245
rect	8	247	9	248
rect	8	250	9	251
rect	8	253	9	254
rect	8	256	9	257
rect	8	259	9	260
rect	8	262	9	263
rect	8	265	9	266
rect	8	268	9	269
rect	8	271	9	272
rect	8	274	9	275
rect	8	277	9	278
rect	8	280	9	281
rect	8	283	9	284
rect	8	286	9	287
rect	8	289	9	290
rect	8	292	9	293
rect	8	295	9	296
rect	8	298	9	299
rect	8	301	9	302
rect	8	304	9	305
rect	8	307	9	308
rect	8	310	9	311
rect	8	313	9	314
rect	8	316	9	317
rect	8	319	9	320
rect	8	322	9	323
rect	8	325	9	326
rect	8	328	9	329
rect	8	331	9	332
rect	8	334	9	335
rect	8	337	9	338
rect	8	340	9	341
rect	8	343	9	344
rect	8	346	9	347
rect	8	349	9	350
rect	8	352	9	353
rect	8	355	9	356
rect	8	358	9	359
rect	8	361	9	362
rect	8	364	9	365
rect	8	367	9	368
rect	8	373	9	374
rect	8	376	9	377
rect	8	379	9	380
rect	8	385	9	386
rect	9	1	10	2
rect	9	4	10	5
rect	9	7	10	8
rect	9	10	10	11
rect	9	13	10	14
rect	9	16	10	17
rect	9	19	10	20
rect	9	22	10	23
rect	9	25	10	26
rect	9	28	10	29
rect	9	31	10	32
rect	9	34	10	35
rect	9	37	10	38
rect	9	40	10	41
rect	9	43	10	44
rect	9	46	10	47
rect	9	49	10	50
rect	9	52	10	53
rect	9	55	10	56
rect	9	58	10	59
rect	9	61	10	62
rect	9	64	10	65
rect	9	67	10	68
rect	9	70	10	71
rect	9	73	10	74
rect	9	76	10	77
rect	9	79	10	80
rect	9	82	10	83
rect	9	85	10	86
rect	9	88	10	89
rect	9	91	10	92
rect	9	94	10	95
rect	9	97	10	98
rect	9	100	10	101
rect	9	103	10	104
rect	9	106	10	107
rect	9	109	10	110
rect	9	112	10	113
rect	9	115	10	116
rect	9	118	10	119
rect	9	121	10	122
rect	9	124	10	125
rect	9	127	10	128
rect	9	130	10	131
rect	9	133	10	134
rect	9	136	10	137
rect	9	139	10	140
rect	9	142	10	143
rect	9	145	10	146
rect	9	148	10	149
rect	9	151	10	152
rect	9	154	10	155
rect	9	157	10	158
rect	9	160	10	161
rect	9	163	10	164
rect	9	166	10	167
rect	9	169	10	170
rect	9	172	10	173
rect	9	175	10	176
rect	9	178	10	179
rect	9	181	10	182
rect	9	184	10	185
rect	9	187	10	188
rect	9	190	10	191
rect	9	193	10	194
rect	9	196	10	197
rect	9	199	10	200
rect	9	202	10	203
rect	9	205	10	206
rect	9	208	10	209
rect	9	211	10	212
rect	9	214	10	215
rect	9	217	10	218
rect	9	220	10	221
rect	9	223	10	224
rect	9	226	10	227
rect	9	229	10	230
rect	9	232	10	233
rect	9	235	10	236
rect	9	238	10	239
rect	9	241	10	242
rect	9	244	10	245
rect	9	247	10	248
rect	9	250	10	251
rect	9	253	10	254
rect	9	256	10	257
rect	9	259	10	260
rect	9	262	10	263
rect	9	265	10	266
rect	9	268	10	269
rect	9	271	10	272
rect	9	274	10	275
rect	9	277	10	278
rect	9	280	10	281
rect	9	283	10	284
rect	9	286	10	287
rect	9	289	10	290
rect	9	292	10	293
rect	9	295	10	296
rect	9	298	10	299
rect	9	301	10	302
rect	9	304	10	305
rect	9	307	10	308
rect	9	310	10	311
rect	9	313	10	314
rect	9	316	10	317
rect	9	319	10	320
rect	9	322	10	323
rect	9	325	10	326
rect	9	328	10	329
rect	9	331	10	332
rect	9	334	10	335
rect	9	337	10	338
rect	9	340	10	341
rect	9	343	10	344
rect	9	346	10	347
rect	9	349	10	350
rect	9	352	10	353
rect	9	355	10	356
rect	9	358	10	359
rect	9	361	10	362
rect	9	364	10	365
rect	9	367	10	368
rect	9	373	10	374
rect	9	376	10	377
rect	9	379	10	380
rect	9	385	10	386
rect	10	1	11	2
rect	10	4	11	5
rect	10	7	11	8
rect	10	10	11	11
rect	10	13	11	14
rect	10	16	11	17
rect	10	19	11	20
rect	10	22	11	23
rect	10	25	11	26
rect	10	28	11	29
rect	10	31	11	32
rect	10	34	11	35
rect	10	37	11	38
rect	10	40	11	41
rect	10	43	11	44
rect	10	46	11	47
rect	10	49	11	50
rect	10	52	11	53
rect	10	55	11	56
rect	10	58	11	59
rect	10	61	11	62
rect	10	64	11	65
rect	10	67	11	68
rect	10	70	11	71
rect	10	73	11	74
rect	10	76	11	77
rect	10	79	11	80
rect	10	82	11	83
rect	10	85	11	86
rect	10	88	11	89
rect	10	91	11	92
rect	10	94	11	95
rect	10	97	11	98
rect	10	100	11	101
rect	10	103	11	104
rect	10	106	11	107
rect	10	109	11	110
rect	10	112	11	113
rect	10	115	11	116
rect	10	118	11	119
rect	10	121	11	122
rect	10	124	11	125
rect	10	127	11	128
rect	10	130	11	131
rect	10	133	11	134
rect	10	136	11	137
rect	10	139	11	140
rect	10	142	11	143
rect	10	145	11	146
rect	10	148	11	149
rect	10	151	11	152
rect	10	154	11	155
rect	10	157	11	158
rect	10	160	11	161
rect	10	163	11	164
rect	10	166	11	167
rect	10	169	11	170
rect	10	172	11	173
rect	10	175	11	176
rect	10	178	11	179
rect	10	181	11	182
rect	10	184	11	185
rect	10	187	11	188
rect	10	190	11	191
rect	10	193	11	194
rect	10	196	11	197
rect	10	199	11	200
rect	10	202	11	203
rect	10	205	11	206
rect	10	208	11	209
rect	10	211	11	212
rect	10	214	11	215
rect	10	217	11	218
rect	10	220	11	221
rect	10	223	11	224
rect	10	226	11	227
rect	10	229	11	230
rect	10	232	11	233
rect	10	235	11	236
rect	10	238	11	239
rect	10	241	11	242
rect	10	244	11	245
rect	10	247	11	248
rect	10	250	11	251
rect	10	253	11	254
rect	10	256	11	257
rect	10	259	11	260
rect	10	262	11	263
rect	10	265	11	266
rect	10	268	11	269
rect	10	271	11	272
rect	10	274	11	275
rect	10	277	11	278
rect	10	280	11	281
rect	10	283	11	284
rect	10	286	11	287
rect	10	289	11	290
rect	10	292	11	293
rect	10	295	11	296
rect	10	298	11	299
rect	10	301	11	302
rect	10	304	11	305
rect	10	307	11	308
rect	10	310	11	311
rect	10	313	11	314
rect	10	316	11	317
rect	10	319	11	320
rect	10	322	11	323
rect	10	325	11	326
rect	10	328	11	329
rect	10	331	11	332
rect	10	334	11	335
rect	10	337	11	338
rect	10	340	11	341
rect	10	343	11	344
rect	10	346	11	347
rect	10	349	11	350
rect	10	352	11	353
rect	10	355	11	356
rect	10	358	11	359
rect	10	361	11	362
rect	10	364	11	365
rect	10	367	11	368
rect	10	373	11	374
rect	10	376	11	377
rect	10	379	11	380
rect	10	385	11	386
rect	11	1	12	2
rect	11	4	12	5
rect	11	7	12	8
rect	11	10	12	11
rect	11	13	12	14
rect	11	16	12	17
rect	11	19	12	20
rect	11	22	12	23
rect	11	25	12	26
rect	11	28	12	29
rect	11	31	12	32
rect	11	34	12	35
rect	11	37	12	38
rect	11	40	12	41
rect	11	43	12	44
rect	11	46	12	47
rect	11	49	12	50
rect	11	52	12	53
rect	11	55	12	56
rect	11	58	12	59
rect	11	61	12	62
rect	11	64	12	65
rect	11	67	12	68
rect	11	70	12	71
rect	11	73	12	74
rect	11	76	12	77
rect	11	79	12	80
rect	11	82	12	83
rect	11	85	12	86
rect	11	88	12	89
rect	11	91	12	92
rect	11	94	12	95
rect	11	97	12	98
rect	11	100	12	101
rect	11	103	12	104
rect	11	106	12	107
rect	11	109	12	110
rect	11	112	12	113
rect	11	115	12	116
rect	11	118	12	119
rect	11	121	12	122
rect	11	124	12	125
rect	11	127	12	128
rect	11	130	12	131
rect	11	133	12	134
rect	11	136	12	137
rect	11	139	12	140
rect	11	142	12	143
rect	11	145	12	146
rect	11	148	12	149
rect	11	151	12	152
rect	11	154	12	155
rect	11	157	12	158
rect	11	160	12	161
rect	11	163	12	164
rect	11	166	12	167
rect	11	169	12	170
rect	11	172	12	173
rect	11	175	12	176
rect	11	178	12	179
rect	11	181	12	182
rect	11	184	12	185
rect	11	187	12	188
rect	11	190	12	191
rect	11	193	12	194
rect	11	196	12	197
rect	11	199	12	200
rect	11	202	12	203
rect	11	205	12	206
rect	11	208	12	209
rect	11	211	12	212
rect	11	214	12	215
rect	11	217	12	218
rect	11	220	12	221
rect	11	223	12	224
rect	11	226	12	227
rect	11	229	12	230
rect	11	232	12	233
rect	11	235	12	236
rect	11	238	12	239
rect	11	241	12	242
rect	11	244	12	245
rect	11	247	12	248
rect	11	250	12	251
rect	11	253	12	254
rect	11	256	12	257
rect	11	259	12	260
rect	11	262	12	263
rect	11	265	12	266
rect	11	268	12	269
rect	11	271	12	272
rect	11	274	12	275
rect	11	277	12	278
rect	11	280	12	281
rect	11	283	12	284
rect	11	286	12	287
rect	11	289	12	290
rect	11	292	12	293
rect	11	295	12	296
rect	11	298	12	299
rect	11	301	12	302
rect	11	304	12	305
rect	11	307	12	308
rect	11	310	12	311
rect	11	313	12	314
rect	11	316	12	317
rect	11	319	12	320
rect	11	322	12	323
rect	11	325	12	326
rect	11	328	12	329
rect	11	331	12	332
rect	11	334	12	335
rect	11	337	12	338
rect	11	340	12	341
rect	11	343	12	344
rect	11	346	12	347
rect	11	349	12	350
rect	11	352	12	353
rect	11	355	12	356
rect	11	358	12	359
rect	11	361	12	362
rect	11	364	12	365
rect	11	367	12	368
rect	11	373	12	374
rect	11	376	12	377
rect	11	379	12	380
rect	11	385	12	386
rect	12	1	13	2
rect	12	4	13	5
rect	12	7	13	8
rect	12	10	13	11
rect	12	13	13	14
rect	12	16	13	17
rect	12	19	13	20
rect	12	22	13	23
rect	12	25	13	26
rect	12	28	13	29
rect	12	31	13	32
rect	12	34	13	35
rect	12	37	13	38
rect	12	40	13	41
rect	12	43	13	44
rect	12	46	13	47
rect	12	49	13	50
rect	12	52	13	53
rect	12	55	13	56
rect	12	58	13	59
rect	12	61	13	62
rect	12	64	13	65
rect	12	67	13	68
rect	12	70	13	71
rect	12	73	13	74
rect	12	76	13	77
rect	12	79	13	80
rect	12	82	13	83
rect	12	85	13	86
rect	12	88	13	89
rect	12	91	13	92
rect	12	94	13	95
rect	12	97	13	98
rect	12	100	13	101
rect	12	103	13	104
rect	12	106	13	107
rect	12	109	13	110
rect	12	112	13	113
rect	12	115	13	116
rect	12	118	13	119
rect	12	121	13	122
rect	12	124	13	125
rect	12	127	13	128
rect	12	130	13	131
rect	12	133	13	134
rect	12	136	13	137
rect	12	139	13	140
rect	12	142	13	143
rect	12	145	13	146
rect	12	148	13	149
rect	12	151	13	152
rect	12	154	13	155
rect	12	157	13	158
rect	12	160	13	161
rect	12	163	13	164
rect	12	166	13	167
rect	12	169	13	170
rect	12	172	13	173
rect	12	175	13	176
rect	12	178	13	179
rect	12	181	13	182
rect	12	184	13	185
rect	12	187	13	188
rect	12	190	13	191
rect	12	193	13	194
rect	12	196	13	197
rect	12	199	13	200
rect	12	202	13	203
rect	12	205	13	206
rect	12	208	13	209
rect	12	211	13	212
rect	12	214	13	215
rect	12	217	13	218
rect	12	220	13	221
rect	12	223	13	224
rect	12	226	13	227
rect	12	229	13	230
rect	12	232	13	233
rect	12	235	13	236
rect	12	238	13	239
rect	12	241	13	242
rect	12	244	13	245
rect	12	247	13	248
rect	12	250	13	251
rect	12	253	13	254
rect	12	256	13	257
rect	12	259	13	260
rect	12	262	13	263
rect	12	265	13	266
rect	12	268	13	269
rect	12	271	13	272
rect	12	274	13	275
rect	12	277	13	278
rect	12	280	13	281
rect	12	283	13	284
rect	12	286	13	287
rect	12	289	13	290
rect	12	292	13	293
rect	12	295	13	296
rect	12	298	13	299
rect	12	301	13	302
rect	12	304	13	305
rect	12	307	13	308
rect	12	310	13	311
rect	12	313	13	314
rect	12	316	13	317
rect	12	319	13	320
rect	12	322	13	323
rect	12	325	13	326
rect	12	328	13	329
rect	12	331	13	332
rect	12	334	13	335
rect	12	337	13	338
rect	12	340	13	341
rect	12	343	13	344
rect	12	346	13	347
rect	12	349	13	350
rect	12	352	13	353
rect	12	355	13	356
rect	12	358	13	359
rect	12	361	13	362
rect	12	364	13	365
rect	12	367	13	368
rect	12	373	13	374
rect	12	376	13	377
rect	12	379	13	380
rect	12	385	13	386
rect	13	1	14	2
rect	13	4	14	5
rect	13	7	14	8
rect	13	10	14	11
rect	13	13	14	14
rect	13	16	14	17
rect	13	19	14	20
rect	13	22	14	23
rect	13	25	14	26
rect	13	28	14	29
rect	13	31	14	32
rect	13	34	14	35
rect	13	37	14	38
rect	13	40	14	41
rect	13	43	14	44
rect	13	46	14	47
rect	13	49	14	50
rect	13	52	14	53
rect	13	55	14	56
rect	13	58	14	59
rect	13	61	14	62
rect	13	64	14	65
rect	13	67	14	68
rect	13	70	14	71
rect	13	73	14	74
rect	13	76	14	77
rect	13	79	14	80
rect	13	82	14	83
rect	13	85	14	86
rect	13	88	14	89
rect	13	91	14	92
rect	13	94	14	95
rect	13	97	14	98
rect	13	100	14	101
rect	13	103	14	104
rect	13	106	14	107
rect	13	109	14	110
rect	13	112	14	113
rect	13	115	14	116
rect	13	118	14	119
rect	13	121	14	122
rect	13	124	14	125
rect	13	127	14	128
rect	13	130	14	131
rect	13	133	14	134
rect	13	136	14	137
rect	13	139	14	140
rect	13	142	14	143
rect	13	145	14	146
rect	13	148	14	149
rect	13	151	14	152
rect	13	154	14	155
rect	13	157	14	158
rect	13	160	14	161
rect	13	163	14	164
rect	13	166	14	167
rect	13	169	14	170
rect	13	172	14	173
rect	13	175	14	176
rect	13	178	14	179
rect	13	181	14	182
rect	13	184	14	185
rect	13	187	14	188
rect	13	190	14	191
rect	13	193	14	194
rect	13	196	14	197
rect	13	199	14	200
rect	13	202	14	203
rect	13	205	14	206
rect	13	208	14	209
rect	13	211	14	212
rect	13	214	14	215
rect	13	217	14	218
rect	13	220	14	221
rect	13	223	14	224
rect	13	226	14	227
rect	13	229	14	230
rect	13	232	14	233
rect	13	235	14	236
rect	13	238	14	239
rect	13	241	14	242
rect	13	244	14	245
rect	13	247	14	248
rect	13	250	14	251
rect	13	253	14	254
rect	13	256	14	257
rect	13	259	14	260
rect	13	262	14	263
rect	13	265	14	266
rect	13	268	14	269
rect	13	271	14	272
rect	13	274	14	275
rect	13	277	14	278
rect	13	280	14	281
rect	13	283	14	284
rect	13	286	14	287
rect	13	289	14	290
rect	13	292	14	293
rect	13	295	14	296
rect	13	298	14	299
rect	13	301	14	302
rect	13	304	14	305
rect	13	307	14	308
rect	13	310	14	311
rect	13	313	14	314
rect	13	316	14	317
rect	13	319	14	320
rect	13	322	14	323
rect	13	325	14	326
rect	13	328	14	329
rect	13	331	14	332
rect	13	334	14	335
rect	13	337	14	338
rect	13	340	14	341
rect	13	343	14	344
rect	13	346	14	347
rect	13	349	14	350
rect	13	352	14	353
rect	13	355	14	356
rect	13	358	14	359
rect	13	361	14	362
rect	13	364	14	365
rect	13	367	14	368
rect	13	373	14	374
rect	13	376	14	377
rect	13	379	14	380
rect	13	385	14	386
rect	14	1	15	2
rect	14	4	15	5
rect	14	7	15	8
rect	14	10	15	11
rect	14	13	15	14
rect	14	16	15	17
rect	14	19	15	20
rect	14	22	15	23
rect	14	25	15	26
rect	14	28	15	29
rect	14	31	15	32
rect	14	34	15	35
rect	14	37	15	38
rect	14	40	15	41
rect	14	43	15	44
rect	14	46	15	47
rect	14	49	15	50
rect	14	52	15	53
rect	14	55	15	56
rect	14	58	15	59
rect	14	61	15	62
rect	14	64	15	65
rect	14	67	15	68
rect	14	70	15	71
rect	14	73	15	74
rect	14	76	15	77
rect	14	79	15	80
rect	14	82	15	83
rect	14	85	15	86
rect	14	88	15	89
rect	14	91	15	92
rect	14	94	15	95
rect	14	97	15	98
rect	14	100	15	101
rect	14	103	15	104
rect	14	106	15	107
rect	14	109	15	110
rect	14	112	15	113
rect	14	115	15	116
rect	14	118	15	119
rect	14	121	15	122
rect	14	124	15	125
rect	14	127	15	128
rect	14	130	15	131
rect	14	133	15	134
rect	14	136	15	137
rect	14	139	15	140
rect	14	142	15	143
rect	14	145	15	146
rect	14	148	15	149
rect	14	151	15	152
rect	14	154	15	155
rect	14	157	15	158
rect	14	160	15	161
rect	14	163	15	164
rect	14	166	15	167
rect	14	169	15	170
rect	14	172	15	173
rect	14	175	15	176
rect	14	178	15	179
rect	14	181	15	182
rect	14	184	15	185
rect	14	187	15	188
rect	14	190	15	191
rect	14	193	15	194
rect	14	196	15	197
rect	14	199	15	200
rect	14	202	15	203
rect	14	205	15	206
rect	14	208	15	209
rect	14	211	15	212
rect	14	214	15	215
rect	14	217	15	218
rect	14	220	15	221
rect	14	223	15	224
rect	14	226	15	227
rect	14	229	15	230
rect	14	232	15	233
rect	14	235	15	236
rect	14	238	15	239
rect	14	241	15	242
rect	14	244	15	245
rect	14	247	15	248
rect	14	250	15	251
rect	14	253	15	254
rect	14	256	15	257
rect	14	259	15	260
rect	14	262	15	263
rect	14	265	15	266
rect	14	268	15	269
rect	14	271	15	272
rect	14	274	15	275
rect	14	277	15	278
rect	14	280	15	281
rect	14	283	15	284
rect	14	286	15	287
rect	14	289	15	290
rect	14	292	15	293
rect	14	295	15	296
rect	14	298	15	299
rect	14	301	15	302
rect	14	304	15	305
rect	14	307	15	308
rect	14	310	15	311
rect	14	313	15	314
rect	14	316	15	317
rect	14	319	15	320
rect	14	322	15	323
rect	14	325	15	326
rect	14	328	15	329
rect	14	331	15	332
rect	14	334	15	335
rect	14	337	15	338
rect	14	340	15	341
rect	14	343	15	344
rect	14	346	15	347
rect	14	349	15	350
rect	14	352	15	353
rect	14	355	15	356
rect	14	358	15	359
rect	14	361	15	362
rect	14	364	15	365
rect	14	367	15	368
rect	14	373	15	374
rect	14	376	15	377
rect	14	379	15	380
rect	14	385	15	386
rect	15	1	16	2
rect	15	4	16	5
rect	15	7	16	8
rect	15	10	16	11
rect	15	13	16	14
rect	15	16	16	17
rect	15	19	16	20
rect	15	22	16	23
rect	15	25	16	26
rect	15	28	16	29
rect	15	31	16	32
rect	15	34	16	35
rect	15	37	16	38
rect	15	40	16	41
rect	15	43	16	44
rect	15	46	16	47
rect	15	49	16	50
rect	15	52	16	53
rect	15	55	16	56
rect	15	58	16	59
rect	15	61	16	62
rect	15	64	16	65
rect	15	67	16	68
rect	15	70	16	71
rect	15	73	16	74
rect	15	76	16	77
rect	15	79	16	80
rect	15	82	16	83
rect	15	85	16	86
rect	15	88	16	89
rect	15	91	16	92
rect	15	94	16	95
rect	15	97	16	98
rect	15	100	16	101
rect	15	103	16	104
rect	15	106	16	107
rect	15	109	16	110
rect	15	112	16	113
rect	15	115	16	116
rect	15	118	16	119
rect	15	121	16	122
rect	15	124	16	125
rect	15	127	16	128
rect	15	130	16	131
rect	15	133	16	134
rect	15	136	16	137
rect	15	139	16	140
rect	15	142	16	143
rect	15	145	16	146
rect	15	148	16	149
rect	15	151	16	152
rect	15	154	16	155
rect	15	157	16	158
rect	15	160	16	161
rect	15	163	16	164
rect	15	166	16	167
rect	15	169	16	170
rect	15	172	16	173
rect	15	175	16	176
rect	15	178	16	179
rect	15	181	16	182
rect	15	184	16	185
rect	15	187	16	188
rect	15	190	16	191
rect	15	193	16	194
rect	15	196	16	197
rect	15	199	16	200
rect	15	202	16	203
rect	15	205	16	206
rect	15	208	16	209
rect	15	211	16	212
rect	15	214	16	215
rect	15	217	16	218
rect	15	220	16	221
rect	15	223	16	224
rect	15	226	16	227
rect	15	229	16	230
rect	15	232	16	233
rect	15	235	16	236
rect	15	238	16	239
rect	15	241	16	242
rect	15	244	16	245
rect	15	247	16	248
rect	15	250	16	251
rect	15	253	16	254
rect	15	256	16	257
rect	15	259	16	260
rect	15	262	16	263
rect	15	265	16	266
rect	15	268	16	269
rect	15	271	16	272
rect	15	274	16	275
rect	15	277	16	278
rect	15	280	16	281
rect	15	283	16	284
rect	15	286	16	287
rect	15	289	16	290
rect	15	292	16	293
rect	15	295	16	296
rect	15	298	16	299
rect	15	301	16	302
rect	15	304	16	305
rect	15	307	16	308
rect	15	310	16	311
rect	15	313	16	314
rect	15	316	16	317
rect	15	319	16	320
rect	15	322	16	323
rect	15	325	16	326
rect	15	328	16	329
rect	15	331	16	332
rect	15	334	16	335
rect	15	337	16	338
rect	15	340	16	341
rect	15	343	16	344
rect	15	346	16	347
rect	15	349	16	350
rect	15	352	16	353
rect	15	355	16	356
rect	15	358	16	359
rect	15	361	16	362
rect	15	364	16	365
rect	15	367	16	368
rect	15	373	16	374
rect	15	376	16	377
rect	15	379	16	380
rect	15	385	16	386
rect	16	1	17	2
rect	16	4	17	5
rect	16	7	17	8
rect	16	10	17	11
rect	16	13	17	14
rect	16	16	17	17
rect	16	19	17	20
rect	16	22	17	23
rect	16	25	17	26
rect	16	28	17	29
rect	16	31	17	32
rect	16	34	17	35
rect	16	37	17	38
rect	16	40	17	41
rect	16	43	17	44
rect	16	46	17	47
rect	16	49	17	50
rect	16	52	17	53
rect	16	55	17	56
rect	16	58	17	59
rect	16	61	17	62
rect	16	64	17	65
rect	16	67	17	68
rect	16	70	17	71
rect	16	73	17	74
rect	16	76	17	77
rect	16	79	17	80
rect	16	82	17	83
rect	16	85	17	86
rect	16	88	17	89
rect	16	91	17	92
rect	16	94	17	95
rect	16	97	17	98
rect	16	100	17	101
rect	16	103	17	104
rect	16	106	17	107
rect	16	109	17	110
rect	16	112	17	113
rect	16	115	17	116
rect	16	118	17	119
rect	16	121	17	122
rect	16	124	17	125
rect	16	127	17	128
rect	16	130	17	131
rect	16	133	17	134
rect	16	136	17	137
rect	16	139	17	140
rect	16	142	17	143
rect	16	145	17	146
rect	16	148	17	149
rect	16	151	17	152
rect	16	154	17	155
rect	16	157	17	158
rect	16	160	17	161
rect	16	163	17	164
rect	16	166	17	167
rect	16	169	17	170
rect	16	172	17	173
rect	16	175	17	176
rect	16	178	17	179
rect	16	181	17	182
rect	16	184	17	185
rect	16	187	17	188
rect	16	190	17	191
rect	16	193	17	194
rect	16	196	17	197
rect	16	199	17	200
rect	16	202	17	203
rect	16	205	17	206
rect	16	208	17	209
rect	16	211	17	212
rect	16	214	17	215
rect	16	217	17	218
rect	16	220	17	221
rect	16	223	17	224
rect	16	226	17	227
rect	16	229	17	230
rect	16	232	17	233
rect	16	235	17	236
rect	16	238	17	239
rect	16	241	17	242
rect	16	244	17	245
rect	16	247	17	248
rect	16	250	17	251
rect	16	253	17	254
rect	16	256	17	257
rect	16	259	17	260
rect	16	262	17	263
rect	16	265	17	266
rect	16	268	17	269
rect	16	271	17	272
rect	16	274	17	275
rect	16	277	17	278
rect	16	280	17	281
rect	16	283	17	284
rect	16	286	17	287
rect	16	289	17	290
rect	16	292	17	293
rect	16	295	17	296
rect	16	298	17	299
rect	16	301	17	302
rect	16	304	17	305
rect	16	307	17	308
rect	16	310	17	311
rect	16	313	17	314
rect	16	316	17	317
rect	16	319	17	320
rect	16	322	17	323
rect	16	325	17	326
rect	16	328	17	329
rect	16	331	17	332
rect	16	334	17	335
rect	16	337	17	338
rect	16	340	17	341
rect	16	343	17	344
rect	16	346	17	347
rect	16	349	17	350
rect	16	352	17	353
rect	16	355	17	356
rect	16	358	17	359
rect	16	361	17	362
rect	16	364	17	365
rect	16	367	17	368
rect	16	373	17	374
rect	16	376	17	377
rect	16	379	17	380
rect	16	385	17	386
rect	17	1	18	2
rect	17	4	18	5
rect	17	7	18	8
rect	17	10	18	11
rect	17	13	18	14
rect	17	16	18	17
rect	17	19	18	20
rect	17	22	18	23
rect	17	25	18	26
rect	17	28	18	29
rect	17	31	18	32
rect	17	34	18	35
rect	17	37	18	38
rect	17	40	18	41
rect	17	43	18	44
rect	17	46	18	47
rect	17	49	18	50
rect	17	52	18	53
rect	17	55	18	56
rect	17	58	18	59
rect	17	61	18	62
rect	17	64	18	65
rect	17	67	18	68
rect	17	70	18	71
rect	17	73	18	74
rect	17	76	18	77
rect	17	79	18	80
rect	17	82	18	83
rect	17	85	18	86
rect	17	88	18	89
rect	17	91	18	92
rect	17	94	18	95
rect	17	97	18	98
rect	17	100	18	101
rect	17	103	18	104
rect	17	106	18	107
rect	17	109	18	110
rect	17	112	18	113
rect	17	115	18	116
rect	17	118	18	119
rect	17	121	18	122
rect	17	124	18	125
rect	17	127	18	128
rect	17	130	18	131
rect	17	133	18	134
rect	17	136	18	137
rect	17	139	18	140
rect	17	142	18	143
rect	17	145	18	146
rect	17	148	18	149
rect	17	151	18	152
rect	17	154	18	155
rect	17	157	18	158
rect	17	160	18	161
rect	17	163	18	164
rect	17	166	18	167
rect	17	169	18	170
rect	17	172	18	173
rect	17	175	18	176
rect	17	178	18	179
rect	17	181	18	182
rect	17	184	18	185
rect	17	187	18	188
rect	17	190	18	191
rect	17	193	18	194
rect	17	196	18	197
rect	17	199	18	200
rect	17	202	18	203
rect	17	205	18	206
rect	17	208	18	209
rect	17	211	18	212
rect	17	214	18	215
rect	17	217	18	218
rect	17	220	18	221
rect	17	223	18	224
rect	17	226	18	227
rect	17	229	18	230
rect	17	232	18	233
rect	17	235	18	236
rect	17	238	18	239
rect	17	241	18	242
rect	17	244	18	245
rect	17	247	18	248
rect	17	250	18	251
rect	17	253	18	254
rect	17	256	18	257
rect	17	259	18	260
rect	17	262	18	263
rect	17	265	18	266
rect	17	268	18	269
rect	17	271	18	272
rect	17	274	18	275
rect	17	277	18	278
rect	17	280	18	281
rect	17	283	18	284
rect	17	286	18	287
rect	17	289	18	290
rect	17	292	18	293
rect	17	295	18	296
rect	17	298	18	299
rect	17	301	18	302
rect	17	304	18	305
rect	17	307	18	308
rect	17	310	18	311
rect	17	313	18	314
rect	17	316	18	317
rect	17	319	18	320
rect	17	322	18	323
rect	17	325	18	326
rect	17	328	18	329
rect	17	331	18	332
rect	17	334	18	335
rect	17	337	18	338
rect	17	340	18	341
rect	17	343	18	344
rect	17	346	18	347
rect	17	349	18	350
rect	17	352	18	353
rect	17	355	18	356
rect	17	358	18	359
rect	17	361	18	362
rect	17	364	18	365
rect	17	367	18	368
rect	17	373	18	374
rect	17	376	18	377
rect	17	379	18	380
rect	17	385	18	386
rect	18	1	19	2
rect	18	4	19	5
rect	18	7	19	8
rect	18	10	19	11
rect	18	13	19	14
rect	18	16	19	17
rect	18	19	19	20
rect	18	22	19	23
rect	18	25	19	26
rect	18	28	19	29
rect	18	31	19	32
rect	18	34	19	35
rect	18	37	19	38
rect	18	40	19	41
rect	18	43	19	44
rect	18	46	19	47
rect	18	49	19	50
rect	18	52	19	53
rect	18	55	19	56
rect	18	58	19	59
rect	18	61	19	62
rect	18	64	19	65
rect	18	67	19	68
rect	18	70	19	71
rect	18	73	19	74
rect	18	76	19	77
rect	18	79	19	80
rect	18	82	19	83
rect	18	85	19	86
rect	18	88	19	89
rect	18	91	19	92
rect	18	94	19	95
rect	18	97	19	98
rect	18	100	19	101
rect	18	103	19	104
rect	18	106	19	107
rect	18	109	19	110
rect	18	112	19	113
rect	18	115	19	116
rect	18	118	19	119
rect	18	121	19	122
rect	18	124	19	125
rect	18	127	19	128
rect	18	130	19	131
rect	18	133	19	134
rect	18	136	19	137
rect	18	139	19	140
rect	18	142	19	143
rect	18	145	19	146
rect	18	148	19	149
rect	18	151	19	152
rect	18	154	19	155
rect	18	157	19	158
rect	18	160	19	161
rect	18	163	19	164
rect	18	166	19	167
rect	18	169	19	170
rect	18	172	19	173
rect	18	175	19	176
rect	18	178	19	179
rect	18	181	19	182
rect	18	184	19	185
rect	18	187	19	188
rect	18	190	19	191
rect	18	193	19	194
rect	18	196	19	197
rect	18	199	19	200
rect	18	202	19	203
rect	18	205	19	206
rect	18	208	19	209
rect	18	211	19	212
rect	18	214	19	215
rect	18	217	19	218
rect	18	220	19	221
rect	18	223	19	224
rect	18	226	19	227
rect	18	229	19	230
rect	18	232	19	233
rect	18	235	19	236
rect	18	238	19	239
rect	18	241	19	242
rect	18	244	19	245
rect	18	247	19	248
rect	18	250	19	251
rect	18	253	19	254
rect	18	256	19	257
rect	18	259	19	260
rect	18	262	19	263
rect	18	265	19	266
rect	18	268	19	269
rect	18	271	19	272
rect	18	274	19	275
rect	18	277	19	278
rect	18	280	19	281
rect	18	283	19	284
rect	18	286	19	287
rect	18	289	19	290
rect	18	292	19	293
rect	18	295	19	296
rect	18	298	19	299
rect	18	301	19	302
rect	18	304	19	305
rect	18	307	19	308
rect	18	310	19	311
rect	18	313	19	314
rect	18	316	19	317
rect	18	319	19	320
rect	18	322	19	323
rect	18	325	19	326
rect	18	328	19	329
rect	18	331	19	332
rect	18	334	19	335
rect	18	337	19	338
rect	18	340	19	341
rect	18	343	19	344
rect	18	346	19	347
rect	18	349	19	350
rect	18	352	19	353
rect	18	355	19	356
rect	18	358	19	359
rect	18	361	19	362
rect	18	364	19	365
rect	18	367	19	368
rect	18	373	19	374
rect	18	376	19	377
rect	18	379	19	380
rect	18	385	19	386
rect	19	1	20	2
rect	19	4	20	5
rect	19	7	20	8
rect	19	10	20	11
rect	19	13	20	14
rect	19	16	20	17
rect	19	19	20	20
rect	19	22	20	23
rect	19	25	20	26
rect	19	28	20	29
rect	19	31	20	32
rect	19	34	20	35
rect	19	37	20	38
rect	19	40	20	41
rect	19	43	20	44
rect	19	46	20	47
rect	19	49	20	50
rect	19	52	20	53
rect	19	55	20	56
rect	19	58	20	59
rect	19	61	20	62
rect	19	64	20	65
rect	19	67	20	68
rect	19	70	20	71
rect	19	73	20	74
rect	19	76	20	77
rect	19	79	20	80
rect	19	82	20	83
rect	19	85	20	86
rect	19	88	20	89
rect	19	91	20	92
rect	19	94	20	95
rect	19	97	20	98
rect	19	100	20	101
rect	19	103	20	104
rect	19	106	20	107
rect	19	109	20	110
rect	19	112	20	113
rect	19	115	20	116
rect	19	118	20	119
rect	19	121	20	122
rect	19	124	20	125
rect	19	127	20	128
rect	19	130	20	131
rect	19	133	20	134
rect	19	136	20	137
rect	19	139	20	140
rect	19	142	20	143
rect	19	145	20	146
rect	19	148	20	149
rect	19	151	20	152
rect	19	154	20	155
rect	19	157	20	158
rect	19	160	20	161
rect	19	163	20	164
rect	19	166	20	167
rect	19	169	20	170
rect	19	172	20	173
rect	19	175	20	176
rect	19	178	20	179
rect	19	181	20	182
rect	19	184	20	185
rect	19	187	20	188
rect	19	190	20	191
rect	19	193	20	194
rect	19	196	20	197
rect	19	199	20	200
rect	19	202	20	203
rect	19	205	20	206
rect	19	208	20	209
rect	19	211	20	212
rect	19	214	20	215
rect	19	217	20	218
rect	19	220	20	221
rect	19	223	20	224
rect	19	226	20	227
rect	19	229	20	230
rect	19	232	20	233
rect	19	235	20	236
rect	19	238	20	239
rect	19	241	20	242
rect	19	244	20	245
rect	19	247	20	248
rect	19	250	20	251
rect	19	253	20	254
rect	19	256	20	257
rect	19	259	20	260
rect	19	262	20	263
rect	19	265	20	266
rect	19	268	20	269
rect	19	271	20	272
rect	19	274	20	275
rect	19	277	20	278
rect	19	280	20	281
rect	19	283	20	284
rect	19	286	20	287
rect	19	289	20	290
rect	19	292	20	293
rect	19	295	20	296
rect	19	298	20	299
rect	19	301	20	302
rect	19	304	20	305
rect	19	307	20	308
rect	19	310	20	311
rect	19	313	20	314
rect	19	316	20	317
rect	19	319	20	320
rect	19	322	20	323
rect	19	325	20	326
rect	19	328	20	329
rect	19	331	20	332
rect	19	334	20	335
rect	19	337	20	338
rect	19	340	20	341
rect	19	343	20	344
rect	19	346	20	347
rect	19	349	20	350
rect	19	352	20	353
rect	19	355	20	356
rect	19	358	20	359
rect	19	361	20	362
rect	19	364	20	365
rect	19	367	20	368
rect	19	373	20	374
rect	19	376	20	377
rect	19	379	20	380
rect	19	385	20	386
rect	20	1	21	2
rect	20	4	21	5
rect	20	7	21	8
rect	20	10	21	11
rect	20	13	21	14
rect	20	16	21	17
rect	20	19	21	20
rect	20	22	21	23
rect	20	25	21	26
rect	20	28	21	29
rect	20	31	21	32
rect	20	34	21	35
rect	20	37	21	38
rect	20	40	21	41
rect	20	43	21	44
rect	20	46	21	47
rect	20	49	21	50
rect	20	52	21	53
rect	20	55	21	56
rect	20	58	21	59
rect	20	61	21	62
rect	20	64	21	65
rect	20	67	21	68
rect	20	70	21	71
rect	20	73	21	74
rect	20	76	21	77
rect	20	79	21	80
rect	20	82	21	83
rect	20	85	21	86
rect	20	88	21	89
rect	20	91	21	92
rect	20	94	21	95
rect	20	97	21	98
rect	20	100	21	101
rect	20	103	21	104
rect	20	106	21	107
rect	20	109	21	110
rect	20	112	21	113
rect	20	115	21	116
rect	20	118	21	119
rect	20	121	21	122
rect	20	124	21	125
rect	20	127	21	128
rect	20	130	21	131
rect	20	133	21	134
rect	20	136	21	137
rect	20	139	21	140
rect	20	142	21	143
rect	20	145	21	146
rect	20	148	21	149
rect	20	151	21	152
rect	20	154	21	155
rect	20	157	21	158
rect	20	160	21	161
rect	20	163	21	164
rect	20	166	21	167
rect	20	169	21	170
rect	20	172	21	173
rect	20	175	21	176
rect	20	178	21	179
rect	20	181	21	182
rect	20	184	21	185
rect	20	187	21	188
rect	20	190	21	191
rect	20	193	21	194
rect	20	196	21	197
rect	20	199	21	200
rect	20	202	21	203
rect	20	205	21	206
rect	20	208	21	209
rect	20	211	21	212
rect	20	214	21	215
rect	20	217	21	218
rect	20	220	21	221
rect	20	223	21	224
rect	20	226	21	227
rect	20	229	21	230
rect	20	232	21	233
rect	20	235	21	236
rect	20	238	21	239
rect	20	241	21	242
rect	20	244	21	245
rect	20	247	21	248
rect	20	250	21	251
rect	20	253	21	254
rect	20	256	21	257
rect	20	259	21	260
rect	20	262	21	263
rect	20	265	21	266
rect	20	268	21	269
rect	20	271	21	272
rect	20	274	21	275
rect	20	277	21	278
rect	20	280	21	281
rect	20	283	21	284
rect	20	286	21	287
rect	20	289	21	290
rect	20	292	21	293
rect	20	295	21	296
rect	20	298	21	299
rect	20	301	21	302
rect	20	304	21	305
rect	20	307	21	308
rect	20	310	21	311
rect	20	313	21	314
rect	20	316	21	317
rect	20	319	21	320
rect	20	322	21	323
rect	20	325	21	326
rect	20	328	21	329
rect	20	331	21	332
rect	20	334	21	335
rect	20	337	21	338
rect	20	340	21	341
rect	20	343	21	344
rect	20	346	21	347
rect	20	349	21	350
rect	20	352	21	353
rect	20	355	21	356
rect	20	358	21	359
rect	20	361	21	362
rect	20	364	21	365
rect	20	367	21	368
rect	20	373	21	374
rect	20	376	21	377
rect	20	379	21	380
rect	20	385	21	386
rect	21	1	22	2
rect	21	4	22	5
rect	21	7	22	8
rect	21	10	22	11
rect	21	13	22	14
rect	21	16	22	17
rect	21	19	22	20
rect	21	22	22	23
rect	21	25	22	26
rect	21	28	22	29
rect	21	31	22	32
rect	21	34	22	35
rect	21	37	22	38
rect	21	40	22	41
rect	21	43	22	44
rect	21	46	22	47
rect	21	49	22	50
rect	21	52	22	53
rect	21	55	22	56
rect	21	58	22	59
rect	21	61	22	62
rect	21	64	22	65
rect	21	67	22	68
rect	21	70	22	71
rect	21	73	22	74
rect	21	76	22	77
rect	21	79	22	80
rect	21	82	22	83
rect	21	85	22	86
rect	21	88	22	89
rect	21	91	22	92
rect	21	94	22	95
rect	21	97	22	98
rect	21	100	22	101
rect	21	103	22	104
rect	21	106	22	107
rect	21	109	22	110
rect	21	112	22	113
rect	21	115	22	116
rect	21	118	22	119
rect	21	121	22	122
rect	21	124	22	125
rect	21	127	22	128
rect	21	130	22	131
rect	21	133	22	134
rect	21	136	22	137
rect	21	139	22	140
rect	21	142	22	143
rect	21	145	22	146
rect	21	148	22	149
rect	21	151	22	152
rect	21	154	22	155
rect	21	157	22	158
rect	21	160	22	161
rect	21	163	22	164
rect	21	166	22	167
rect	21	169	22	170
rect	21	172	22	173
rect	21	175	22	176
rect	21	178	22	179
rect	21	181	22	182
rect	21	184	22	185
rect	21	187	22	188
rect	21	190	22	191
rect	21	193	22	194
rect	21	196	22	197
rect	21	199	22	200
rect	21	202	22	203
rect	21	205	22	206
rect	21	208	22	209
rect	21	211	22	212
rect	21	214	22	215
rect	21	217	22	218
rect	21	220	22	221
rect	21	223	22	224
rect	21	226	22	227
rect	21	229	22	230
rect	21	232	22	233
rect	21	235	22	236
rect	21	238	22	239
rect	21	241	22	242
rect	21	244	22	245
rect	21	247	22	248
rect	21	250	22	251
rect	21	253	22	254
rect	21	256	22	257
rect	21	259	22	260
rect	21	262	22	263
rect	21	265	22	266
rect	21	268	22	269
rect	21	271	22	272
rect	21	274	22	275
rect	21	277	22	278
rect	21	280	22	281
rect	21	283	22	284
rect	21	286	22	287
rect	21	289	22	290
rect	21	292	22	293
rect	21	295	22	296
rect	21	298	22	299
rect	21	301	22	302
rect	21	304	22	305
rect	21	307	22	308
rect	21	310	22	311
rect	21	313	22	314
rect	21	316	22	317
rect	21	319	22	320
rect	21	322	22	323
rect	21	325	22	326
rect	21	328	22	329
rect	21	331	22	332
rect	21	334	22	335
rect	21	337	22	338
rect	21	340	22	341
rect	21	343	22	344
rect	21	346	22	347
rect	21	349	22	350
rect	21	352	22	353
rect	21	355	22	356
rect	21	358	22	359
rect	21	361	22	362
rect	21	364	22	365
rect	21	367	22	368
rect	21	373	22	374
rect	21	376	22	377
rect	21	379	22	380
rect	21	385	22	386
rect	22	1	23	2
rect	22	4	23	5
rect	22	7	23	8
rect	22	10	23	11
rect	22	13	23	14
rect	22	16	23	17
rect	22	19	23	20
rect	22	22	23	23
rect	22	25	23	26
rect	22	28	23	29
rect	22	31	23	32
rect	22	34	23	35
rect	22	37	23	38
rect	22	40	23	41
rect	22	43	23	44
rect	22	46	23	47
rect	22	49	23	50
rect	22	52	23	53
rect	22	55	23	56
rect	22	58	23	59
rect	22	61	23	62
rect	22	64	23	65
rect	22	67	23	68
rect	22	70	23	71
rect	22	73	23	74
rect	22	76	23	77
rect	22	79	23	80
rect	22	82	23	83
rect	22	85	23	86
rect	22	88	23	89
rect	22	91	23	92
rect	22	94	23	95
rect	22	97	23	98
rect	22	100	23	101
rect	22	103	23	104
rect	22	106	23	107
rect	22	109	23	110
rect	22	112	23	113
rect	22	115	23	116
rect	22	118	23	119
rect	22	121	23	122
rect	22	124	23	125
rect	22	127	23	128
rect	22	130	23	131
rect	22	133	23	134
rect	22	136	23	137
rect	22	139	23	140
rect	22	142	23	143
rect	22	145	23	146
rect	22	148	23	149
rect	22	151	23	152
rect	22	154	23	155
rect	22	157	23	158
rect	22	160	23	161
rect	22	163	23	164
rect	22	166	23	167
rect	22	169	23	170
rect	22	172	23	173
rect	22	175	23	176
rect	22	178	23	179
rect	22	181	23	182
rect	22	184	23	185
rect	22	187	23	188
rect	22	190	23	191
rect	22	193	23	194
rect	22	196	23	197
rect	22	199	23	200
rect	22	202	23	203
rect	22	205	23	206
rect	22	208	23	209
rect	22	211	23	212
rect	22	214	23	215
rect	22	217	23	218
rect	22	220	23	221
rect	22	223	23	224
rect	22	226	23	227
rect	22	229	23	230
rect	22	232	23	233
rect	22	235	23	236
rect	22	238	23	239
rect	22	241	23	242
rect	22	244	23	245
rect	22	247	23	248
rect	22	250	23	251
rect	22	253	23	254
rect	22	256	23	257
rect	22	259	23	260
rect	22	262	23	263
rect	22	265	23	266
rect	22	268	23	269
rect	22	271	23	272
rect	22	274	23	275
rect	22	277	23	278
rect	22	280	23	281
rect	22	283	23	284
rect	22	286	23	287
rect	22	289	23	290
rect	22	292	23	293
rect	22	295	23	296
rect	22	298	23	299
rect	22	301	23	302
rect	22	304	23	305
rect	22	307	23	308
rect	22	310	23	311
rect	22	313	23	314
rect	22	316	23	317
rect	22	319	23	320
rect	22	322	23	323
rect	22	325	23	326
rect	22	328	23	329
rect	22	331	23	332
rect	22	334	23	335
rect	22	337	23	338
rect	22	340	23	341
rect	22	343	23	344
rect	22	346	23	347
rect	22	349	23	350
rect	22	352	23	353
rect	22	355	23	356
rect	22	358	23	359
rect	22	361	23	362
rect	22	364	23	365
rect	22	367	23	368
rect	22	373	23	374
rect	22	376	23	377
rect	22	379	23	380
rect	22	385	23	386
rect	23	1	24	2
rect	23	4	24	5
rect	23	7	24	8
rect	23	10	24	11
rect	23	13	24	14
rect	23	16	24	17
rect	23	19	24	20
rect	23	22	24	23
rect	23	25	24	26
rect	23	28	24	29
rect	23	31	24	32
rect	23	34	24	35
rect	23	37	24	38
rect	23	40	24	41
rect	23	43	24	44
rect	23	46	24	47
rect	23	49	24	50
rect	23	52	24	53
rect	23	55	24	56
rect	23	58	24	59
rect	23	61	24	62
rect	23	64	24	65
rect	23	67	24	68
rect	23	70	24	71
rect	23	73	24	74
rect	23	76	24	77
rect	23	79	24	80
rect	23	82	24	83
rect	23	85	24	86
rect	23	88	24	89
rect	23	91	24	92
rect	23	94	24	95
rect	23	97	24	98
rect	23	100	24	101
rect	23	103	24	104
rect	23	106	24	107
rect	23	109	24	110
rect	23	112	24	113
rect	23	115	24	116
rect	23	118	24	119
rect	23	121	24	122
rect	23	124	24	125
rect	23	127	24	128
rect	23	130	24	131
rect	23	133	24	134
rect	23	136	24	137
rect	23	139	24	140
rect	23	142	24	143
rect	23	145	24	146
rect	23	148	24	149
rect	23	151	24	152
rect	23	154	24	155
rect	23	157	24	158
rect	23	160	24	161
rect	23	163	24	164
rect	23	166	24	167
rect	23	169	24	170
rect	23	172	24	173
rect	23	175	24	176
rect	23	178	24	179
rect	23	181	24	182
rect	23	184	24	185
rect	23	187	24	188
rect	23	190	24	191
rect	23	193	24	194
rect	23	196	24	197
rect	23	199	24	200
rect	23	202	24	203
rect	23	205	24	206
rect	23	208	24	209
rect	23	211	24	212
rect	23	214	24	215
rect	23	217	24	218
rect	23	220	24	221
rect	23	223	24	224
rect	23	226	24	227
rect	23	229	24	230
rect	23	232	24	233
rect	23	235	24	236
rect	23	238	24	239
rect	23	241	24	242
rect	23	244	24	245
rect	23	247	24	248
rect	23	250	24	251
rect	23	253	24	254
rect	23	256	24	257
rect	23	259	24	260
rect	23	262	24	263
rect	23	265	24	266
rect	23	268	24	269
rect	23	271	24	272
rect	23	274	24	275
rect	23	277	24	278
rect	23	280	24	281
rect	23	283	24	284
rect	23	286	24	287
rect	23	289	24	290
rect	23	292	24	293
rect	23	295	24	296
rect	23	298	24	299
rect	23	301	24	302
rect	23	304	24	305
rect	23	307	24	308
rect	23	310	24	311
rect	23	313	24	314
rect	23	316	24	317
rect	23	319	24	320
rect	23	322	24	323
rect	23	325	24	326
rect	23	328	24	329
rect	23	331	24	332
rect	23	334	24	335
rect	23	337	24	338
rect	23	340	24	341
rect	23	343	24	344
rect	23	346	24	347
rect	23	349	24	350
rect	23	352	24	353
rect	23	355	24	356
rect	23	358	24	359
rect	23	361	24	362
rect	23	364	24	365
rect	23	367	24	368
rect	23	373	24	374
rect	23	376	24	377
rect	23	379	24	380
rect	23	385	24	386
rect	24	1	25	2
rect	24	4	25	5
rect	24	7	25	8
rect	24	10	25	11
rect	24	13	25	14
rect	24	16	25	17
rect	24	19	25	20
rect	24	22	25	23
rect	24	25	25	26
rect	24	28	25	29
rect	24	31	25	32
rect	24	34	25	35
rect	24	37	25	38
rect	24	40	25	41
rect	24	43	25	44
rect	24	46	25	47
rect	24	49	25	50
rect	24	52	25	53
rect	24	55	25	56
rect	24	58	25	59
rect	24	61	25	62
rect	24	64	25	65
rect	24	67	25	68
rect	24	70	25	71
rect	24	73	25	74
rect	24	76	25	77
rect	24	79	25	80
rect	24	82	25	83
rect	24	85	25	86
rect	24	88	25	89
rect	24	91	25	92
rect	24	94	25	95
rect	24	97	25	98
rect	24	100	25	101
rect	24	103	25	104
rect	24	106	25	107
rect	24	109	25	110
rect	24	112	25	113
rect	24	115	25	116
rect	24	118	25	119
rect	24	121	25	122
rect	24	124	25	125
rect	24	127	25	128
rect	24	130	25	131
rect	24	133	25	134
rect	24	136	25	137
rect	24	139	25	140
rect	24	142	25	143
rect	24	145	25	146
rect	24	148	25	149
rect	24	151	25	152
rect	24	154	25	155
rect	24	157	25	158
rect	24	160	25	161
rect	24	163	25	164
rect	24	166	25	167
rect	24	169	25	170
rect	24	172	25	173
rect	24	175	25	176
rect	24	178	25	179
rect	24	181	25	182
rect	24	184	25	185
rect	24	187	25	188
rect	24	190	25	191
rect	24	193	25	194
rect	24	196	25	197
rect	24	199	25	200
rect	24	202	25	203
rect	24	205	25	206
rect	24	208	25	209
rect	24	211	25	212
rect	24	214	25	215
rect	24	217	25	218
rect	24	220	25	221
rect	24	223	25	224
rect	24	226	25	227
rect	24	229	25	230
rect	24	232	25	233
rect	24	235	25	236
rect	24	238	25	239
rect	24	241	25	242
rect	24	244	25	245
rect	24	247	25	248
rect	24	250	25	251
rect	24	253	25	254
rect	24	256	25	257
rect	24	259	25	260
rect	24	262	25	263
rect	24	265	25	266
rect	24	268	25	269
rect	24	271	25	272
rect	24	274	25	275
rect	24	277	25	278
rect	24	280	25	281
rect	24	283	25	284
rect	24	286	25	287
rect	24	289	25	290
rect	24	292	25	293
rect	24	295	25	296
rect	24	298	25	299
rect	24	301	25	302
rect	24	304	25	305
rect	24	307	25	308
rect	24	310	25	311
rect	24	313	25	314
rect	24	316	25	317
rect	24	319	25	320
rect	24	322	25	323
rect	24	325	25	326
rect	24	328	25	329
rect	24	331	25	332
rect	24	334	25	335
rect	24	337	25	338
rect	24	340	25	341
rect	24	343	25	344
rect	24	346	25	347
rect	24	349	25	350
rect	24	352	25	353
rect	24	355	25	356
rect	24	358	25	359
rect	24	361	25	362
rect	24	364	25	365
rect	24	367	25	368
rect	24	373	25	374
rect	24	376	25	377
rect	24	379	25	380
rect	24	385	25	386
rect	25	1	26	2
rect	25	4	26	5
rect	25	7	26	8
rect	25	10	26	11
rect	25	13	26	14
rect	25	16	26	17
rect	25	19	26	20
rect	25	22	26	23
rect	25	25	26	26
rect	25	28	26	29
rect	25	31	26	32
rect	25	34	26	35
rect	25	37	26	38
rect	25	40	26	41
rect	25	43	26	44
rect	25	46	26	47
rect	25	49	26	50
rect	25	52	26	53
rect	25	55	26	56
rect	25	58	26	59
rect	25	61	26	62
rect	25	64	26	65
rect	25	67	26	68
rect	25	70	26	71
rect	25	73	26	74
rect	25	76	26	77
rect	25	79	26	80
rect	25	82	26	83
rect	25	85	26	86
rect	25	88	26	89
rect	25	91	26	92
rect	25	94	26	95
rect	25	97	26	98
rect	25	100	26	101
rect	25	103	26	104
rect	25	106	26	107
rect	25	109	26	110
rect	25	112	26	113
rect	25	115	26	116
rect	25	118	26	119
rect	25	121	26	122
rect	25	124	26	125
rect	25	127	26	128
rect	25	130	26	131
rect	25	133	26	134
rect	25	136	26	137
rect	25	139	26	140
rect	25	142	26	143
rect	25	145	26	146
rect	25	148	26	149
rect	25	151	26	152
rect	25	154	26	155
rect	25	157	26	158
rect	25	160	26	161
rect	25	163	26	164
rect	25	166	26	167
rect	25	169	26	170
rect	25	172	26	173
rect	25	175	26	176
rect	25	178	26	179
rect	25	181	26	182
rect	25	184	26	185
rect	25	187	26	188
rect	25	190	26	191
rect	25	193	26	194
rect	25	196	26	197
rect	25	199	26	200
rect	25	202	26	203
rect	25	205	26	206
rect	25	208	26	209
rect	25	211	26	212
rect	25	214	26	215
rect	25	217	26	218
rect	25	220	26	221
rect	25	223	26	224
rect	25	226	26	227
rect	25	229	26	230
rect	25	232	26	233
rect	25	235	26	236
rect	25	238	26	239
rect	25	241	26	242
rect	25	244	26	245
rect	25	247	26	248
rect	25	250	26	251
rect	25	253	26	254
rect	25	256	26	257
rect	25	259	26	260
rect	25	262	26	263
rect	25	265	26	266
rect	25	268	26	269
rect	25	271	26	272
rect	25	274	26	275
rect	25	277	26	278
rect	25	280	26	281
rect	25	283	26	284
rect	25	286	26	287
rect	25	289	26	290
rect	25	292	26	293
rect	25	295	26	296
rect	25	298	26	299
rect	25	301	26	302
rect	25	304	26	305
rect	25	307	26	308
rect	25	310	26	311
rect	25	313	26	314
rect	25	316	26	317
rect	25	319	26	320
rect	25	322	26	323
rect	25	325	26	326
rect	25	328	26	329
rect	25	331	26	332
rect	25	334	26	335
rect	25	337	26	338
rect	25	340	26	341
rect	25	343	26	344
rect	25	346	26	347
rect	25	349	26	350
rect	25	352	26	353
rect	25	355	26	356
rect	25	358	26	359
rect	25	361	26	362
rect	25	364	26	365
rect	25	367	26	368
rect	25	373	26	374
rect	25	376	26	377
rect	25	379	26	380
rect	25	385	26	386
rect	26	1	27	2
rect	26	4	27	5
rect	26	7	27	8
rect	26	10	27	11
rect	26	13	27	14
rect	26	16	27	17
rect	26	19	27	20
rect	26	22	27	23
rect	26	25	27	26
rect	26	28	27	29
rect	26	31	27	32
rect	26	34	27	35
rect	26	37	27	38
rect	26	40	27	41
rect	26	43	27	44
rect	26	46	27	47
rect	26	49	27	50
rect	26	52	27	53
rect	26	55	27	56
rect	26	58	27	59
rect	26	61	27	62
rect	26	64	27	65
rect	26	67	27	68
rect	26	70	27	71
rect	26	73	27	74
rect	26	76	27	77
rect	26	79	27	80
rect	26	82	27	83
rect	26	85	27	86
rect	26	88	27	89
rect	26	91	27	92
rect	26	94	27	95
rect	26	97	27	98
rect	26	100	27	101
rect	26	103	27	104
rect	26	106	27	107
rect	26	109	27	110
rect	26	112	27	113
rect	26	115	27	116
rect	26	118	27	119
rect	26	121	27	122
rect	26	124	27	125
rect	26	127	27	128
rect	26	130	27	131
rect	26	133	27	134
rect	26	136	27	137
rect	26	139	27	140
rect	26	142	27	143
rect	26	145	27	146
rect	26	148	27	149
rect	26	151	27	152
rect	26	154	27	155
rect	26	157	27	158
rect	26	160	27	161
rect	26	163	27	164
rect	26	166	27	167
rect	26	169	27	170
rect	26	172	27	173
rect	26	175	27	176
rect	26	178	27	179
rect	26	181	27	182
rect	26	184	27	185
rect	26	187	27	188
rect	26	190	27	191
rect	26	193	27	194
rect	26	196	27	197
rect	26	199	27	200
rect	26	202	27	203
rect	26	205	27	206
rect	26	208	27	209
rect	26	211	27	212
rect	26	214	27	215
rect	26	217	27	218
rect	26	220	27	221
rect	26	223	27	224
rect	26	226	27	227
rect	26	229	27	230
rect	26	232	27	233
rect	26	235	27	236
rect	26	238	27	239
rect	26	241	27	242
rect	26	244	27	245
rect	26	247	27	248
rect	26	250	27	251
rect	26	253	27	254
rect	26	256	27	257
rect	26	259	27	260
rect	26	262	27	263
rect	26	265	27	266
rect	26	268	27	269
rect	26	271	27	272
rect	26	274	27	275
rect	26	277	27	278
rect	26	280	27	281
rect	26	283	27	284
rect	26	286	27	287
rect	26	289	27	290
rect	26	292	27	293
rect	26	295	27	296
rect	26	298	27	299
rect	26	301	27	302
rect	26	304	27	305
rect	26	307	27	308
rect	26	310	27	311
rect	26	313	27	314
rect	26	316	27	317
rect	26	319	27	320
rect	26	322	27	323
rect	26	325	27	326
rect	26	328	27	329
rect	26	331	27	332
rect	26	334	27	335
rect	26	337	27	338
rect	26	340	27	341
rect	26	343	27	344
rect	26	346	27	347
rect	26	349	27	350
rect	26	352	27	353
rect	26	355	27	356
rect	26	358	27	359
rect	26	361	27	362
rect	26	364	27	365
rect	26	367	27	368
rect	26	373	27	374
rect	26	376	27	377
rect	26	379	27	380
rect	26	385	27	386
rect	27	1	28	2
rect	27	4	28	5
rect	27	7	28	8
rect	27	10	28	11
rect	27	13	28	14
rect	27	16	28	17
rect	27	19	28	20
rect	27	22	28	23
rect	27	25	28	26
rect	27	28	28	29
rect	27	31	28	32
rect	27	34	28	35
rect	27	37	28	38
rect	27	40	28	41
rect	27	43	28	44
rect	27	46	28	47
rect	27	49	28	50
rect	27	52	28	53
rect	27	55	28	56
rect	27	58	28	59
rect	27	61	28	62
rect	27	64	28	65
rect	27	67	28	68
rect	27	70	28	71
rect	27	73	28	74
rect	27	76	28	77
rect	27	79	28	80
rect	27	82	28	83
rect	27	85	28	86
rect	27	88	28	89
rect	27	91	28	92
rect	27	94	28	95
rect	27	97	28	98
rect	27	100	28	101
rect	27	103	28	104
rect	27	106	28	107
rect	27	109	28	110
rect	27	112	28	113
rect	27	115	28	116
rect	27	118	28	119
rect	27	121	28	122
rect	27	124	28	125
rect	27	127	28	128
rect	27	130	28	131
rect	27	133	28	134
rect	27	136	28	137
rect	27	139	28	140
rect	27	142	28	143
rect	27	145	28	146
rect	27	148	28	149
rect	27	151	28	152
rect	27	154	28	155
rect	27	157	28	158
rect	27	160	28	161
rect	27	163	28	164
rect	27	166	28	167
rect	27	169	28	170
rect	27	172	28	173
rect	27	175	28	176
rect	27	178	28	179
rect	27	181	28	182
rect	27	184	28	185
rect	27	187	28	188
rect	27	190	28	191
rect	27	193	28	194
rect	27	196	28	197
rect	27	199	28	200
rect	27	202	28	203
rect	27	205	28	206
rect	27	208	28	209
rect	27	211	28	212
rect	27	214	28	215
rect	27	217	28	218
rect	27	220	28	221
rect	27	223	28	224
rect	27	226	28	227
rect	27	229	28	230
rect	27	232	28	233
rect	27	235	28	236
rect	27	238	28	239
rect	27	241	28	242
rect	27	244	28	245
rect	27	247	28	248
rect	27	250	28	251
rect	27	253	28	254
rect	27	256	28	257
rect	27	259	28	260
rect	27	262	28	263
rect	27	265	28	266
rect	27	268	28	269
rect	27	271	28	272
rect	27	274	28	275
rect	27	277	28	278
rect	27	280	28	281
rect	27	283	28	284
rect	27	286	28	287
rect	27	289	28	290
rect	27	292	28	293
rect	27	295	28	296
rect	27	298	28	299
rect	27	301	28	302
rect	27	304	28	305
rect	27	307	28	308
rect	27	310	28	311
rect	27	313	28	314
rect	27	316	28	317
rect	27	319	28	320
rect	27	322	28	323
rect	27	325	28	326
rect	27	328	28	329
rect	27	331	28	332
rect	27	334	28	335
rect	27	337	28	338
rect	27	340	28	341
rect	27	343	28	344
rect	27	346	28	347
rect	27	349	28	350
rect	27	352	28	353
rect	27	355	28	356
rect	27	358	28	359
rect	27	361	28	362
rect	27	364	28	365
rect	27	367	28	368
rect	27	373	28	374
rect	27	376	28	377
rect	27	379	28	380
rect	27	385	28	386
rect	28	1	29	2
rect	28	4	29	5
rect	28	7	29	8
rect	28	10	29	11
rect	28	13	29	14
rect	28	16	29	17
rect	28	19	29	20
rect	28	22	29	23
rect	28	25	29	26
rect	28	28	29	29
rect	28	31	29	32
rect	28	34	29	35
rect	28	37	29	38
rect	28	40	29	41
rect	28	43	29	44
rect	28	46	29	47
rect	28	49	29	50
rect	28	52	29	53
rect	28	55	29	56
rect	28	58	29	59
rect	28	61	29	62
rect	28	64	29	65
rect	28	67	29	68
rect	28	70	29	71
rect	28	73	29	74
rect	28	76	29	77
rect	28	79	29	80
rect	28	82	29	83
rect	28	85	29	86
rect	28	88	29	89
rect	28	91	29	92
rect	28	94	29	95
rect	28	97	29	98
rect	28	100	29	101
rect	28	103	29	104
rect	28	106	29	107
rect	28	109	29	110
rect	28	112	29	113
rect	28	115	29	116
rect	28	118	29	119
rect	28	121	29	122
rect	28	124	29	125
rect	28	127	29	128
rect	28	130	29	131
rect	28	133	29	134
rect	28	136	29	137
rect	28	139	29	140
rect	28	142	29	143
rect	28	145	29	146
rect	28	148	29	149
rect	28	151	29	152
rect	28	154	29	155
rect	28	157	29	158
rect	28	160	29	161
rect	28	163	29	164
rect	28	166	29	167
rect	28	169	29	170
rect	28	172	29	173
rect	28	175	29	176
rect	28	178	29	179
rect	28	181	29	182
rect	28	184	29	185
rect	28	187	29	188
rect	28	190	29	191
rect	28	193	29	194
rect	28	196	29	197
rect	28	199	29	200
rect	28	202	29	203
rect	28	205	29	206
rect	28	208	29	209
rect	28	211	29	212
rect	28	214	29	215
rect	28	217	29	218
rect	28	220	29	221
rect	28	223	29	224
rect	28	226	29	227
rect	28	229	29	230
rect	28	232	29	233
rect	28	235	29	236
rect	28	238	29	239
rect	28	241	29	242
rect	28	244	29	245
rect	28	247	29	248
rect	28	250	29	251
rect	28	253	29	254
rect	28	256	29	257
rect	28	259	29	260
rect	28	262	29	263
rect	28	265	29	266
rect	28	268	29	269
rect	28	271	29	272
rect	28	274	29	275
rect	28	277	29	278
rect	28	280	29	281
rect	28	283	29	284
rect	28	286	29	287
rect	28	289	29	290
rect	28	292	29	293
rect	28	295	29	296
rect	28	298	29	299
rect	28	301	29	302
rect	28	304	29	305
rect	28	307	29	308
rect	28	310	29	311
rect	28	313	29	314
rect	28	316	29	317
rect	28	319	29	320
rect	28	322	29	323
rect	28	325	29	326
rect	28	328	29	329
rect	28	331	29	332
rect	28	334	29	335
rect	28	337	29	338
rect	28	340	29	341
rect	28	343	29	344
rect	28	346	29	347
rect	28	349	29	350
rect	28	352	29	353
rect	28	355	29	356
rect	28	358	29	359
rect	28	361	29	362
rect	28	364	29	365
rect	28	367	29	368
rect	28	373	29	374
rect	28	376	29	377
rect	28	379	29	380
rect	28	385	29	386
rect	29	1	30	2
rect	29	4	30	5
rect	29	7	30	8
rect	29	10	30	11
rect	29	13	30	14
rect	29	16	30	17
rect	29	19	30	20
rect	29	22	30	23
rect	29	25	30	26
rect	29	28	30	29
rect	29	31	30	32
rect	29	34	30	35
rect	29	37	30	38
rect	29	40	30	41
rect	29	43	30	44
rect	29	46	30	47
rect	29	49	30	50
rect	29	52	30	53
rect	29	55	30	56
rect	29	58	30	59
rect	29	61	30	62
rect	29	64	30	65
rect	29	67	30	68
rect	29	70	30	71
rect	29	73	30	74
rect	29	76	30	77
rect	29	79	30	80
rect	29	82	30	83
rect	29	85	30	86
rect	29	88	30	89
rect	29	91	30	92
rect	29	94	30	95
rect	29	97	30	98
rect	29	100	30	101
rect	29	103	30	104
rect	29	106	30	107
rect	29	109	30	110
rect	29	112	30	113
rect	29	115	30	116
rect	29	118	30	119
rect	29	121	30	122
rect	29	124	30	125
rect	29	127	30	128
rect	29	130	30	131
rect	29	133	30	134
rect	29	136	30	137
rect	29	139	30	140
rect	29	142	30	143
rect	29	145	30	146
rect	29	148	30	149
rect	29	151	30	152
rect	29	154	30	155
rect	29	157	30	158
rect	29	160	30	161
rect	29	163	30	164
rect	29	166	30	167
rect	29	169	30	170
rect	29	172	30	173
rect	29	175	30	176
rect	29	178	30	179
rect	29	181	30	182
rect	29	184	30	185
rect	29	187	30	188
rect	29	190	30	191
rect	29	193	30	194
rect	29	196	30	197
rect	29	199	30	200
rect	29	202	30	203
rect	29	205	30	206
rect	29	208	30	209
rect	29	211	30	212
rect	29	214	30	215
rect	29	217	30	218
rect	29	220	30	221
rect	29	223	30	224
rect	29	226	30	227
rect	29	229	30	230
rect	29	232	30	233
rect	29	235	30	236
rect	29	238	30	239
rect	29	241	30	242
rect	29	244	30	245
rect	29	247	30	248
rect	29	250	30	251
rect	29	253	30	254
rect	29	256	30	257
rect	29	259	30	260
rect	29	262	30	263
rect	29	265	30	266
rect	29	268	30	269
rect	29	271	30	272
rect	29	274	30	275
rect	29	277	30	278
rect	29	280	30	281
rect	29	283	30	284
rect	29	286	30	287
rect	29	289	30	290
rect	29	292	30	293
rect	29	295	30	296
rect	29	298	30	299
rect	29	301	30	302
rect	29	304	30	305
rect	29	307	30	308
rect	29	310	30	311
rect	29	313	30	314
rect	29	316	30	317
rect	29	319	30	320
rect	29	322	30	323
rect	29	325	30	326
rect	29	328	30	329
rect	29	331	30	332
rect	29	334	30	335
rect	29	337	30	338
rect	29	340	30	341
rect	29	343	30	344
rect	29	346	30	347
rect	29	349	30	350
rect	29	352	30	353
rect	29	355	30	356
rect	29	358	30	359
rect	29	361	30	362
rect	29	364	30	365
rect	29	367	30	368
rect	29	373	30	374
rect	29	376	30	377
rect	29	379	30	380
rect	29	385	30	386
rect	30	1	31	2
rect	30	4	31	5
rect	30	7	31	8
rect	30	10	31	11
rect	30	13	31	14
rect	30	16	31	17
rect	30	19	31	20
rect	30	22	31	23
rect	30	25	31	26
rect	30	28	31	29
rect	30	31	31	32
rect	30	34	31	35
rect	30	37	31	38
rect	30	40	31	41
rect	30	43	31	44
rect	30	46	31	47
rect	30	49	31	50
rect	30	52	31	53
rect	30	55	31	56
rect	30	58	31	59
rect	30	61	31	62
rect	30	64	31	65
rect	30	67	31	68
rect	30	70	31	71
rect	30	73	31	74
rect	30	76	31	77
rect	30	79	31	80
rect	30	82	31	83
rect	30	85	31	86
rect	30	88	31	89
rect	30	91	31	92
rect	30	94	31	95
rect	30	97	31	98
rect	30	100	31	101
rect	30	103	31	104
rect	30	106	31	107
rect	30	109	31	110
rect	30	112	31	113
rect	30	115	31	116
rect	30	118	31	119
rect	30	121	31	122
rect	30	124	31	125
rect	30	127	31	128
rect	30	130	31	131
rect	30	133	31	134
rect	30	136	31	137
rect	30	139	31	140
rect	30	142	31	143
rect	30	145	31	146
rect	30	148	31	149
rect	30	151	31	152
rect	30	154	31	155
rect	30	157	31	158
rect	30	160	31	161
rect	30	163	31	164
rect	30	166	31	167
rect	30	169	31	170
rect	30	172	31	173
rect	30	175	31	176
rect	30	178	31	179
rect	30	181	31	182
rect	30	184	31	185
rect	30	187	31	188
rect	30	190	31	191
rect	30	193	31	194
rect	30	196	31	197
rect	30	199	31	200
rect	30	202	31	203
rect	30	205	31	206
rect	30	208	31	209
rect	30	211	31	212
rect	30	214	31	215
rect	30	217	31	218
rect	30	220	31	221
rect	30	223	31	224
rect	30	226	31	227
rect	30	229	31	230
rect	30	232	31	233
rect	30	235	31	236
rect	30	238	31	239
rect	30	241	31	242
rect	30	244	31	245
rect	30	247	31	248
rect	30	250	31	251
rect	30	253	31	254
rect	30	256	31	257
rect	30	259	31	260
rect	30	262	31	263
rect	30	265	31	266
rect	30	268	31	269
rect	30	271	31	272
rect	30	274	31	275
rect	30	277	31	278
rect	30	280	31	281
rect	30	283	31	284
rect	30	286	31	287
rect	30	289	31	290
rect	30	292	31	293
rect	30	295	31	296
rect	30	298	31	299
rect	30	301	31	302
rect	30	304	31	305
rect	30	307	31	308
rect	30	310	31	311
rect	30	313	31	314
rect	30	316	31	317
rect	30	319	31	320
rect	30	322	31	323
rect	30	325	31	326
rect	30	328	31	329
rect	30	331	31	332
rect	30	334	31	335
rect	30	337	31	338
rect	30	340	31	341
rect	30	343	31	344
rect	30	346	31	347
rect	30	349	31	350
rect	30	352	31	353
rect	30	355	31	356
rect	30	358	31	359
rect	30	361	31	362
rect	30	364	31	365
rect	30	367	31	368
rect	30	373	31	374
rect	30	376	31	377
rect	30	379	31	380
rect	30	385	31	386
rect	31	1	32	2
rect	31	4	32	5
rect	31	7	32	8
rect	31	10	32	11
rect	31	13	32	14
rect	31	16	32	17
rect	31	19	32	20
rect	31	22	32	23
rect	31	25	32	26
rect	31	28	32	29
rect	31	31	32	32
rect	31	34	32	35
rect	31	37	32	38
rect	31	40	32	41
rect	31	43	32	44
rect	31	46	32	47
rect	31	49	32	50
rect	31	52	32	53
rect	31	55	32	56
rect	31	58	32	59
rect	31	61	32	62
rect	31	64	32	65
rect	31	67	32	68
rect	31	70	32	71
rect	31	73	32	74
rect	31	76	32	77
rect	31	79	32	80
rect	31	82	32	83
rect	31	85	32	86
rect	31	88	32	89
rect	31	91	32	92
rect	31	94	32	95
rect	31	97	32	98
rect	31	100	32	101
rect	31	103	32	104
rect	31	106	32	107
rect	31	109	32	110
rect	31	112	32	113
rect	31	115	32	116
rect	31	118	32	119
rect	31	121	32	122
rect	31	124	32	125
rect	31	127	32	128
rect	31	130	32	131
rect	31	133	32	134
rect	31	136	32	137
rect	31	139	32	140
rect	31	142	32	143
rect	31	145	32	146
rect	31	148	32	149
rect	31	151	32	152
rect	31	154	32	155
rect	31	157	32	158
rect	31	160	32	161
rect	31	163	32	164
rect	31	166	32	167
rect	31	169	32	170
rect	31	172	32	173
rect	31	175	32	176
rect	31	178	32	179
rect	31	181	32	182
rect	31	184	32	185
rect	31	187	32	188
rect	31	190	32	191
rect	31	193	32	194
rect	31	196	32	197
rect	31	199	32	200
rect	31	202	32	203
rect	31	205	32	206
rect	31	208	32	209
rect	31	211	32	212
rect	31	214	32	215
rect	31	217	32	218
rect	31	220	32	221
rect	31	223	32	224
rect	31	226	32	227
rect	31	229	32	230
rect	31	232	32	233
rect	31	235	32	236
rect	31	238	32	239
rect	31	241	32	242
rect	31	244	32	245
rect	31	247	32	248
rect	31	250	32	251
rect	31	253	32	254
rect	31	256	32	257
rect	31	259	32	260
rect	31	262	32	263
rect	31	265	32	266
rect	31	268	32	269
rect	31	271	32	272
rect	31	274	32	275
rect	31	277	32	278
rect	31	280	32	281
rect	31	283	32	284
rect	31	286	32	287
rect	31	289	32	290
rect	31	292	32	293
rect	31	295	32	296
rect	31	298	32	299
rect	31	301	32	302
rect	31	304	32	305
rect	31	307	32	308
rect	31	310	32	311
rect	31	313	32	314
rect	31	316	32	317
rect	31	319	32	320
rect	31	322	32	323
rect	31	325	32	326
rect	31	328	32	329
rect	31	331	32	332
rect	31	334	32	335
rect	31	337	32	338
rect	31	340	32	341
rect	31	343	32	344
rect	31	346	32	347
rect	31	349	32	350
rect	31	352	32	353
rect	31	355	32	356
rect	31	358	32	359
rect	31	361	32	362
rect	31	364	32	365
rect	31	367	32	368
rect	31	373	32	374
rect	31	376	32	377
rect	31	379	32	380
rect	31	385	32	386
rect	32	1	33	2
rect	32	4	33	5
rect	32	7	33	8
rect	32	10	33	11
rect	32	13	33	14
rect	32	16	33	17
rect	32	19	33	20
rect	32	22	33	23
rect	32	25	33	26
rect	32	28	33	29
rect	32	31	33	32
rect	32	34	33	35
rect	32	37	33	38
rect	32	40	33	41
rect	32	43	33	44
rect	32	46	33	47
rect	32	49	33	50
rect	32	52	33	53
rect	32	55	33	56
rect	32	58	33	59
rect	32	61	33	62
rect	32	64	33	65
rect	32	67	33	68
rect	32	70	33	71
rect	32	73	33	74
rect	32	76	33	77
rect	32	79	33	80
rect	32	82	33	83
rect	32	85	33	86
rect	32	88	33	89
rect	32	91	33	92
rect	32	94	33	95
rect	32	97	33	98
rect	32	100	33	101
rect	32	103	33	104
rect	32	106	33	107
rect	32	109	33	110
rect	32	112	33	113
rect	32	115	33	116
rect	32	118	33	119
rect	32	121	33	122
rect	32	124	33	125
rect	32	127	33	128
rect	32	130	33	131
rect	32	133	33	134
rect	32	136	33	137
rect	32	139	33	140
rect	32	142	33	143
rect	32	145	33	146
rect	32	148	33	149
rect	32	151	33	152
rect	32	154	33	155
rect	32	157	33	158
rect	32	160	33	161
rect	32	163	33	164
rect	32	166	33	167
rect	32	169	33	170
rect	32	172	33	173
rect	32	175	33	176
rect	32	178	33	179
rect	32	181	33	182
rect	32	184	33	185
rect	32	187	33	188
rect	32	190	33	191
rect	32	193	33	194
rect	32	196	33	197
rect	32	199	33	200
rect	32	202	33	203
rect	32	205	33	206
rect	32	208	33	209
rect	32	211	33	212
rect	32	214	33	215
rect	32	217	33	218
rect	32	220	33	221
rect	32	223	33	224
rect	32	226	33	227
rect	32	229	33	230
rect	32	232	33	233
rect	32	235	33	236
rect	32	238	33	239
rect	32	241	33	242
rect	32	244	33	245
rect	32	247	33	248
rect	32	250	33	251
rect	32	253	33	254
rect	32	256	33	257
rect	32	259	33	260
rect	32	262	33	263
rect	32	265	33	266
rect	32	268	33	269
rect	32	271	33	272
rect	32	274	33	275
rect	32	277	33	278
rect	32	280	33	281
rect	32	283	33	284
rect	32	286	33	287
rect	32	289	33	290
rect	32	292	33	293
rect	32	295	33	296
rect	32	298	33	299
rect	32	301	33	302
rect	32	304	33	305
rect	32	307	33	308
rect	32	310	33	311
rect	32	313	33	314
rect	32	316	33	317
rect	32	319	33	320
rect	32	322	33	323
rect	32	325	33	326
rect	32	328	33	329
rect	32	331	33	332
rect	32	334	33	335
rect	32	337	33	338
rect	32	340	33	341
rect	32	343	33	344
rect	32	346	33	347
rect	32	349	33	350
rect	32	352	33	353
rect	32	355	33	356
rect	32	358	33	359
rect	32	361	33	362
rect	32	364	33	365
rect	32	367	33	368
rect	32	373	33	374
rect	32	376	33	377
rect	32	379	33	380
rect	32	385	33	386
rect	33	1	34	2
rect	33	4	34	5
rect	33	7	34	8
rect	33	10	34	11
rect	33	13	34	14
rect	33	16	34	17
rect	33	19	34	20
rect	33	22	34	23
rect	33	25	34	26
rect	33	28	34	29
rect	33	31	34	32
rect	33	34	34	35
rect	33	37	34	38
rect	33	40	34	41
rect	33	43	34	44
rect	33	46	34	47
rect	33	49	34	50
rect	33	52	34	53
rect	33	55	34	56
rect	33	58	34	59
rect	33	61	34	62
rect	33	64	34	65
rect	33	67	34	68
rect	33	70	34	71
rect	33	73	34	74
rect	33	76	34	77
rect	33	79	34	80
rect	33	82	34	83
rect	33	85	34	86
rect	33	88	34	89
rect	33	91	34	92
rect	33	94	34	95
rect	33	97	34	98
rect	33	100	34	101
rect	33	103	34	104
rect	33	106	34	107
rect	33	109	34	110
rect	33	112	34	113
rect	33	115	34	116
rect	33	118	34	119
rect	33	121	34	122
rect	33	124	34	125
rect	33	127	34	128
rect	33	130	34	131
rect	33	133	34	134
rect	33	136	34	137
rect	33	139	34	140
rect	33	142	34	143
rect	33	145	34	146
rect	33	148	34	149
rect	33	151	34	152
rect	33	154	34	155
rect	33	157	34	158
rect	33	160	34	161
rect	33	163	34	164
rect	33	166	34	167
rect	33	169	34	170
rect	33	172	34	173
rect	33	175	34	176
rect	33	178	34	179
rect	33	181	34	182
rect	33	184	34	185
rect	33	187	34	188
rect	33	190	34	191
rect	33	193	34	194
rect	33	196	34	197
rect	33	199	34	200
rect	33	202	34	203
rect	33	205	34	206
rect	33	208	34	209
rect	33	211	34	212
rect	33	214	34	215
rect	33	217	34	218
rect	33	220	34	221
rect	33	223	34	224
rect	33	226	34	227
rect	33	229	34	230
rect	33	232	34	233
rect	33	235	34	236
rect	33	238	34	239
rect	33	241	34	242
rect	33	244	34	245
rect	33	247	34	248
rect	33	250	34	251
rect	33	253	34	254
rect	33	256	34	257
rect	33	259	34	260
rect	33	262	34	263
rect	33	265	34	266
rect	33	268	34	269
rect	33	271	34	272
rect	33	274	34	275
rect	33	277	34	278
rect	33	280	34	281
rect	33	283	34	284
rect	33	286	34	287
rect	33	289	34	290
rect	33	292	34	293
rect	33	295	34	296
rect	33	298	34	299
rect	33	301	34	302
rect	33	304	34	305
rect	33	307	34	308
rect	33	310	34	311
rect	33	313	34	314
rect	33	316	34	317
rect	33	319	34	320
rect	33	322	34	323
rect	33	325	34	326
rect	33	328	34	329
rect	33	331	34	332
rect	33	334	34	335
rect	33	337	34	338
rect	33	340	34	341
rect	33	343	34	344
rect	33	346	34	347
rect	33	349	34	350
rect	33	352	34	353
rect	33	355	34	356
rect	33	358	34	359
rect	33	361	34	362
rect	33	364	34	365
rect	33	367	34	368
rect	33	373	34	374
rect	33	376	34	377
rect	33	379	34	380
rect	33	385	34	386
rect	34	1	35	2
rect	34	4	35	5
rect	34	7	35	8
rect	34	10	35	11
rect	34	13	35	14
rect	34	16	35	17
rect	34	19	35	20
rect	34	22	35	23
rect	34	25	35	26
rect	34	28	35	29
rect	34	31	35	32
rect	34	34	35	35
rect	34	37	35	38
rect	34	40	35	41
rect	34	43	35	44
rect	34	46	35	47
rect	34	49	35	50
rect	34	52	35	53
rect	34	55	35	56
rect	34	58	35	59
rect	34	61	35	62
rect	34	64	35	65
rect	34	67	35	68
rect	34	70	35	71
rect	34	73	35	74
rect	34	76	35	77
rect	34	79	35	80
rect	34	82	35	83
rect	34	85	35	86
rect	34	88	35	89
rect	34	91	35	92
rect	34	94	35	95
rect	34	97	35	98
rect	34	100	35	101
rect	34	103	35	104
rect	34	106	35	107
rect	34	109	35	110
rect	34	112	35	113
rect	34	115	35	116
rect	34	118	35	119
rect	34	121	35	122
rect	34	124	35	125
rect	34	127	35	128
rect	34	130	35	131
rect	34	133	35	134
rect	34	136	35	137
rect	34	139	35	140
rect	34	142	35	143
rect	34	145	35	146
rect	34	148	35	149
rect	34	151	35	152
rect	34	154	35	155
rect	34	157	35	158
rect	34	160	35	161
rect	34	163	35	164
rect	34	166	35	167
rect	34	169	35	170
rect	34	172	35	173
rect	34	175	35	176
rect	34	178	35	179
rect	34	181	35	182
rect	34	184	35	185
rect	34	187	35	188
rect	34	190	35	191
rect	34	193	35	194
rect	34	196	35	197
rect	34	199	35	200
rect	34	202	35	203
rect	34	205	35	206
rect	34	208	35	209
rect	34	211	35	212
rect	34	214	35	215
rect	34	217	35	218
rect	34	220	35	221
rect	34	223	35	224
rect	34	226	35	227
rect	34	229	35	230
rect	34	232	35	233
rect	34	235	35	236
rect	34	238	35	239
rect	34	241	35	242
rect	34	244	35	245
rect	34	247	35	248
rect	34	250	35	251
rect	34	253	35	254
rect	34	256	35	257
rect	34	259	35	260
rect	34	262	35	263
rect	34	265	35	266
rect	34	268	35	269
rect	34	271	35	272
rect	34	274	35	275
rect	34	277	35	278
rect	34	280	35	281
rect	34	283	35	284
rect	34	286	35	287
rect	34	289	35	290
rect	34	292	35	293
rect	34	295	35	296
rect	34	298	35	299
rect	34	301	35	302
rect	34	304	35	305
rect	34	307	35	308
rect	34	310	35	311
rect	34	313	35	314
rect	34	316	35	317
rect	34	319	35	320
rect	34	322	35	323
rect	34	325	35	326
rect	34	328	35	329
rect	34	331	35	332
rect	34	334	35	335
rect	34	337	35	338
rect	34	340	35	341
rect	34	343	35	344
rect	34	346	35	347
rect	34	349	35	350
rect	34	352	35	353
rect	34	355	35	356
rect	34	358	35	359
rect	34	361	35	362
rect	34	364	35	365
rect	34	367	35	368
rect	34	373	35	374
rect	34	376	35	377
rect	34	379	35	380
rect	34	385	35	386
rect	35	1	36	2
rect	35	4	36	5
rect	35	7	36	8
rect	35	13	36	14
rect	35	16	36	17
rect	35	19	36	20
rect	35	22	36	23
rect	35	25	36	26
rect	35	28	36	29
rect	35	31	36	32
rect	35	34	36	35
rect	35	37	36	38
rect	35	40	36	41
rect	35	43	36	44
rect	35	46	36	47
rect	35	49	36	50
rect	35	52	36	53
rect	35	55	36	56
rect	35	58	36	59
rect	35	61	36	62
rect	35	64	36	65
rect	35	67	36	68
rect	35	70	36	71
rect	35	73	36	74
rect	35	76	36	77
rect	35	79	36	80
rect	35	82	36	83
rect	35	85	36	86
rect	35	88	36	89
rect	35	91	36	92
rect	35	94	36	95
rect	35	97	36	98
rect	35	100	36	101
rect	35	103	36	104
rect	35	106	36	107
rect	35	109	36	110
rect	35	112	36	113
rect	35	115	36	116
rect	35	118	36	119
rect	35	121	36	122
rect	35	124	36	125
rect	35	127	36	128
rect	35	130	36	131
rect	35	133	36	134
rect	35	136	36	137
rect	35	139	36	140
rect	35	142	36	143
rect	35	145	36	146
rect	35	148	36	149
rect	35	151	36	152
rect	35	154	36	155
rect	35	157	36	158
rect	35	160	36	161
rect	35	163	36	164
rect	35	166	36	167
rect	35	169	36	170
rect	35	172	36	173
rect	35	175	36	176
rect	35	178	36	179
rect	35	181	36	182
rect	35	184	36	185
rect	35	187	36	188
rect	35	190	36	191
rect	35	193	36	194
rect	35	196	36	197
rect	35	199	36	200
rect	35	202	36	203
rect	35	205	36	206
rect	35	208	36	209
rect	35	211	36	212
rect	35	214	36	215
rect	35	217	36	218
rect	35	220	36	221
rect	35	223	36	224
rect	35	226	36	227
rect	35	229	36	230
rect	35	232	36	233
rect	35	235	36	236
rect	35	238	36	239
rect	35	241	36	242
rect	35	244	36	245
rect	35	247	36	248
rect	35	250	36	251
rect	35	253	36	254
rect	35	256	36	257
rect	35	259	36	260
rect	35	262	36	263
rect	35	265	36	266
rect	35	268	36	269
rect	35	271	36	272
rect	35	274	36	275
rect	35	277	36	278
rect	35	280	36	281
rect	35	283	36	284
rect	35	286	36	287
rect	35	289	36	290
rect	35	292	36	293
rect	35	295	36	296
rect	35	298	36	299
rect	35	301	36	302
rect	35	304	36	305
rect	35	307	36	308
rect	35	310	36	311
rect	35	313	36	314
rect	35	316	36	317
rect	35	319	36	320
rect	35	322	36	323
rect	35	325	36	326
rect	35	328	36	329
rect	35	331	36	332
rect	35	334	36	335
rect	35	337	36	338
rect	35	340	36	341
rect	35	343	36	344
rect	35	346	36	347
rect	35	349	36	350
rect	35	352	36	353
rect	35	355	36	356
rect	35	358	36	359
rect	35	361	36	362
rect	35	364	36	365
rect	35	367	36	368
rect	35	373	36	374
rect	35	376	36	377
rect	35	379	36	380
rect	35	385	36	386
rect	36	1	37	2
rect	36	4	37	5
rect	36	7	37	8
rect	36	10	37	11
rect	36	13	37	14
rect	36	16	37	17
rect	36	19	37	20
rect	36	22	37	23
rect	36	25	37	26
rect	36	28	37	29
rect	36	31	37	32
rect	36	34	37	35
rect	36	37	37	38
rect	36	40	37	41
rect	36	43	37	44
rect	36	46	37	47
rect	36	49	37	50
rect	36	52	37	53
rect	36	55	37	56
rect	36	58	37	59
rect	36	61	37	62
rect	36	64	37	65
rect	36	67	37	68
rect	36	70	37	71
rect	36	73	37	74
rect	36	76	37	77
rect	36	79	37	80
rect	36	82	37	83
rect	36	85	37	86
rect	36	88	37	89
rect	36	91	37	92
rect	36	94	37	95
rect	36	97	37	98
rect	36	100	37	101
rect	36	103	37	104
rect	36	106	37	107
rect	36	109	37	110
rect	36	112	37	113
rect	36	115	37	116
rect	36	118	37	119
rect	36	121	37	122
rect	36	124	37	125
rect	36	127	37	128
rect	36	130	37	131
rect	36	133	37	134
rect	36	136	37	137
rect	36	139	37	140
rect	36	142	37	143
rect	36	145	37	146
rect	36	148	37	149
rect	36	151	37	152
rect	36	154	37	155
rect	36	157	37	158
rect	36	160	37	161
rect	36	163	37	164
rect	36	166	37	167
rect	36	169	37	170
rect	36	172	37	173
rect	36	175	37	176
rect	36	178	37	179
rect	36	181	37	182
rect	36	184	37	185
rect	36	187	37	188
rect	36	190	37	191
rect	36	193	37	194
rect	36	196	37	197
rect	36	199	37	200
rect	36	202	37	203
rect	36	205	37	206
rect	36	208	37	209
rect	36	211	37	212
rect	36	214	37	215
rect	36	217	37	218
rect	36	220	37	221
rect	36	223	37	224
rect	36	226	37	227
rect	36	229	37	230
rect	36	232	37	233
rect	36	235	37	236
rect	36	238	37	239
rect	36	241	37	242
rect	36	244	37	245
rect	36	247	37	248
rect	36	250	37	251
rect	36	253	37	254
rect	36	256	37	257
rect	36	259	37	260
rect	36	262	37	263
rect	36	265	37	266
rect	36	268	37	269
rect	36	271	37	272
rect	36	274	37	275
rect	36	277	37	278
rect	36	280	37	281
rect	36	283	37	284
rect	36	286	37	287
rect	36	289	37	290
rect	36	292	37	293
rect	36	295	37	296
rect	36	298	37	299
rect	36	301	37	302
rect	36	304	37	305
rect	36	307	37	308
rect	36	310	37	311
rect	36	313	37	314
rect	36	316	37	317
rect	36	319	37	320
rect	36	322	37	323
rect	36	325	37	326
rect	36	328	37	329
rect	36	331	37	332
rect	36	334	37	335
rect	36	337	37	338
rect	36	340	37	341
rect	36	343	37	344
rect	36	346	37	347
rect	36	349	37	350
rect	36	352	37	353
rect	36	355	37	356
rect	36	358	37	359
rect	36	361	37	362
rect	36	364	37	365
rect	36	367	37	368
rect	36	373	37	374
rect	36	376	37	377
rect	36	379	37	380
rect	36	385	37	386
rect	37	1	38	2
rect	37	4	38	5
rect	37	7	38	8
rect	37	10	38	11
rect	37	13	38	14
rect	37	16	38	17
rect	37	19	38	20
rect	37	22	38	23
rect	37	25	38	26
rect	37	28	38	29
rect	37	31	38	32
rect	37	34	38	35
rect	37	37	38	38
rect	37	40	38	41
rect	37	43	38	44
rect	37	46	38	47
rect	37	49	38	50
rect	37	52	38	53
rect	37	55	38	56
rect	37	58	38	59
rect	37	61	38	62
rect	37	64	38	65
rect	37	67	38	68
rect	37	70	38	71
rect	37	73	38	74
rect	37	76	38	77
rect	37	79	38	80
rect	37	82	38	83
rect	37	85	38	86
rect	37	88	38	89
rect	37	91	38	92
rect	37	94	38	95
rect	37	97	38	98
rect	37	100	38	101
rect	37	103	38	104
rect	37	106	38	107
rect	37	109	38	110
rect	37	112	38	113
rect	37	115	38	116
rect	37	118	38	119
rect	37	121	38	122
rect	37	124	38	125
rect	37	127	38	128
rect	37	130	38	131
rect	37	133	38	134
rect	37	136	38	137
rect	37	139	38	140
rect	37	142	38	143
rect	37	145	38	146
rect	37	148	38	149
rect	37	151	38	152
rect	37	154	38	155
rect	37	157	38	158
rect	37	160	38	161
rect	37	163	38	164
rect	37	166	38	167
rect	37	169	38	170
rect	37	172	38	173
rect	37	175	38	176
rect	37	178	38	179
rect	37	181	38	182
rect	37	184	38	185
rect	37	187	38	188
rect	37	190	38	191
rect	37	193	38	194
rect	37	196	38	197
rect	37	199	38	200
rect	37	202	38	203
rect	37	205	38	206
rect	37	208	38	209
rect	37	211	38	212
rect	37	214	38	215
rect	37	217	38	218
rect	37	220	38	221
rect	37	223	38	224
rect	37	226	38	227
rect	37	229	38	230
rect	37	232	38	233
rect	37	235	38	236
rect	37	238	38	239
rect	37	241	38	242
rect	37	244	38	245
rect	37	247	38	248
rect	37	250	38	251
rect	37	253	38	254
rect	37	256	38	257
rect	37	259	38	260
rect	37	262	38	263
rect	37	265	38	266
rect	37	268	38	269
rect	37	271	38	272
rect	37	274	38	275
rect	37	277	38	278
rect	37	280	38	281
rect	37	283	38	284
rect	37	286	38	287
rect	37	289	38	290
rect	37	292	38	293
rect	37	295	38	296
rect	37	298	38	299
rect	37	301	38	302
rect	37	304	38	305
rect	37	307	38	308
rect	37	310	38	311
rect	37	313	38	314
rect	37	316	38	317
rect	37	319	38	320
rect	37	322	38	323
rect	37	325	38	326
rect	37	328	38	329
rect	37	331	38	332
rect	37	334	38	335
rect	37	337	38	338
rect	37	340	38	341
rect	37	343	38	344
rect	37	346	38	347
rect	37	349	38	350
rect	37	352	38	353
rect	37	355	38	356
rect	37	358	38	359
rect	37	361	38	362
rect	37	364	38	365
rect	37	367	38	368
rect	37	373	38	374
rect	37	376	38	377
rect	37	379	38	380
rect	37	385	38	386
rect	38	1	39	2
rect	38	4	39	5
rect	38	7	39	8
rect	38	10	39	11
rect	38	13	39	14
rect	38	16	39	17
rect	38	19	39	20
rect	38	22	39	23
rect	38	25	39	26
rect	38	28	39	29
rect	38	31	39	32
rect	38	34	39	35
rect	38	37	39	38
rect	38	40	39	41
rect	38	43	39	44
rect	38	46	39	47
rect	38	49	39	50
rect	38	52	39	53
rect	38	55	39	56
rect	38	58	39	59
rect	38	61	39	62
rect	38	64	39	65
rect	38	67	39	68
rect	38	70	39	71
rect	38	73	39	74
rect	38	76	39	77
rect	38	79	39	80
rect	38	82	39	83
rect	38	85	39	86
rect	38	88	39	89
rect	38	91	39	92
rect	38	94	39	95
rect	38	97	39	98
rect	38	100	39	101
rect	38	103	39	104
rect	38	106	39	107
rect	38	109	39	110
rect	38	112	39	113
rect	38	115	39	116
rect	38	118	39	119
rect	38	121	39	122
rect	38	124	39	125
rect	38	127	39	128
rect	38	130	39	131
rect	38	133	39	134
rect	38	136	39	137
rect	38	139	39	140
rect	38	142	39	143
rect	38	145	39	146
rect	38	148	39	149
rect	38	151	39	152
rect	38	154	39	155
rect	38	157	39	158
rect	38	160	39	161
rect	38	163	39	164
rect	38	166	39	167
rect	38	169	39	170
rect	38	172	39	173
rect	38	175	39	176
rect	38	178	39	179
rect	38	181	39	182
rect	38	184	39	185
rect	38	187	39	188
rect	38	190	39	191
rect	38	193	39	194
rect	38	196	39	197
rect	38	199	39	200
rect	38	202	39	203
rect	38	205	39	206
rect	38	208	39	209
rect	38	211	39	212
rect	38	214	39	215
rect	38	217	39	218
rect	38	220	39	221
rect	38	223	39	224
rect	38	226	39	227
rect	38	229	39	230
rect	38	232	39	233
rect	38	235	39	236
rect	38	238	39	239
rect	38	241	39	242
rect	38	244	39	245
rect	38	247	39	248
rect	38	250	39	251
rect	38	253	39	254
rect	38	256	39	257
rect	38	259	39	260
rect	38	262	39	263
rect	38	265	39	266
rect	38	268	39	269
rect	38	271	39	272
rect	38	274	39	275
rect	38	277	39	278
rect	38	280	39	281
rect	38	283	39	284
rect	38	286	39	287
rect	38	289	39	290
rect	38	292	39	293
rect	38	295	39	296
rect	38	298	39	299
rect	38	301	39	302
rect	38	304	39	305
rect	38	307	39	308
rect	38	310	39	311
rect	38	313	39	314
rect	38	316	39	317
rect	38	319	39	320
rect	38	322	39	323
rect	38	325	39	326
rect	38	328	39	329
rect	38	331	39	332
rect	38	334	39	335
rect	38	337	39	338
rect	38	340	39	341
rect	38	343	39	344
rect	38	346	39	347
rect	38	349	39	350
rect	38	352	39	353
rect	38	355	39	356
rect	38	358	39	359
rect	38	361	39	362
rect	38	364	39	365
rect	38	367	39	368
rect	38	373	39	374
rect	38	376	39	377
rect	38	379	39	380
rect	38	385	39	386
rect	39	1	40	2
rect	39	4	40	5
rect	39	7	40	8
rect	39	10	40	11
rect	39	13	40	14
rect	39	16	40	17
rect	39	19	40	20
rect	39	22	40	23
rect	39	25	40	26
rect	39	28	40	29
rect	39	31	40	32
rect	39	34	40	35
rect	39	37	40	38
rect	39	40	40	41
rect	39	43	40	44
rect	39	46	40	47
rect	39	49	40	50
rect	39	52	40	53
rect	39	55	40	56
rect	39	58	40	59
rect	39	61	40	62
rect	39	64	40	65
rect	39	67	40	68
rect	39	70	40	71
rect	39	73	40	74
rect	39	76	40	77
rect	39	79	40	80
rect	39	82	40	83
rect	39	85	40	86
rect	39	88	40	89
rect	39	91	40	92
rect	39	94	40	95
rect	39	97	40	98
rect	39	100	40	101
rect	39	103	40	104
rect	39	106	40	107
rect	39	109	40	110
rect	39	112	40	113
rect	39	115	40	116
rect	39	118	40	119
rect	39	121	40	122
rect	39	124	40	125
rect	39	127	40	128
rect	39	130	40	131
rect	39	133	40	134
rect	39	136	40	137
rect	39	139	40	140
rect	39	142	40	143
rect	39	145	40	146
rect	39	148	40	149
rect	39	151	40	152
rect	39	154	40	155
rect	39	157	40	158
rect	39	160	40	161
rect	39	163	40	164
rect	39	166	40	167
rect	39	169	40	170
rect	39	172	40	173
rect	39	175	40	176
rect	39	178	40	179
rect	39	181	40	182
rect	39	184	40	185
rect	39	187	40	188
rect	39	190	40	191
rect	39	193	40	194
rect	39	196	40	197
rect	39	199	40	200
rect	39	202	40	203
rect	39	205	40	206
rect	39	208	40	209
rect	39	211	40	212
rect	39	214	40	215
rect	39	217	40	218
rect	39	220	40	221
rect	39	223	40	224
rect	39	226	40	227
rect	39	229	40	230
rect	39	232	40	233
rect	39	235	40	236
rect	39	238	40	239
rect	39	241	40	242
rect	39	244	40	245
rect	39	247	40	248
rect	39	250	40	251
rect	39	253	40	254
rect	39	256	40	257
rect	39	259	40	260
rect	39	262	40	263
rect	39	265	40	266
rect	39	268	40	269
rect	39	271	40	272
rect	39	274	40	275
rect	39	277	40	278
rect	39	280	40	281
rect	39	283	40	284
rect	39	286	40	287
rect	39	289	40	290
rect	39	292	40	293
rect	39	295	40	296
rect	39	298	40	299
rect	39	301	40	302
rect	39	304	40	305
rect	39	307	40	308
rect	39	310	40	311
rect	39	313	40	314
rect	39	316	40	317
rect	39	319	40	320
rect	39	322	40	323
rect	39	325	40	326
rect	39	328	40	329
rect	39	331	40	332
rect	39	334	40	335
rect	39	337	40	338
rect	39	340	40	341
rect	39	343	40	344
rect	39	346	40	347
rect	39	349	40	350
rect	39	352	40	353
rect	39	355	40	356
rect	39	358	40	359
rect	39	361	40	362
rect	39	364	40	365
rect	39	367	40	368
rect	39	373	40	374
rect	39	376	40	377
rect	39	379	40	380
rect	39	385	40	386
rect	40	1	41	2
rect	40	4	41	5
rect	40	7	41	8
rect	40	10	41	11
rect	40	13	41	14
rect	40	16	41	17
rect	40	19	41	20
rect	40	22	41	23
rect	40	25	41	26
rect	40	28	41	29
rect	40	31	41	32
rect	40	34	41	35
rect	40	37	41	38
rect	40	40	41	41
rect	40	43	41	44
rect	40	46	41	47
rect	40	49	41	50
rect	40	52	41	53
rect	40	55	41	56
rect	40	58	41	59
rect	40	61	41	62
rect	40	64	41	65
rect	40	67	41	68
rect	40	70	41	71
rect	40	73	41	74
rect	40	76	41	77
rect	40	79	41	80
rect	40	82	41	83
rect	40	85	41	86
rect	40	88	41	89
rect	40	91	41	92
rect	40	94	41	95
rect	40	97	41	98
rect	40	100	41	101
rect	40	103	41	104
rect	40	106	41	107
rect	40	109	41	110
rect	40	112	41	113
rect	40	115	41	116
rect	40	118	41	119
rect	40	121	41	122
rect	40	124	41	125
rect	40	127	41	128
rect	40	130	41	131
rect	40	133	41	134
rect	40	136	41	137
rect	40	139	41	140
rect	40	142	41	143
rect	40	145	41	146
rect	40	148	41	149
rect	40	151	41	152
rect	40	154	41	155
rect	40	157	41	158
rect	40	160	41	161
rect	40	163	41	164
rect	40	166	41	167
rect	40	169	41	170
rect	40	172	41	173
rect	40	175	41	176
rect	40	178	41	179
rect	40	181	41	182
rect	40	184	41	185
rect	40	187	41	188
rect	40	190	41	191
rect	40	193	41	194
rect	40	196	41	197
rect	40	199	41	200
rect	40	202	41	203
rect	40	205	41	206
rect	40	208	41	209
rect	40	211	41	212
rect	40	214	41	215
rect	40	217	41	218
rect	40	220	41	221
rect	40	223	41	224
rect	40	226	41	227
rect	40	229	41	230
rect	40	232	41	233
rect	40	235	41	236
rect	40	238	41	239
rect	40	241	41	242
rect	40	244	41	245
rect	40	247	41	248
rect	40	250	41	251
rect	40	253	41	254
rect	40	256	41	257
rect	40	259	41	260
rect	40	262	41	263
rect	40	265	41	266
rect	40	268	41	269
rect	40	271	41	272
rect	40	274	41	275
rect	40	277	41	278
rect	40	280	41	281
rect	40	283	41	284
rect	40	286	41	287
rect	40	289	41	290
rect	40	292	41	293
rect	40	295	41	296
rect	40	298	41	299
rect	40	301	41	302
rect	40	304	41	305
rect	40	307	41	308
rect	40	310	41	311
rect	40	313	41	314
rect	40	316	41	317
rect	40	319	41	320
rect	40	322	41	323
rect	40	325	41	326
rect	40	328	41	329
rect	40	331	41	332
rect	40	334	41	335
rect	40	337	41	338
rect	40	340	41	341
rect	40	343	41	344
rect	40	346	41	347
rect	40	349	41	350
rect	40	352	41	353
rect	40	355	41	356
rect	40	358	41	359
rect	40	361	41	362
rect	40	364	41	365
rect	40	367	41	368
rect	40	373	41	374
rect	40	376	41	377
rect	40	379	41	380
rect	40	385	41	386
rect	41	1	42	2
rect	41	4	42	5
rect	41	7	42	8
rect	41	10	42	11
rect	41	13	42	14
rect	41	16	42	17
rect	41	19	42	20
rect	41	22	42	23
rect	41	25	42	26
rect	41	28	42	29
rect	41	31	42	32
rect	41	34	42	35
rect	41	37	42	38
rect	41	40	42	41
rect	41	43	42	44
rect	41	46	42	47
rect	41	49	42	50
rect	41	52	42	53
rect	41	55	42	56
rect	41	58	42	59
rect	41	61	42	62
rect	41	64	42	65
rect	41	67	42	68
rect	41	70	42	71
rect	41	73	42	74
rect	41	76	42	77
rect	41	79	42	80
rect	41	82	42	83
rect	41	85	42	86
rect	41	88	42	89
rect	41	91	42	92
rect	41	94	42	95
rect	41	97	42	98
rect	41	100	42	101
rect	41	103	42	104
rect	41	106	42	107
rect	41	109	42	110
rect	41	112	42	113
rect	41	115	42	116
rect	41	118	42	119
rect	41	121	42	122
rect	41	124	42	125
rect	41	127	42	128
rect	41	130	42	131
rect	41	133	42	134
rect	41	136	42	137
rect	41	139	42	140
rect	41	142	42	143
rect	41	145	42	146
rect	41	148	42	149
rect	41	151	42	152
rect	41	154	42	155
rect	41	157	42	158
rect	41	160	42	161
rect	41	163	42	164
rect	41	166	42	167
rect	41	169	42	170
rect	41	172	42	173
rect	41	175	42	176
rect	41	178	42	179
rect	41	181	42	182
rect	41	184	42	185
rect	41	187	42	188
rect	41	190	42	191
rect	41	193	42	194
rect	41	196	42	197
rect	41	199	42	200
rect	41	202	42	203
rect	41	205	42	206
rect	41	208	42	209
rect	41	211	42	212
rect	41	214	42	215
rect	41	217	42	218
rect	41	220	42	221
rect	41	223	42	224
rect	41	226	42	227
rect	41	229	42	230
rect	41	232	42	233
rect	41	235	42	236
rect	41	238	42	239
rect	41	241	42	242
rect	41	244	42	245
rect	41	247	42	248
rect	41	250	42	251
rect	41	253	42	254
rect	41	256	42	257
rect	41	259	42	260
rect	41	262	42	263
rect	41	265	42	266
rect	41	268	42	269
rect	41	271	42	272
rect	41	274	42	275
rect	41	277	42	278
rect	41	280	42	281
rect	41	283	42	284
rect	41	286	42	287
rect	41	289	42	290
rect	41	292	42	293
rect	41	295	42	296
rect	41	298	42	299
rect	41	301	42	302
rect	41	304	42	305
rect	41	307	42	308
rect	41	310	42	311
rect	41	313	42	314
rect	41	316	42	317
rect	41	319	42	320
rect	41	322	42	323
rect	41	325	42	326
rect	41	328	42	329
rect	41	331	42	332
rect	41	334	42	335
rect	41	337	42	338
rect	41	340	42	341
rect	41	343	42	344
rect	41	346	42	347
rect	41	349	42	350
rect	41	352	42	353
rect	41	355	42	356
rect	41	358	42	359
rect	41	361	42	362
rect	41	364	42	365
rect	41	367	42	368
rect	41	373	42	374
rect	41	376	42	377
rect	41	379	42	380
rect	41	385	42	386
rect	42	1	43	2
rect	42	4	43	5
rect	42	7	43	8
rect	42	10	43	11
rect	42	13	43	14
rect	42	16	43	17
rect	42	19	43	20
rect	42	22	43	23
rect	42	25	43	26
rect	42	28	43	29
rect	42	31	43	32
rect	42	34	43	35
rect	42	37	43	38
rect	42	40	43	41
rect	42	43	43	44
rect	42	46	43	47
rect	42	49	43	50
rect	42	52	43	53
rect	42	55	43	56
rect	42	58	43	59
rect	42	61	43	62
rect	42	64	43	65
rect	42	67	43	68
rect	42	70	43	71
rect	42	73	43	74
rect	42	76	43	77
rect	42	79	43	80
rect	42	82	43	83
rect	42	85	43	86
rect	42	88	43	89
rect	42	91	43	92
rect	42	94	43	95
rect	42	97	43	98
rect	42	100	43	101
rect	42	103	43	104
rect	42	106	43	107
rect	42	109	43	110
rect	42	112	43	113
rect	42	115	43	116
rect	42	118	43	119
rect	42	121	43	122
rect	42	124	43	125
rect	42	127	43	128
rect	42	130	43	131
rect	42	133	43	134
rect	42	136	43	137
rect	42	139	43	140
rect	42	142	43	143
rect	42	145	43	146
rect	42	148	43	149
rect	42	151	43	152
rect	42	154	43	155
rect	42	157	43	158
rect	42	160	43	161
rect	42	163	43	164
rect	42	166	43	167
rect	42	169	43	170
rect	42	172	43	173
rect	42	175	43	176
rect	42	178	43	179
rect	42	181	43	182
rect	42	184	43	185
rect	42	187	43	188
rect	42	190	43	191
rect	42	193	43	194
rect	42	196	43	197
rect	42	199	43	200
rect	42	202	43	203
rect	42	205	43	206
rect	42	208	43	209
rect	42	211	43	212
rect	42	214	43	215
rect	42	217	43	218
rect	42	220	43	221
rect	42	223	43	224
rect	42	226	43	227
rect	42	229	43	230
rect	42	232	43	233
rect	42	235	43	236
rect	42	238	43	239
rect	42	241	43	242
rect	42	244	43	245
rect	42	247	43	248
rect	42	250	43	251
rect	42	253	43	254
rect	42	256	43	257
rect	42	259	43	260
rect	42	262	43	263
rect	42	265	43	266
rect	42	268	43	269
rect	42	271	43	272
rect	42	274	43	275
rect	42	277	43	278
rect	42	280	43	281
rect	42	283	43	284
rect	42	286	43	287
rect	42	289	43	290
rect	42	292	43	293
rect	42	295	43	296
rect	42	298	43	299
rect	42	301	43	302
rect	42	304	43	305
rect	42	307	43	308
rect	42	310	43	311
rect	42	313	43	314
rect	42	316	43	317
rect	42	319	43	320
rect	42	322	43	323
rect	42	325	43	326
rect	42	328	43	329
rect	42	331	43	332
rect	42	334	43	335
rect	42	337	43	338
rect	42	340	43	341
rect	42	343	43	344
rect	42	346	43	347
rect	42	349	43	350
rect	42	352	43	353
rect	42	355	43	356
rect	42	358	43	359
rect	42	361	43	362
rect	42	364	43	365
rect	42	367	43	368
rect	42	373	43	374
rect	42	376	43	377
rect	42	379	43	380
rect	42	385	43	386
rect	43	1	44	2
rect	43	4	44	5
rect	43	7	44	8
rect	43	10	44	11
rect	43	13	44	14
rect	43	16	44	17
rect	43	19	44	20
rect	43	22	44	23
rect	43	25	44	26
rect	43	28	44	29
rect	43	31	44	32
rect	43	34	44	35
rect	43	37	44	38
rect	43	40	44	41
rect	43	43	44	44
rect	43	46	44	47
rect	43	49	44	50
rect	43	52	44	53
rect	43	55	44	56
rect	43	58	44	59
rect	43	61	44	62
rect	43	64	44	65
rect	43	67	44	68
rect	43	70	44	71
rect	43	73	44	74
rect	43	76	44	77
rect	43	79	44	80
rect	43	82	44	83
rect	43	85	44	86
rect	43	88	44	89
rect	43	91	44	92
rect	43	94	44	95
rect	43	97	44	98
rect	43	100	44	101
rect	43	103	44	104
rect	43	106	44	107
rect	43	109	44	110
rect	43	112	44	113
rect	43	115	44	116
rect	43	118	44	119
rect	43	121	44	122
rect	43	124	44	125
rect	43	127	44	128
rect	43	130	44	131
rect	43	133	44	134
rect	43	136	44	137
rect	43	139	44	140
rect	43	142	44	143
rect	43	145	44	146
rect	43	148	44	149
rect	43	151	44	152
rect	43	154	44	155
rect	43	157	44	158
rect	43	160	44	161
rect	43	163	44	164
rect	43	166	44	167
rect	43	169	44	170
rect	43	172	44	173
rect	43	175	44	176
rect	43	178	44	179
rect	43	181	44	182
rect	43	184	44	185
rect	43	187	44	188
rect	43	190	44	191
rect	43	193	44	194
rect	43	196	44	197
rect	43	199	44	200
rect	43	202	44	203
rect	43	205	44	206
rect	43	208	44	209
rect	43	211	44	212
rect	43	214	44	215
rect	43	217	44	218
rect	43	220	44	221
rect	43	223	44	224
rect	43	226	44	227
rect	43	229	44	230
rect	43	232	44	233
rect	43	235	44	236
rect	43	238	44	239
rect	43	241	44	242
rect	43	244	44	245
rect	43	247	44	248
rect	43	250	44	251
rect	43	253	44	254
rect	43	256	44	257
rect	43	259	44	260
rect	43	262	44	263
rect	43	265	44	266
rect	43	268	44	269
rect	43	271	44	272
rect	43	274	44	275
rect	43	277	44	278
rect	43	280	44	281
rect	43	283	44	284
rect	43	286	44	287
rect	43	289	44	290
rect	43	292	44	293
rect	43	295	44	296
rect	43	298	44	299
rect	43	301	44	302
rect	43	304	44	305
rect	43	307	44	308
rect	43	310	44	311
rect	43	313	44	314
rect	43	316	44	317
rect	43	319	44	320
rect	43	322	44	323
rect	43	325	44	326
rect	43	328	44	329
rect	43	331	44	332
rect	43	334	44	335
rect	43	337	44	338
rect	43	340	44	341
rect	43	343	44	344
rect	43	346	44	347
rect	43	349	44	350
rect	43	352	44	353
rect	43	355	44	356
rect	43	358	44	359
rect	43	361	44	362
rect	43	364	44	365
rect	43	367	44	368
rect	43	373	44	374
rect	43	376	44	377
rect	43	379	44	380
rect	43	385	44	386
rect	44	1	45	2
rect	44	4	45	5
rect	44	7	45	8
rect	44	10	45	11
rect	44	13	45	14
rect	44	16	45	17
rect	44	19	45	20
rect	44	22	45	23
rect	44	25	45	26
rect	44	28	45	29
rect	44	31	45	32
rect	44	34	45	35
rect	44	37	45	38
rect	44	40	45	41
rect	44	43	45	44
rect	44	46	45	47
rect	44	49	45	50
rect	44	52	45	53
rect	44	55	45	56
rect	44	58	45	59
rect	44	61	45	62
rect	44	64	45	65
rect	44	67	45	68
rect	44	70	45	71
rect	44	73	45	74
rect	44	76	45	77
rect	44	79	45	80
rect	44	82	45	83
rect	44	85	45	86
rect	44	88	45	89
rect	44	91	45	92
rect	44	94	45	95
rect	44	97	45	98
rect	44	100	45	101
rect	44	103	45	104
rect	44	106	45	107
rect	44	109	45	110
rect	44	112	45	113
rect	44	115	45	116
rect	44	118	45	119
rect	44	121	45	122
rect	44	124	45	125
rect	44	127	45	128
rect	44	130	45	131
rect	44	133	45	134
rect	44	136	45	137
rect	44	139	45	140
rect	44	142	45	143
rect	44	145	45	146
rect	44	148	45	149
rect	44	151	45	152
rect	44	154	45	155
rect	44	157	45	158
rect	44	160	45	161
rect	44	163	45	164
rect	44	166	45	167
rect	44	169	45	170
rect	44	172	45	173
rect	44	175	45	176
rect	44	178	45	179
rect	44	181	45	182
rect	44	184	45	185
rect	44	187	45	188
rect	44	190	45	191
rect	44	193	45	194
rect	44	196	45	197
rect	44	199	45	200
rect	44	202	45	203
rect	44	205	45	206
rect	44	208	45	209
rect	44	211	45	212
rect	44	214	45	215
rect	44	217	45	218
rect	44	220	45	221
rect	44	223	45	224
rect	44	226	45	227
rect	44	229	45	230
rect	44	232	45	233
rect	44	235	45	236
rect	44	238	45	239
rect	44	241	45	242
rect	44	244	45	245
rect	44	247	45	248
rect	44	250	45	251
rect	44	253	45	254
rect	44	256	45	257
rect	44	259	45	260
rect	44	262	45	263
rect	44	265	45	266
rect	44	268	45	269
rect	44	271	45	272
rect	44	274	45	275
rect	44	277	45	278
rect	44	280	45	281
rect	44	283	45	284
rect	44	286	45	287
rect	44	289	45	290
rect	44	292	45	293
rect	44	295	45	296
rect	44	298	45	299
rect	44	301	45	302
rect	44	304	45	305
rect	44	307	45	308
rect	44	310	45	311
rect	44	313	45	314
rect	44	316	45	317
rect	44	319	45	320
rect	44	322	45	323
rect	44	325	45	326
rect	44	328	45	329
rect	44	331	45	332
rect	44	334	45	335
rect	44	337	45	338
rect	44	340	45	341
rect	44	343	45	344
rect	44	346	45	347
rect	44	349	45	350
rect	44	352	45	353
rect	44	355	45	356
rect	44	358	45	359
rect	44	361	45	362
rect	44	364	45	365
rect	44	367	45	368
rect	44	373	45	374
rect	44	376	45	377
rect	44	379	45	380
rect	44	385	45	386
rect	45	1	46	2
rect	45	4	46	5
rect	45	7	46	8
rect	45	10	46	11
rect	45	13	46	14
rect	45	16	46	17
rect	45	19	46	20
rect	45	22	46	23
rect	45	25	46	26
rect	45	28	46	29
rect	45	31	46	32
rect	45	34	46	35
rect	45	37	46	38
rect	45	40	46	41
rect	45	43	46	44
rect	45	46	46	47
rect	45	49	46	50
rect	45	52	46	53
rect	45	55	46	56
rect	45	58	46	59
rect	45	61	46	62
rect	45	64	46	65
rect	45	67	46	68
rect	45	70	46	71
rect	45	73	46	74
rect	45	76	46	77
rect	45	79	46	80
rect	45	82	46	83
rect	45	85	46	86
rect	45	88	46	89
rect	45	91	46	92
rect	45	94	46	95
rect	45	97	46	98
rect	45	100	46	101
rect	45	103	46	104
rect	45	106	46	107
rect	45	109	46	110
rect	45	112	46	113
rect	45	115	46	116
rect	45	118	46	119
rect	45	121	46	122
rect	45	124	46	125
rect	45	127	46	128
rect	45	130	46	131
rect	45	133	46	134
rect	45	136	46	137
rect	45	139	46	140
rect	45	142	46	143
rect	45	145	46	146
rect	45	148	46	149
rect	45	151	46	152
rect	45	154	46	155
rect	45	157	46	158
rect	45	160	46	161
rect	45	163	46	164
rect	45	166	46	167
rect	45	169	46	170
rect	45	172	46	173
rect	45	175	46	176
rect	45	178	46	179
rect	45	181	46	182
rect	45	184	46	185
rect	45	187	46	188
rect	45	190	46	191
rect	45	193	46	194
rect	45	196	46	197
rect	45	199	46	200
rect	45	202	46	203
rect	45	205	46	206
rect	45	208	46	209
rect	45	211	46	212
rect	45	214	46	215
rect	45	217	46	218
rect	45	220	46	221
rect	45	223	46	224
rect	45	226	46	227
rect	45	229	46	230
rect	45	232	46	233
rect	45	235	46	236
rect	45	238	46	239
rect	45	241	46	242
rect	45	244	46	245
rect	45	247	46	248
rect	45	250	46	251
rect	45	253	46	254
rect	45	256	46	257
rect	45	259	46	260
rect	45	262	46	263
rect	45	265	46	266
rect	45	268	46	269
rect	45	271	46	272
rect	45	274	46	275
rect	45	277	46	278
rect	45	280	46	281
rect	45	283	46	284
rect	45	286	46	287
rect	45	289	46	290
rect	45	292	46	293
rect	45	295	46	296
rect	45	298	46	299
rect	45	301	46	302
rect	45	304	46	305
rect	45	307	46	308
rect	45	310	46	311
rect	45	313	46	314
rect	45	316	46	317
rect	45	319	46	320
rect	45	322	46	323
rect	45	325	46	326
rect	45	328	46	329
rect	45	331	46	332
rect	45	334	46	335
rect	45	337	46	338
rect	45	340	46	341
rect	45	343	46	344
rect	45	346	46	347
rect	45	349	46	350
rect	45	352	46	353
rect	45	355	46	356
rect	45	358	46	359
rect	45	361	46	362
rect	45	364	46	365
rect	45	367	46	368
rect	45	373	46	374
rect	45	376	46	377
rect	45	379	46	380
rect	45	385	46	386
rect	46	1	47	2
rect	46	4	47	5
rect	46	7	47	8
rect	46	10	47	11
rect	46	13	47	14
rect	46	16	47	17
rect	46	19	47	20
rect	46	22	47	23
rect	46	25	47	26
rect	46	28	47	29
rect	46	31	47	32
rect	46	34	47	35
rect	46	37	47	38
rect	46	40	47	41
rect	46	43	47	44
rect	46	46	47	47
rect	46	49	47	50
rect	46	52	47	53
rect	46	55	47	56
rect	46	58	47	59
rect	46	61	47	62
rect	46	64	47	65
rect	46	67	47	68
rect	46	70	47	71
rect	46	73	47	74
rect	46	76	47	77
rect	46	79	47	80
rect	46	82	47	83
rect	46	85	47	86
rect	46	88	47	89
rect	46	91	47	92
rect	46	94	47	95
rect	46	97	47	98
rect	46	100	47	101
rect	46	103	47	104
rect	46	106	47	107
rect	46	109	47	110
rect	46	112	47	113
rect	46	115	47	116
rect	46	118	47	119
rect	46	121	47	122
rect	46	124	47	125
rect	46	127	47	128
rect	46	130	47	131
rect	46	133	47	134
rect	46	136	47	137
rect	46	139	47	140
rect	46	142	47	143
rect	46	145	47	146
rect	46	148	47	149
rect	46	151	47	152
rect	46	154	47	155
rect	46	157	47	158
rect	46	160	47	161
rect	46	163	47	164
rect	46	166	47	167
rect	46	169	47	170
rect	46	172	47	173
rect	46	175	47	176
rect	46	178	47	179
rect	46	184	47	185
rect	46	187	47	188
rect	46	190	47	191
rect	46	193	47	194
rect	46	196	47	197
rect	46	199	47	200
rect	46	202	47	203
rect	46	205	47	206
rect	46	208	47	209
rect	46	211	47	212
rect	46	214	47	215
rect	46	217	47	218
rect	46	220	47	221
rect	46	223	47	224
rect	46	226	47	227
rect	46	229	47	230
rect	46	232	47	233
rect	46	235	47	236
rect	46	238	47	239
rect	46	244	47	245
rect	46	247	47	248
rect	46	250	47	251
rect	46	253	47	254
rect	46	256	47	257
rect	46	259	47	260
rect	46	262	47	263
rect	46	265	47	266
rect	46	268	47	269
rect	46	271	47	272
rect	46	274	47	275
rect	46	277	47	278
rect	46	280	47	281
rect	46	283	47	284
rect	46	286	47	287
rect	46	289	47	290
rect	46	292	47	293
rect	46	295	47	296
rect	46	298	47	299
rect	46	301	47	302
rect	46	304	47	305
rect	46	307	47	308
rect	46	310	47	311
rect	46	313	47	314
rect	46	316	47	317
rect	46	319	47	320
rect	46	322	47	323
rect	46	325	47	326
rect	46	328	47	329
rect	46	331	47	332
rect	46	334	47	335
rect	46	337	47	338
rect	46	340	47	341
rect	46	343	47	344
rect	46	346	47	347
rect	46	349	47	350
rect	46	352	47	353
rect	46	355	47	356
rect	46	358	47	359
rect	46	361	47	362
rect	46	364	47	365
rect	46	367	47	368
rect	46	373	47	374
rect	46	376	47	377
rect	46	379	47	380
rect	46	385	47	386
rect	47	1	48	2
rect	47	4	48	5
rect	47	7	48	8
rect	47	10	48	11
rect	47	13	48	14
rect	47	16	48	17
rect	47	19	48	20
rect	47	22	48	23
rect	47	25	48	26
rect	47	28	48	29
rect	47	31	48	32
rect	47	34	48	35
rect	47	37	48	38
rect	47	40	48	41
rect	47	43	48	44
rect	47	46	48	47
rect	47	49	48	50
rect	47	52	48	53
rect	47	55	48	56
rect	47	58	48	59
rect	47	61	48	62
rect	47	64	48	65
rect	47	67	48	68
rect	47	70	48	71
rect	47	73	48	74
rect	47	76	48	77
rect	47	79	48	80
rect	47	82	48	83
rect	47	85	48	86
rect	47	88	48	89
rect	47	91	48	92
rect	47	94	48	95
rect	47	97	48	98
rect	47	100	48	101
rect	47	103	48	104
rect	47	106	48	107
rect	47	109	48	110
rect	47	112	48	113
rect	47	115	48	116
rect	47	118	48	119
rect	47	121	48	122
rect	47	124	48	125
rect	47	127	48	128
rect	47	130	48	131
rect	47	133	48	134
rect	47	136	48	137
rect	47	139	48	140
rect	47	142	48	143
rect	47	145	48	146
rect	47	148	48	149
rect	47	151	48	152
rect	47	154	48	155
rect	47	157	48	158
rect	47	160	48	161
rect	47	163	48	164
rect	47	166	48	167
rect	47	169	48	170
rect	47	172	48	173
rect	47	175	48	176
rect	47	178	48	179
rect	47	181	48	182
rect	47	184	48	185
rect	47	187	48	188
rect	47	190	48	191
rect	47	193	48	194
rect	47	196	48	197
rect	47	199	48	200
rect	47	202	48	203
rect	47	205	48	206
rect	47	208	48	209
rect	47	211	48	212
rect	47	214	48	215
rect	47	217	48	218
rect	47	220	48	221
rect	47	223	48	224
rect	47	226	48	227
rect	47	229	48	230
rect	47	232	48	233
rect	47	235	48	236
rect	47	238	48	239
rect	47	241	48	242
rect	47	244	48	245
rect	47	247	48	248
rect	47	250	48	251
rect	47	253	48	254
rect	47	256	48	257
rect	47	259	48	260
rect	47	262	48	263
rect	47	265	48	266
rect	47	268	48	269
rect	47	271	48	272
rect	47	274	48	275
rect	47	277	48	278
rect	47	280	48	281
rect	47	283	48	284
rect	47	286	48	287
rect	47	289	48	290
rect	47	292	48	293
rect	47	295	48	296
rect	47	298	48	299
rect	47	301	48	302
rect	47	304	48	305
rect	47	307	48	308
rect	47	310	48	311
rect	47	313	48	314
rect	47	316	48	317
rect	47	319	48	320
rect	47	322	48	323
rect	47	325	48	326
rect	47	328	48	329
rect	47	331	48	332
rect	47	334	48	335
rect	47	337	48	338
rect	47	340	48	341
rect	47	343	48	344
rect	47	346	48	347
rect	47	349	48	350
rect	47	352	48	353
rect	47	355	48	356
rect	47	358	48	359
rect	47	361	48	362
rect	47	364	48	365
rect	47	367	48	368
rect	47	373	48	374
rect	47	376	48	377
rect	47	379	48	380
rect	47	385	48	386
rect	48	1	49	2
rect	48	4	49	5
rect	48	7	49	8
rect	48	10	49	11
rect	48	13	49	14
rect	48	16	49	17
rect	48	19	49	20
rect	48	22	49	23
rect	48	25	49	26
rect	48	28	49	29
rect	48	31	49	32
rect	48	34	49	35
rect	48	37	49	38
rect	48	40	49	41
rect	48	43	49	44
rect	48	46	49	47
rect	48	49	49	50
rect	48	52	49	53
rect	48	55	49	56
rect	48	58	49	59
rect	48	61	49	62
rect	48	64	49	65
rect	48	67	49	68
rect	48	70	49	71
rect	48	73	49	74
rect	48	76	49	77
rect	48	79	49	80
rect	48	82	49	83
rect	48	85	49	86
rect	48	88	49	89
rect	48	91	49	92
rect	48	94	49	95
rect	48	97	49	98
rect	48	100	49	101
rect	48	103	49	104
rect	48	106	49	107
rect	48	109	49	110
rect	48	112	49	113
rect	48	115	49	116
rect	48	118	49	119
rect	48	121	49	122
rect	48	124	49	125
rect	48	127	49	128
rect	48	130	49	131
rect	48	133	49	134
rect	48	136	49	137
rect	48	139	49	140
rect	48	142	49	143
rect	48	145	49	146
rect	48	148	49	149
rect	48	151	49	152
rect	48	154	49	155
rect	48	157	49	158
rect	48	160	49	161
rect	48	163	49	164
rect	48	166	49	167
rect	48	169	49	170
rect	48	172	49	173
rect	48	175	49	176
rect	48	178	49	179
rect	48	181	49	182
rect	48	184	49	185
rect	48	187	49	188
rect	48	190	49	191
rect	48	193	49	194
rect	48	196	49	197
rect	48	199	49	200
rect	48	202	49	203
rect	48	205	49	206
rect	48	208	49	209
rect	48	211	49	212
rect	48	214	49	215
rect	48	217	49	218
rect	48	220	49	221
rect	48	223	49	224
rect	48	226	49	227
rect	48	229	49	230
rect	48	232	49	233
rect	48	235	49	236
rect	48	238	49	239
rect	48	241	49	242
rect	48	244	49	245
rect	48	247	49	248
rect	48	250	49	251
rect	48	253	49	254
rect	48	256	49	257
rect	48	259	49	260
rect	48	262	49	263
rect	48	265	49	266
rect	48	268	49	269
rect	48	271	49	272
rect	48	274	49	275
rect	48	277	49	278
rect	48	280	49	281
rect	48	283	49	284
rect	48	286	49	287
rect	48	289	49	290
rect	48	292	49	293
rect	48	295	49	296
rect	48	298	49	299
rect	48	301	49	302
rect	48	304	49	305
rect	48	307	49	308
rect	48	310	49	311
rect	48	313	49	314
rect	48	316	49	317
rect	48	319	49	320
rect	48	322	49	323
rect	48	325	49	326
rect	48	328	49	329
rect	48	331	49	332
rect	48	334	49	335
rect	48	337	49	338
rect	48	340	49	341
rect	48	343	49	344
rect	48	346	49	347
rect	48	349	49	350
rect	48	352	49	353
rect	48	355	49	356
rect	48	358	49	359
rect	48	361	49	362
rect	48	364	49	365
rect	48	367	49	368
rect	48	373	49	374
rect	48	376	49	377
rect	48	379	49	380
rect	48	385	49	386
rect	49	1	50	2
rect	49	4	50	5
rect	49	7	50	8
rect	49	10	50	11
rect	49	13	50	14
rect	49	16	50	17
rect	49	19	50	20
rect	49	22	50	23
rect	49	25	50	26
rect	49	28	50	29
rect	49	31	50	32
rect	49	34	50	35
rect	49	37	50	38
rect	49	40	50	41
rect	49	43	50	44
rect	49	46	50	47
rect	49	49	50	50
rect	49	52	50	53
rect	49	55	50	56
rect	49	58	50	59
rect	49	61	50	62
rect	49	64	50	65
rect	49	67	50	68
rect	49	70	50	71
rect	49	73	50	74
rect	49	76	50	77
rect	49	79	50	80
rect	49	82	50	83
rect	49	85	50	86
rect	49	88	50	89
rect	49	91	50	92
rect	49	94	50	95
rect	49	97	50	98
rect	49	100	50	101
rect	49	103	50	104
rect	49	106	50	107
rect	49	109	50	110
rect	49	112	50	113
rect	49	115	50	116
rect	49	118	50	119
rect	49	121	50	122
rect	49	124	50	125
rect	49	127	50	128
rect	49	130	50	131
rect	49	133	50	134
rect	49	136	50	137
rect	49	139	50	140
rect	49	142	50	143
rect	49	145	50	146
rect	49	148	50	149
rect	49	151	50	152
rect	49	154	50	155
rect	49	157	50	158
rect	49	160	50	161
rect	49	163	50	164
rect	49	166	50	167
rect	49	169	50	170
rect	49	172	50	173
rect	49	175	50	176
rect	49	178	50	179
rect	49	181	50	182
rect	49	184	50	185
rect	49	187	50	188
rect	49	190	50	191
rect	49	193	50	194
rect	49	196	50	197
rect	49	199	50	200
rect	49	202	50	203
rect	49	205	50	206
rect	49	208	50	209
rect	49	211	50	212
rect	49	214	50	215
rect	49	217	50	218
rect	49	220	50	221
rect	49	223	50	224
rect	49	226	50	227
rect	49	229	50	230
rect	49	232	50	233
rect	49	235	50	236
rect	49	238	50	239
rect	49	241	50	242
rect	49	244	50	245
rect	49	247	50	248
rect	49	250	50	251
rect	49	253	50	254
rect	49	256	50	257
rect	49	259	50	260
rect	49	262	50	263
rect	49	265	50	266
rect	49	268	50	269
rect	49	271	50	272
rect	49	274	50	275
rect	49	277	50	278
rect	49	280	50	281
rect	49	283	50	284
rect	49	286	50	287
rect	49	289	50	290
rect	49	292	50	293
rect	49	295	50	296
rect	49	298	50	299
rect	49	301	50	302
rect	49	304	50	305
rect	49	307	50	308
rect	49	310	50	311
rect	49	313	50	314
rect	49	316	50	317
rect	49	319	50	320
rect	49	322	50	323
rect	49	325	50	326
rect	49	328	50	329
rect	49	331	50	332
rect	49	334	50	335
rect	49	337	50	338
rect	49	340	50	341
rect	49	343	50	344
rect	49	346	50	347
rect	49	349	50	350
rect	49	352	50	353
rect	49	355	50	356
rect	49	358	50	359
rect	49	361	50	362
rect	49	364	50	365
rect	49	367	50	368
rect	49	373	50	374
rect	49	376	50	377
rect	49	379	50	380
rect	49	385	50	386
rect	50	1	51	2
rect	50	4	51	5
rect	50	7	51	8
rect	50	10	51	11
rect	50	13	51	14
rect	50	16	51	17
rect	50	19	51	20
rect	50	22	51	23
rect	50	25	51	26
rect	50	28	51	29
rect	50	31	51	32
rect	50	34	51	35
rect	50	37	51	38
rect	50	40	51	41
rect	50	43	51	44
rect	50	46	51	47
rect	50	49	51	50
rect	50	52	51	53
rect	50	55	51	56
rect	50	58	51	59
rect	50	61	51	62
rect	50	64	51	65
rect	50	67	51	68
rect	50	70	51	71
rect	50	73	51	74
rect	50	76	51	77
rect	50	79	51	80
rect	50	82	51	83
rect	50	85	51	86
rect	50	88	51	89
rect	50	91	51	92
rect	50	94	51	95
rect	50	97	51	98
rect	50	100	51	101
rect	50	103	51	104
rect	50	106	51	107
rect	50	109	51	110
rect	50	112	51	113
rect	50	115	51	116
rect	50	118	51	119
rect	50	121	51	122
rect	50	124	51	125
rect	50	127	51	128
rect	50	130	51	131
rect	50	133	51	134
rect	50	136	51	137
rect	50	139	51	140
rect	50	142	51	143
rect	50	145	51	146
rect	50	148	51	149
rect	50	151	51	152
rect	50	154	51	155
rect	50	157	51	158
rect	50	160	51	161
rect	50	163	51	164
rect	50	166	51	167
rect	50	169	51	170
rect	50	172	51	173
rect	50	175	51	176
rect	50	178	51	179
rect	50	181	51	182
rect	50	184	51	185
rect	50	187	51	188
rect	50	190	51	191
rect	50	193	51	194
rect	50	196	51	197
rect	50	199	51	200
rect	50	202	51	203
rect	50	205	51	206
rect	50	208	51	209
rect	50	211	51	212
rect	50	214	51	215
rect	50	217	51	218
rect	50	220	51	221
rect	50	223	51	224
rect	50	226	51	227
rect	50	229	51	230
rect	50	232	51	233
rect	50	235	51	236
rect	50	238	51	239
rect	50	241	51	242
rect	50	244	51	245
rect	50	247	51	248
rect	50	250	51	251
rect	50	253	51	254
rect	50	256	51	257
rect	50	259	51	260
rect	50	262	51	263
rect	50	265	51	266
rect	50	268	51	269
rect	50	271	51	272
rect	50	274	51	275
rect	50	277	51	278
rect	50	280	51	281
rect	50	283	51	284
rect	50	286	51	287
rect	50	289	51	290
rect	50	292	51	293
rect	50	295	51	296
rect	50	298	51	299
rect	50	301	51	302
rect	50	304	51	305
rect	50	307	51	308
rect	50	310	51	311
rect	50	313	51	314
rect	50	316	51	317
rect	50	319	51	320
rect	50	322	51	323
rect	50	325	51	326
rect	50	328	51	329
rect	50	331	51	332
rect	50	334	51	335
rect	50	337	51	338
rect	50	340	51	341
rect	50	343	51	344
rect	50	346	51	347
rect	50	349	51	350
rect	50	352	51	353
rect	50	355	51	356
rect	50	358	51	359
rect	50	361	51	362
rect	50	364	51	365
rect	50	367	51	368
rect	50	373	51	374
rect	50	376	51	377
rect	50	379	51	380
rect	50	385	51	386
rect	51	1	52	2
rect	51	4	52	5
rect	51	7	52	8
rect	51	10	52	11
rect	51	13	52	14
rect	51	16	52	17
rect	51	19	52	20
rect	51	22	52	23
rect	51	25	52	26
rect	51	28	52	29
rect	51	31	52	32
rect	51	34	52	35
rect	51	37	52	38
rect	51	40	52	41
rect	51	43	52	44
rect	51	46	52	47
rect	51	49	52	50
rect	51	52	52	53
rect	51	55	52	56
rect	51	58	52	59
rect	51	61	52	62
rect	51	64	52	65
rect	51	67	52	68
rect	51	70	52	71
rect	51	73	52	74
rect	51	76	52	77
rect	51	79	52	80
rect	51	82	52	83
rect	51	85	52	86
rect	51	88	52	89
rect	51	91	52	92
rect	51	94	52	95
rect	51	97	52	98
rect	51	100	52	101
rect	51	103	52	104
rect	51	106	52	107
rect	51	109	52	110
rect	51	112	52	113
rect	51	115	52	116
rect	51	118	52	119
rect	51	121	52	122
rect	51	124	52	125
rect	51	127	52	128
rect	51	130	52	131
rect	51	133	52	134
rect	51	136	52	137
rect	51	139	52	140
rect	51	142	52	143
rect	51	145	52	146
rect	51	148	52	149
rect	51	151	52	152
rect	51	154	52	155
rect	51	157	52	158
rect	51	160	52	161
rect	51	163	52	164
rect	51	166	52	167
rect	51	169	52	170
rect	51	172	52	173
rect	51	175	52	176
rect	51	178	52	179
rect	51	181	52	182
rect	51	184	52	185
rect	51	187	52	188
rect	51	190	52	191
rect	51	193	52	194
rect	51	196	52	197
rect	51	199	52	200
rect	51	202	52	203
rect	51	205	52	206
rect	51	208	52	209
rect	51	211	52	212
rect	51	214	52	215
rect	51	217	52	218
rect	51	220	52	221
rect	51	223	52	224
rect	51	226	52	227
rect	51	229	52	230
rect	51	232	52	233
rect	51	235	52	236
rect	51	238	52	239
rect	51	241	52	242
rect	51	244	52	245
rect	51	247	52	248
rect	51	250	52	251
rect	51	253	52	254
rect	51	256	52	257
rect	51	259	52	260
rect	51	262	52	263
rect	51	265	52	266
rect	51	268	52	269
rect	51	271	52	272
rect	51	274	52	275
rect	51	277	52	278
rect	51	280	52	281
rect	51	283	52	284
rect	51	286	52	287
rect	51	289	52	290
rect	51	292	52	293
rect	51	295	52	296
rect	51	298	52	299
rect	51	301	52	302
rect	51	304	52	305
rect	51	307	52	308
rect	51	310	52	311
rect	51	313	52	314
rect	51	316	52	317
rect	51	319	52	320
rect	51	322	52	323
rect	51	325	52	326
rect	51	328	52	329
rect	51	331	52	332
rect	51	334	52	335
rect	51	337	52	338
rect	51	340	52	341
rect	51	343	52	344
rect	51	346	52	347
rect	51	349	52	350
rect	51	352	52	353
rect	51	355	52	356
rect	51	358	52	359
rect	51	361	52	362
rect	51	364	52	365
rect	51	367	52	368
rect	51	373	52	374
rect	51	376	52	377
rect	51	379	52	380
rect	51	385	52	386
rect	52	1	53	2
rect	52	4	53	5
rect	52	7	53	8
rect	52	10	53	11
rect	52	13	53	14
rect	52	16	53	17
rect	52	19	53	20
rect	52	22	53	23
rect	52	25	53	26
rect	52	28	53	29
rect	52	31	53	32
rect	52	34	53	35
rect	52	37	53	38
rect	52	40	53	41
rect	52	43	53	44
rect	52	46	53	47
rect	52	49	53	50
rect	52	52	53	53
rect	52	55	53	56
rect	52	58	53	59
rect	52	61	53	62
rect	52	64	53	65
rect	52	67	53	68
rect	52	70	53	71
rect	52	73	53	74
rect	52	76	53	77
rect	52	79	53	80
rect	52	82	53	83
rect	52	85	53	86
rect	52	88	53	89
rect	52	91	53	92
rect	52	94	53	95
rect	52	97	53	98
rect	52	100	53	101
rect	52	103	53	104
rect	52	106	53	107
rect	52	109	53	110
rect	52	112	53	113
rect	52	115	53	116
rect	52	118	53	119
rect	52	121	53	122
rect	52	124	53	125
rect	52	127	53	128
rect	52	130	53	131
rect	52	133	53	134
rect	52	136	53	137
rect	52	139	53	140
rect	52	142	53	143
rect	52	145	53	146
rect	52	148	53	149
rect	52	151	53	152
rect	52	154	53	155
rect	52	157	53	158
rect	52	160	53	161
rect	52	163	53	164
rect	52	166	53	167
rect	52	169	53	170
rect	52	172	53	173
rect	52	175	53	176
rect	52	178	53	179
rect	52	181	53	182
rect	52	184	53	185
rect	52	187	53	188
rect	52	190	53	191
rect	52	193	53	194
rect	52	196	53	197
rect	52	199	53	200
rect	52	202	53	203
rect	52	205	53	206
rect	52	208	53	209
rect	52	211	53	212
rect	52	214	53	215
rect	52	217	53	218
rect	52	220	53	221
rect	52	223	53	224
rect	52	226	53	227
rect	52	229	53	230
rect	52	232	53	233
rect	52	235	53	236
rect	52	238	53	239
rect	52	241	53	242
rect	52	244	53	245
rect	52	247	53	248
rect	52	250	53	251
rect	52	253	53	254
rect	52	256	53	257
rect	52	259	53	260
rect	52	262	53	263
rect	52	265	53	266
rect	52	268	53	269
rect	52	271	53	272
rect	52	274	53	275
rect	52	277	53	278
rect	52	280	53	281
rect	52	283	53	284
rect	52	286	53	287
rect	52	289	53	290
rect	52	292	53	293
rect	52	295	53	296
rect	52	298	53	299
rect	52	301	53	302
rect	52	304	53	305
rect	52	307	53	308
rect	52	310	53	311
rect	52	313	53	314
rect	52	316	53	317
rect	52	319	53	320
rect	52	322	53	323
rect	52	325	53	326
rect	52	328	53	329
rect	52	331	53	332
rect	52	334	53	335
rect	52	337	53	338
rect	52	340	53	341
rect	52	343	53	344
rect	52	346	53	347
rect	52	349	53	350
rect	52	352	53	353
rect	52	355	53	356
rect	52	358	53	359
rect	52	361	53	362
rect	52	364	53	365
rect	52	367	53	368
rect	52	373	53	374
rect	52	376	53	377
rect	52	379	53	380
rect	52	385	53	386
rect	53	1	54	2
rect	53	4	54	5
rect	53	7	54	8
rect	53	10	54	11
rect	53	13	54	14
rect	53	16	54	17
rect	53	19	54	20
rect	53	22	54	23
rect	53	25	54	26
rect	53	28	54	29
rect	53	31	54	32
rect	53	34	54	35
rect	53	37	54	38
rect	53	40	54	41
rect	53	43	54	44
rect	53	46	54	47
rect	53	49	54	50
rect	53	52	54	53
rect	53	55	54	56
rect	53	58	54	59
rect	53	61	54	62
rect	53	64	54	65
rect	53	67	54	68
rect	53	70	54	71
rect	53	73	54	74
rect	53	76	54	77
rect	53	79	54	80
rect	53	82	54	83
rect	53	85	54	86
rect	53	88	54	89
rect	53	91	54	92
rect	53	94	54	95
rect	53	97	54	98
rect	53	100	54	101
rect	53	103	54	104
rect	53	106	54	107
rect	53	109	54	110
rect	53	112	54	113
rect	53	115	54	116
rect	53	118	54	119
rect	53	121	54	122
rect	53	124	54	125
rect	53	127	54	128
rect	53	130	54	131
rect	53	133	54	134
rect	53	136	54	137
rect	53	139	54	140
rect	53	142	54	143
rect	53	145	54	146
rect	53	148	54	149
rect	53	151	54	152
rect	53	154	54	155
rect	53	157	54	158
rect	53	160	54	161
rect	53	163	54	164
rect	53	166	54	167
rect	53	169	54	170
rect	53	172	54	173
rect	53	175	54	176
rect	53	178	54	179
rect	53	181	54	182
rect	53	184	54	185
rect	53	187	54	188
rect	53	190	54	191
rect	53	193	54	194
rect	53	196	54	197
rect	53	199	54	200
rect	53	202	54	203
rect	53	205	54	206
rect	53	208	54	209
rect	53	211	54	212
rect	53	214	54	215
rect	53	217	54	218
rect	53	220	54	221
rect	53	223	54	224
rect	53	226	54	227
rect	53	229	54	230
rect	53	232	54	233
rect	53	235	54	236
rect	53	238	54	239
rect	53	241	54	242
rect	53	244	54	245
rect	53	247	54	248
rect	53	250	54	251
rect	53	253	54	254
rect	53	256	54	257
rect	53	259	54	260
rect	53	262	54	263
rect	53	265	54	266
rect	53	268	54	269
rect	53	271	54	272
rect	53	274	54	275
rect	53	277	54	278
rect	53	280	54	281
rect	53	283	54	284
rect	53	286	54	287
rect	53	289	54	290
rect	53	292	54	293
rect	53	295	54	296
rect	53	298	54	299
rect	53	301	54	302
rect	53	304	54	305
rect	53	307	54	308
rect	53	310	54	311
rect	53	313	54	314
rect	53	316	54	317
rect	53	319	54	320
rect	53	322	54	323
rect	53	325	54	326
rect	53	328	54	329
rect	53	331	54	332
rect	53	334	54	335
rect	53	337	54	338
rect	53	340	54	341
rect	53	343	54	344
rect	53	346	54	347
rect	53	349	54	350
rect	53	352	54	353
rect	53	355	54	356
rect	53	358	54	359
rect	53	361	54	362
rect	53	364	54	365
rect	53	367	54	368
rect	53	373	54	374
rect	53	376	54	377
rect	53	379	54	380
rect	53	385	54	386
rect	54	1	55	2
rect	54	4	55	5
rect	54	7	55	8
rect	54	10	55	11
rect	54	13	55	14
rect	54	16	55	17
rect	54	19	55	20
rect	54	22	55	23
rect	54	25	55	26
rect	54	28	55	29
rect	54	31	55	32
rect	54	34	55	35
rect	54	37	55	38
rect	54	40	55	41
rect	54	43	55	44
rect	54	46	55	47
rect	54	49	55	50
rect	54	52	55	53
rect	54	55	55	56
rect	54	58	55	59
rect	54	61	55	62
rect	54	64	55	65
rect	54	67	55	68
rect	54	70	55	71
rect	54	73	55	74
rect	54	76	55	77
rect	54	79	55	80
rect	54	82	55	83
rect	54	85	55	86
rect	54	88	55	89
rect	54	91	55	92
rect	54	94	55	95
rect	54	97	55	98
rect	54	100	55	101
rect	54	103	55	104
rect	54	106	55	107
rect	54	109	55	110
rect	54	112	55	113
rect	54	115	55	116
rect	54	118	55	119
rect	54	121	55	122
rect	54	124	55	125
rect	54	127	55	128
rect	54	130	55	131
rect	54	133	55	134
rect	54	136	55	137
rect	54	139	55	140
rect	54	142	55	143
rect	54	145	55	146
rect	54	148	55	149
rect	54	151	55	152
rect	54	154	55	155
rect	54	157	55	158
rect	54	160	55	161
rect	54	163	55	164
rect	54	166	55	167
rect	54	169	55	170
rect	54	172	55	173
rect	54	175	55	176
rect	54	178	55	179
rect	54	181	55	182
rect	54	184	55	185
rect	54	187	55	188
rect	54	190	55	191
rect	54	193	55	194
rect	54	196	55	197
rect	54	199	55	200
rect	54	202	55	203
rect	54	205	55	206
rect	54	208	55	209
rect	54	211	55	212
rect	54	214	55	215
rect	54	217	55	218
rect	54	220	55	221
rect	54	223	55	224
rect	54	226	55	227
rect	54	229	55	230
rect	54	232	55	233
rect	54	235	55	236
rect	54	238	55	239
rect	54	241	55	242
rect	54	244	55	245
rect	54	247	55	248
rect	54	250	55	251
rect	54	253	55	254
rect	54	256	55	257
rect	54	259	55	260
rect	54	262	55	263
rect	54	265	55	266
rect	54	268	55	269
rect	54	271	55	272
rect	54	274	55	275
rect	54	277	55	278
rect	54	280	55	281
rect	54	283	55	284
rect	54	286	55	287
rect	54	289	55	290
rect	54	292	55	293
rect	54	295	55	296
rect	54	298	55	299
rect	54	301	55	302
rect	54	304	55	305
rect	54	307	55	308
rect	54	310	55	311
rect	54	313	55	314
rect	54	316	55	317
rect	54	319	55	320
rect	54	322	55	323
rect	54	325	55	326
rect	54	328	55	329
rect	54	331	55	332
rect	54	334	55	335
rect	54	337	55	338
rect	54	340	55	341
rect	54	343	55	344
rect	54	346	55	347
rect	54	349	55	350
rect	54	352	55	353
rect	54	355	55	356
rect	54	358	55	359
rect	54	361	55	362
rect	54	364	55	365
rect	54	367	55	368
rect	54	373	55	374
rect	54	376	55	377
rect	54	379	55	380
rect	54	385	55	386
rect	55	1	56	2
rect	55	4	56	5
rect	55	7	56	8
rect	55	10	56	11
rect	55	13	56	14
rect	55	16	56	17
rect	55	19	56	20
rect	55	22	56	23
rect	55	25	56	26
rect	55	28	56	29
rect	55	31	56	32
rect	55	34	56	35
rect	55	37	56	38
rect	55	40	56	41
rect	55	43	56	44
rect	55	46	56	47
rect	55	49	56	50
rect	55	52	56	53
rect	55	55	56	56
rect	55	58	56	59
rect	55	61	56	62
rect	55	64	56	65
rect	55	67	56	68
rect	55	70	56	71
rect	55	73	56	74
rect	55	76	56	77
rect	55	79	56	80
rect	55	82	56	83
rect	55	85	56	86
rect	55	88	56	89
rect	55	91	56	92
rect	55	94	56	95
rect	55	97	56	98
rect	55	100	56	101
rect	55	103	56	104
rect	55	106	56	107
rect	55	109	56	110
rect	55	112	56	113
rect	55	115	56	116
rect	55	118	56	119
rect	55	121	56	122
rect	55	124	56	125
rect	55	127	56	128
rect	55	130	56	131
rect	55	133	56	134
rect	55	136	56	137
rect	55	139	56	140
rect	55	142	56	143
rect	55	145	56	146
rect	55	148	56	149
rect	55	151	56	152
rect	55	154	56	155
rect	55	157	56	158
rect	55	160	56	161
rect	55	163	56	164
rect	55	166	56	167
rect	55	169	56	170
rect	55	172	56	173
rect	55	175	56	176
rect	55	178	56	179
rect	55	181	56	182
rect	55	184	56	185
rect	55	187	56	188
rect	55	190	56	191
rect	55	193	56	194
rect	55	196	56	197
rect	55	199	56	200
rect	55	202	56	203
rect	55	205	56	206
rect	55	208	56	209
rect	55	211	56	212
rect	55	214	56	215
rect	55	217	56	218
rect	55	220	56	221
rect	55	223	56	224
rect	55	226	56	227
rect	55	229	56	230
rect	55	232	56	233
rect	55	235	56	236
rect	55	238	56	239
rect	55	241	56	242
rect	55	244	56	245
rect	55	247	56	248
rect	55	250	56	251
rect	55	253	56	254
rect	55	256	56	257
rect	55	259	56	260
rect	55	262	56	263
rect	55	265	56	266
rect	55	268	56	269
rect	55	271	56	272
rect	55	274	56	275
rect	55	277	56	278
rect	55	280	56	281
rect	55	283	56	284
rect	55	286	56	287
rect	55	289	56	290
rect	55	292	56	293
rect	55	295	56	296
rect	55	298	56	299
rect	55	301	56	302
rect	55	304	56	305
rect	55	307	56	308
rect	55	310	56	311
rect	55	313	56	314
rect	55	316	56	317
rect	55	319	56	320
rect	55	322	56	323
rect	55	325	56	326
rect	55	328	56	329
rect	55	331	56	332
rect	55	334	56	335
rect	55	337	56	338
rect	55	340	56	341
rect	55	343	56	344
rect	55	346	56	347
rect	55	349	56	350
rect	55	352	56	353
rect	55	355	56	356
rect	55	358	56	359
rect	55	361	56	362
rect	55	364	56	365
rect	55	367	56	368
rect	55	373	56	374
rect	55	376	56	377
rect	55	379	56	380
rect	55	385	56	386
rect	56	1	57	2
rect	56	4	57	5
rect	56	7	57	8
rect	56	10	57	11
rect	56	13	57	14
rect	56	16	57	17
rect	56	19	57	20
rect	56	22	57	23
rect	56	25	57	26
rect	56	28	57	29
rect	56	31	57	32
rect	56	34	57	35
rect	56	37	57	38
rect	56	40	57	41
rect	56	43	57	44
rect	56	46	57	47
rect	56	49	57	50
rect	56	52	57	53
rect	56	55	57	56
rect	56	58	57	59
rect	56	61	57	62
rect	56	64	57	65
rect	56	67	57	68
rect	56	70	57	71
rect	56	73	57	74
rect	56	76	57	77
rect	56	79	57	80
rect	56	82	57	83
rect	56	85	57	86
rect	56	88	57	89
rect	56	91	57	92
rect	56	94	57	95
rect	56	97	57	98
rect	56	100	57	101
rect	56	103	57	104
rect	56	106	57	107
rect	56	109	57	110
rect	56	112	57	113
rect	56	115	57	116
rect	56	118	57	119
rect	56	121	57	122
rect	56	124	57	125
rect	56	127	57	128
rect	56	130	57	131
rect	56	133	57	134
rect	56	136	57	137
rect	56	139	57	140
rect	56	142	57	143
rect	56	145	57	146
rect	56	148	57	149
rect	56	151	57	152
rect	56	154	57	155
rect	56	157	57	158
rect	56	160	57	161
rect	56	163	57	164
rect	56	166	57	167
rect	56	169	57	170
rect	56	172	57	173
rect	56	175	57	176
rect	56	178	57	179
rect	56	181	57	182
rect	56	184	57	185
rect	56	187	57	188
rect	56	190	57	191
rect	56	193	57	194
rect	56	196	57	197
rect	56	199	57	200
rect	56	202	57	203
rect	56	205	57	206
rect	56	208	57	209
rect	56	211	57	212
rect	56	214	57	215
rect	56	217	57	218
rect	56	220	57	221
rect	56	223	57	224
rect	56	226	57	227
rect	56	229	57	230
rect	56	232	57	233
rect	56	235	57	236
rect	56	238	57	239
rect	56	241	57	242
rect	56	244	57	245
rect	56	247	57	248
rect	56	250	57	251
rect	56	253	57	254
rect	56	256	57	257
rect	56	259	57	260
rect	56	262	57	263
rect	56	265	57	266
rect	56	268	57	269
rect	56	271	57	272
rect	56	274	57	275
rect	56	277	57	278
rect	56	280	57	281
rect	56	283	57	284
rect	56	286	57	287
rect	56	289	57	290
rect	56	292	57	293
rect	56	295	57	296
rect	56	298	57	299
rect	56	301	57	302
rect	56	304	57	305
rect	56	307	57	308
rect	56	310	57	311
rect	56	313	57	314
rect	56	316	57	317
rect	56	319	57	320
rect	56	322	57	323
rect	56	325	57	326
rect	56	328	57	329
rect	56	331	57	332
rect	56	334	57	335
rect	56	337	57	338
rect	56	340	57	341
rect	56	343	57	344
rect	56	346	57	347
rect	56	349	57	350
rect	56	352	57	353
rect	56	355	57	356
rect	56	358	57	359
rect	56	361	57	362
rect	56	364	57	365
rect	56	367	57	368
rect	56	373	57	374
rect	56	376	57	377
rect	56	379	57	380
rect	56	385	57	386
rect	57	1	58	2
rect	57	4	58	5
rect	57	7	58	8
rect	57	10	58	11
rect	57	13	58	14
rect	57	16	58	17
rect	57	19	58	20
rect	57	22	58	23
rect	57	25	58	26
rect	57	28	58	29
rect	57	31	58	32
rect	57	34	58	35
rect	57	37	58	38
rect	57	40	58	41
rect	57	43	58	44
rect	57	46	58	47
rect	57	49	58	50
rect	57	52	58	53
rect	57	55	58	56
rect	57	58	58	59
rect	57	61	58	62
rect	57	64	58	65
rect	57	67	58	68
rect	57	70	58	71
rect	57	73	58	74
rect	57	76	58	77
rect	57	79	58	80
rect	57	82	58	83
rect	57	85	58	86
rect	57	88	58	89
rect	57	91	58	92
rect	57	94	58	95
rect	57	97	58	98
rect	57	100	58	101
rect	57	103	58	104
rect	57	106	58	107
rect	57	109	58	110
rect	57	112	58	113
rect	57	115	58	116
rect	57	118	58	119
rect	57	121	58	122
rect	57	124	58	125
rect	57	127	58	128
rect	57	130	58	131
rect	57	133	58	134
rect	57	136	58	137
rect	57	139	58	140
rect	57	142	58	143
rect	57	145	58	146
rect	57	148	58	149
rect	57	151	58	152
rect	57	154	58	155
rect	57	157	58	158
rect	57	160	58	161
rect	57	163	58	164
rect	57	166	58	167
rect	57	169	58	170
rect	57	172	58	173
rect	57	175	58	176
rect	57	178	58	179
rect	57	181	58	182
rect	57	184	58	185
rect	57	187	58	188
rect	57	190	58	191
rect	57	193	58	194
rect	57	196	58	197
rect	57	199	58	200
rect	57	202	58	203
rect	57	205	58	206
rect	57	208	58	209
rect	57	211	58	212
rect	57	214	58	215
rect	57	217	58	218
rect	57	220	58	221
rect	57	223	58	224
rect	57	226	58	227
rect	57	229	58	230
rect	57	232	58	233
rect	57	235	58	236
rect	57	238	58	239
rect	57	241	58	242
rect	57	244	58	245
rect	57	247	58	248
rect	57	250	58	251
rect	57	253	58	254
rect	57	256	58	257
rect	57	259	58	260
rect	57	262	58	263
rect	57	265	58	266
rect	57	268	58	269
rect	57	271	58	272
rect	57	274	58	275
rect	57	277	58	278
rect	57	280	58	281
rect	57	283	58	284
rect	57	286	58	287
rect	57	289	58	290
rect	57	292	58	293
rect	57	295	58	296
rect	57	298	58	299
rect	57	301	58	302
rect	57	304	58	305
rect	57	307	58	308
rect	57	310	58	311
rect	57	313	58	314
rect	57	316	58	317
rect	57	319	58	320
rect	57	322	58	323
rect	57	325	58	326
rect	57	328	58	329
rect	57	331	58	332
rect	57	334	58	335
rect	57	337	58	338
rect	57	340	58	341
rect	57	343	58	344
rect	57	346	58	347
rect	57	349	58	350
rect	57	352	58	353
rect	57	355	58	356
rect	57	358	58	359
rect	57	361	58	362
rect	57	364	58	365
rect	57	367	58	368
rect	57	373	58	374
rect	57	376	58	377
rect	57	379	58	380
rect	57	385	58	386
rect	58	1	59	2
rect	58	4	59	5
rect	58	7	59	8
rect	58	10	59	11
rect	58	13	59	14
rect	58	16	59	17
rect	58	19	59	20
rect	58	22	59	23
rect	58	25	59	26
rect	58	28	59	29
rect	58	31	59	32
rect	58	34	59	35
rect	58	37	59	38
rect	58	40	59	41
rect	58	43	59	44
rect	58	46	59	47
rect	58	49	59	50
rect	58	52	59	53
rect	58	55	59	56
rect	58	58	59	59
rect	58	61	59	62
rect	58	64	59	65
rect	58	67	59	68
rect	58	70	59	71
rect	58	73	59	74
rect	58	76	59	77
rect	58	79	59	80
rect	58	82	59	83
rect	58	85	59	86
rect	58	88	59	89
rect	58	91	59	92
rect	58	94	59	95
rect	58	97	59	98
rect	58	100	59	101
rect	58	103	59	104
rect	58	106	59	107
rect	58	109	59	110
rect	58	112	59	113
rect	58	115	59	116
rect	58	118	59	119
rect	58	121	59	122
rect	58	124	59	125
rect	58	127	59	128
rect	58	130	59	131
rect	58	133	59	134
rect	58	136	59	137
rect	58	139	59	140
rect	58	142	59	143
rect	58	145	59	146
rect	58	148	59	149
rect	58	151	59	152
rect	58	154	59	155
rect	58	157	59	158
rect	58	160	59	161
rect	58	163	59	164
rect	58	166	59	167
rect	58	169	59	170
rect	58	172	59	173
rect	58	175	59	176
rect	58	178	59	179
rect	58	181	59	182
rect	58	184	59	185
rect	58	187	59	188
rect	58	190	59	191
rect	58	193	59	194
rect	58	196	59	197
rect	58	199	59	200
rect	58	202	59	203
rect	58	205	59	206
rect	58	208	59	209
rect	58	211	59	212
rect	58	214	59	215
rect	58	217	59	218
rect	58	220	59	221
rect	58	223	59	224
rect	58	226	59	227
rect	58	229	59	230
rect	58	232	59	233
rect	58	235	59	236
rect	58	238	59	239
rect	58	241	59	242
rect	58	244	59	245
rect	58	247	59	248
rect	58	250	59	251
rect	58	253	59	254
rect	58	256	59	257
rect	58	259	59	260
rect	58	262	59	263
rect	58	265	59	266
rect	58	268	59	269
rect	58	271	59	272
rect	58	274	59	275
rect	58	277	59	278
rect	58	280	59	281
rect	58	283	59	284
rect	58	286	59	287
rect	58	289	59	290
rect	58	292	59	293
rect	58	295	59	296
rect	58	298	59	299
rect	58	301	59	302
rect	58	304	59	305
rect	58	307	59	308
rect	58	310	59	311
rect	58	313	59	314
rect	58	316	59	317
rect	58	319	59	320
rect	58	322	59	323
rect	58	325	59	326
rect	58	328	59	329
rect	58	331	59	332
rect	58	334	59	335
rect	58	337	59	338
rect	58	340	59	341
rect	58	343	59	344
rect	58	346	59	347
rect	58	349	59	350
rect	58	352	59	353
rect	58	355	59	356
rect	58	358	59	359
rect	58	361	59	362
rect	58	364	59	365
rect	58	367	59	368
rect	58	373	59	374
rect	58	376	59	377
rect	58	379	59	380
rect	58	385	59	386
rect	59	1	60	2
rect	59	4	60	5
rect	59	7	60	8
rect	59	10	60	11
rect	59	13	60	14
rect	59	16	60	17
rect	59	19	60	20
rect	59	22	60	23
rect	59	25	60	26
rect	59	28	60	29
rect	59	31	60	32
rect	59	34	60	35
rect	59	37	60	38
rect	59	40	60	41
rect	59	43	60	44
rect	59	46	60	47
rect	59	49	60	50
rect	59	52	60	53
rect	59	55	60	56
rect	59	58	60	59
rect	59	61	60	62
rect	59	64	60	65
rect	59	67	60	68
rect	59	70	60	71
rect	59	73	60	74
rect	59	76	60	77
rect	59	79	60	80
rect	59	82	60	83
rect	59	85	60	86
rect	59	88	60	89
rect	59	91	60	92
rect	59	94	60	95
rect	59	97	60	98
rect	59	100	60	101
rect	59	103	60	104
rect	59	106	60	107
rect	59	109	60	110
rect	59	112	60	113
rect	59	115	60	116
rect	59	118	60	119
rect	59	121	60	122
rect	59	124	60	125
rect	59	127	60	128
rect	59	130	60	131
rect	59	133	60	134
rect	59	136	60	137
rect	59	139	60	140
rect	59	142	60	143
rect	59	145	60	146
rect	59	148	60	149
rect	59	151	60	152
rect	59	154	60	155
rect	59	157	60	158
rect	59	160	60	161
rect	59	163	60	164
rect	59	166	60	167
rect	59	169	60	170
rect	59	172	60	173
rect	59	175	60	176
rect	59	178	60	179
rect	59	181	60	182
rect	59	184	60	185
rect	59	187	60	188
rect	59	190	60	191
rect	59	193	60	194
rect	59	196	60	197
rect	59	199	60	200
rect	59	202	60	203
rect	59	205	60	206
rect	59	208	60	209
rect	59	211	60	212
rect	59	214	60	215
rect	59	217	60	218
rect	59	220	60	221
rect	59	223	60	224
rect	59	226	60	227
rect	59	229	60	230
rect	59	232	60	233
rect	59	235	60	236
rect	59	238	60	239
rect	59	241	60	242
rect	59	244	60	245
rect	59	247	60	248
rect	59	250	60	251
rect	59	253	60	254
rect	59	256	60	257
rect	59	259	60	260
rect	59	262	60	263
rect	59	265	60	266
rect	59	268	60	269
rect	59	271	60	272
rect	59	274	60	275
rect	59	277	60	278
rect	59	280	60	281
rect	59	283	60	284
rect	59	286	60	287
rect	59	289	60	290
rect	59	292	60	293
rect	59	295	60	296
rect	59	298	60	299
rect	59	301	60	302
rect	59	304	60	305
rect	59	307	60	308
rect	59	310	60	311
rect	59	313	60	314
rect	59	316	60	317
rect	59	319	60	320
rect	59	322	60	323
rect	59	325	60	326
rect	59	328	60	329
rect	59	331	60	332
rect	59	334	60	335
rect	59	337	60	338
rect	59	340	60	341
rect	59	343	60	344
rect	59	346	60	347
rect	59	349	60	350
rect	59	352	60	353
rect	59	355	60	356
rect	59	358	60	359
rect	59	361	60	362
rect	59	364	60	365
rect	59	367	60	368
rect	59	373	60	374
rect	59	376	60	377
rect	59	379	60	380
rect	59	385	60	386
rect	60	1	61	2
rect	60	4	61	5
rect	60	7	61	8
rect	60	10	61	11
rect	60	13	61	14
rect	60	16	61	17
rect	60	19	61	20
rect	60	22	61	23
rect	60	25	61	26
rect	60	28	61	29
rect	60	31	61	32
rect	60	34	61	35
rect	60	37	61	38
rect	60	40	61	41
rect	60	43	61	44
rect	60	46	61	47
rect	60	49	61	50
rect	60	52	61	53
rect	60	55	61	56
rect	60	58	61	59
rect	60	61	61	62
rect	60	64	61	65
rect	60	67	61	68
rect	60	70	61	71
rect	60	73	61	74
rect	60	76	61	77
rect	60	79	61	80
rect	60	82	61	83
rect	60	85	61	86
rect	60	88	61	89
rect	60	91	61	92
rect	60	94	61	95
rect	60	97	61	98
rect	60	100	61	101
rect	60	103	61	104
rect	60	106	61	107
rect	60	109	61	110
rect	60	112	61	113
rect	60	115	61	116
rect	60	118	61	119
rect	60	121	61	122
rect	60	124	61	125
rect	60	127	61	128
rect	60	130	61	131
rect	60	133	61	134
rect	60	136	61	137
rect	60	139	61	140
rect	60	142	61	143
rect	60	145	61	146
rect	60	148	61	149
rect	60	151	61	152
rect	60	154	61	155
rect	60	157	61	158
rect	60	160	61	161
rect	60	163	61	164
rect	60	166	61	167
rect	60	169	61	170
rect	60	172	61	173
rect	60	175	61	176
rect	60	178	61	179
rect	60	181	61	182
rect	60	184	61	185
rect	60	187	61	188
rect	60	190	61	191
rect	60	193	61	194
rect	60	196	61	197
rect	60	199	61	200
rect	60	202	61	203
rect	60	205	61	206
rect	60	208	61	209
rect	60	211	61	212
rect	60	214	61	215
rect	60	217	61	218
rect	60	220	61	221
rect	60	223	61	224
rect	60	226	61	227
rect	60	229	61	230
rect	60	232	61	233
rect	60	235	61	236
rect	60	238	61	239
rect	60	241	61	242
rect	60	244	61	245
rect	60	247	61	248
rect	60	250	61	251
rect	60	253	61	254
rect	60	256	61	257
rect	60	259	61	260
rect	60	262	61	263
rect	60	265	61	266
rect	60	268	61	269
rect	60	271	61	272
rect	60	274	61	275
rect	60	277	61	278
rect	60	280	61	281
rect	60	283	61	284
rect	60	286	61	287
rect	60	289	61	290
rect	60	292	61	293
rect	60	295	61	296
rect	60	298	61	299
rect	60	301	61	302
rect	60	304	61	305
rect	60	307	61	308
rect	60	310	61	311
rect	60	313	61	314
rect	60	316	61	317
rect	60	319	61	320
rect	60	322	61	323
rect	60	325	61	326
rect	60	328	61	329
rect	60	331	61	332
rect	60	334	61	335
rect	60	337	61	338
rect	60	340	61	341
rect	60	343	61	344
rect	60	346	61	347
rect	60	349	61	350
rect	60	352	61	353
rect	60	355	61	356
rect	60	358	61	359
rect	60	361	61	362
rect	60	364	61	365
rect	60	367	61	368
rect	60	373	61	374
rect	60	376	61	377
rect	60	379	61	380
rect	60	385	61	386
rect	61	1	62	2
rect	61	4	62	5
rect	61	7	62	8
rect	61	10	62	11
rect	61	13	62	14
rect	61	16	62	17
rect	61	19	62	20
rect	61	22	62	23
rect	61	25	62	26
rect	61	28	62	29
rect	61	37	62	38
rect	61	40	62	41
rect	61	43	62	44
rect	61	46	62	47
rect	61	49	62	50
rect	61	52	62	53
rect	61	55	62	56
rect	61	58	62	59
rect	61	61	62	62
rect	61	64	62	65
rect	61	67	62	68
rect	61	70	62	71
rect	61	73	62	74
rect	61	76	62	77
rect	61	79	62	80
rect	61	82	62	83
rect	61	85	62	86
rect	61	88	62	89
rect	61	91	62	92
rect	61	94	62	95
rect	61	97	62	98
rect	61	100	62	101
rect	61	103	62	104
rect	61	106	62	107
rect	61	109	62	110
rect	61	112	62	113
rect	61	115	62	116
rect	61	118	62	119
rect	61	121	62	122
rect	61	124	62	125
rect	61	127	62	128
rect	61	130	62	131
rect	61	133	62	134
rect	61	136	62	137
rect	61	139	62	140
rect	61	142	62	143
rect	61	145	62	146
rect	61	148	62	149
rect	61	151	62	152
rect	61	154	62	155
rect	61	157	62	158
rect	61	160	62	161
rect	61	163	62	164
rect	61	166	62	167
rect	61	169	62	170
rect	61	172	62	173
rect	61	175	62	176
rect	61	178	62	179
rect	61	181	62	182
rect	61	184	62	185
rect	61	187	62	188
rect	61	190	62	191
rect	61	193	62	194
rect	61	196	62	197
rect	61	199	62	200
rect	61	202	62	203
rect	61	205	62	206
rect	61	208	62	209
rect	61	211	62	212
rect	61	214	62	215
rect	61	217	62	218
rect	61	220	62	221
rect	61	223	62	224
rect	61	226	62	227
rect	61	229	62	230
rect	61	232	62	233
rect	61	235	62	236
rect	61	238	62	239
rect	61	241	62	242
rect	61	244	62	245
rect	61	247	62	248
rect	61	250	62	251
rect	61	253	62	254
rect	61	256	62	257
rect	61	259	62	260
rect	61	262	62	263
rect	61	265	62	266
rect	61	268	62	269
rect	61	271	62	272
rect	61	274	62	275
rect	61	277	62	278
rect	61	280	62	281
rect	61	283	62	284
rect	61	286	62	287
rect	61	289	62	290
rect	61	292	62	293
rect	61	295	62	296
rect	61	298	62	299
rect	61	301	62	302
rect	61	304	62	305
rect	61	307	62	308
rect	61	310	62	311
rect	61	313	62	314
rect	61	316	62	317
rect	61	319	62	320
rect	61	322	62	323
rect	61	325	62	326
rect	61	328	62	329
rect	61	331	62	332
rect	61	334	62	335
rect	61	337	62	338
rect	61	340	62	341
rect	61	343	62	344
rect	61	346	62	347
rect	61	349	62	350
rect	61	352	62	353
rect	61	355	62	356
rect	61	358	62	359
rect	61	361	62	362
rect	61	364	62	365
rect	61	367	62	368
rect	61	373	62	374
rect	61	376	62	377
rect	61	379	62	380
rect	61	385	62	386
rect	62	1	63	2
rect	62	4	63	5
rect	62	7	63	8
rect	62	10	63	11
rect	62	13	63	14
rect	62	16	63	17
rect	62	19	63	20
rect	62	22	63	23
rect	62	25	63	26
rect	62	28	63	29
rect	62	31	63	32
rect	62	34	63	35
rect	62	37	63	38
rect	62	40	63	41
rect	62	43	63	44
rect	62	46	63	47
rect	62	49	63	50
rect	62	52	63	53
rect	62	55	63	56
rect	62	58	63	59
rect	62	61	63	62
rect	62	64	63	65
rect	62	67	63	68
rect	62	70	63	71
rect	62	73	63	74
rect	62	76	63	77
rect	62	79	63	80
rect	62	82	63	83
rect	62	85	63	86
rect	62	88	63	89
rect	62	91	63	92
rect	62	94	63	95
rect	62	97	63	98
rect	62	100	63	101
rect	62	103	63	104
rect	62	106	63	107
rect	62	109	63	110
rect	62	112	63	113
rect	62	115	63	116
rect	62	118	63	119
rect	62	121	63	122
rect	62	124	63	125
rect	62	127	63	128
rect	62	130	63	131
rect	62	133	63	134
rect	62	136	63	137
rect	62	139	63	140
rect	62	142	63	143
rect	62	145	63	146
rect	62	148	63	149
rect	62	151	63	152
rect	62	154	63	155
rect	62	157	63	158
rect	62	160	63	161
rect	62	163	63	164
rect	62	166	63	167
rect	62	169	63	170
rect	62	172	63	173
rect	62	175	63	176
rect	62	178	63	179
rect	62	181	63	182
rect	62	184	63	185
rect	62	187	63	188
rect	62	190	63	191
rect	62	193	63	194
rect	62	196	63	197
rect	62	199	63	200
rect	62	202	63	203
rect	62	205	63	206
rect	62	208	63	209
rect	62	211	63	212
rect	62	214	63	215
rect	62	217	63	218
rect	62	220	63	221
rect	62	223	63	224
rect	62	226	63	227
rect	62	229	63	230
rect	62	232	63	233
rect	62	235	63	236
rect	62	238	63	239
rect	62	241	63	242
rect	62	244	63	245
rect	62	247	63	248
rect	62	250	63	251
rect	62	253	63	254
rect	62	256	63	257
rect	62	259	63	260
rect	62	262	63	263
rect	62	265	63	266
rect	62	268	63	269
rect	62	271	63	272
rect	62	274	63	275
rect	62	277	63	278
rect	62	280	63	281
rect	62	283	63	284
rect	62	286	63	287
rect	62	289	63	290
rect	62	292	63	293
rect	62	295	63	296
rect	62	298	63	299
rect	62	301	63	302
rect	62	304	63	305
rect	62	307	63	308
rect	62	310	63	311
rect	62	313	63	314
rect	62	316	63	317
rect	62	319	63	320
rect	62	322	63	323
rect	62	325	63	326
rect	62	328	63	329
rect	62	331	63	332
rect	62	334	63	335
rect	62	337	63	338
rect	62	340	63	341
rect	62	343	63	344
rect	62	346	63	347
rect	62	349	63	350
rect	62	352	63	353
rect	62	355	63	356
rect	62	358	63	359
rect	62	361	63	362
rect	62	364	63	365
rect	62	367	63	368
rect	62	373	63	374
rect	62	376	63	377
rect	62	379	63	380
rect	62	385	63	386
rect	63	1	64	2
rect	63	4	64	5
rect	63	7	64	8
rect	63	10	64	11
rect	63	13	64	14
rect	63	16	64	17
rect	63	19	64	20
rect	63	22	64	23
rect	63	25	64	26
rect	63	28	64	29
rect	63	31	64	32
rect	63	34	64	35
rect	63	37	64	38
rect	63	40	64	41
rect	63	43	64	44
rect	63	46	64	47
rect	63	49	64	50
rect	63	52	64	53
rect	63	55	64	56
rect	63	58	64	59
rect	63	61	64	62
rect	63	64	64	65
rect	63	67	64	68
rect	63	70	64	71
rect	63	73	64	74
rect	63	76	64	77
rect	63	79	64	80
rect	63	82	64	83
rect	63	85	64	86
rect	63	88	64	89
rect	63	91	64	92
rect	63	94	64	95
rect	63	97	64	98
rect	63	100	64	101
rect	63	103	64	104
rect	63	106	64	107
rect	63	109	64	110
rect	63	112	64	113
rect	63	115	64	116
rect	63	118	64	119
rect	63	121	64	122
rect	63	124	64	125
rect	63	127	64	128
rect	63	130	64	131
rect	63	133	64	134
rect	63	136	64	137
rect	63	139	64	140
rect	63	142	64	143
rect	63	145	64	146
rect	63	148	64	149
rect	63	151	64	152
rect	63	154	64	155
rect	63	157	64	158
rect	63	160	64	161
rect	63	163	64	164
rect	63	166	64	167
rect	63	169	64	170
rect	63	172	64	173
rect	63	175	64	176
rect	63	178	64	179
rect	63	181	64	182
rect	63	184	64	185
rect	63	187	64	188
rect	63	190	64	191
rect	63	193	64	194
rect	63	196	64	197
rect	63	199	64	200
rect	63	202	64	203
rect	63	205	64	206
rect	63	208	64	209
rect	63	211	64	212
rect	63	214	64	215
rect	63	217	64	218
rect	63	220	64	221
rect	63	223	64	224
rect	63	226	64	227
rect	63	229	64	230
rect	63	232	64	233
rect	63	235	64	236
rect	63	238	64	239
rect	63	241	64	242
rect	63	244	64	245
rect	63	247	64	248
rect	63	250	64	251
rect	63	253	64	254
rect	63	256	64	257
rect	63	259	64	260
rect	63	262	64	263
rect	63	265	64	266
rect	63	268	64	269
rect	63	271	64	272
rect	63	274	64	275
rect	63	277	64	278
rect	63	280	64	281
rect	63	283	64	284
rect	63	286	64	287
rect	63	289	64	290
rect	63	292	64	293
rect	63	295	64	296
rect	63	298	64	299
rect	63	301	64	302
rect	63	304	64	305
rect	63	307	64	308
rect	63	310	64	311
rect	63	313	64	314
rect	63	316	64	317
rect	63	319	64	320
rect	63	322	64	323
rect	63	325	64	326
rect	63	328	64	329
rect	63	331	64	332
rect	63	334	64	335
rect	63	337	64	338
rect	63	340	64	341
rect	63	343	64	344
rect	63	346	64	347
rect	63	349	64	350
rect	63	352	64	353
rect	63	355	64	356
rect	63	358	64	359
rect	63	361	64	362
rect	63	364	64	365
rect	63	367	64	368
rect	63	373	64	374
rect	63	376	64	377
rect	63	379	64	380
rect	63	385	64	386
rect	64	1	65	2
rect	64	4	65	5
rect	64	7	65	8
rect	64	10	65	11
rect	64	13	65	14
rect	64	16	65	17
rect	64	19	65	20
rect	64	22	65	23
rect	64	25	65	26
rect	64	28	65	29
rect	64	31	65	32
rect	64	34	65	35
rect	64	37	65	38
rect	64	40	65	41
rect	64	43	65	44
rect	64	46	65	47
rect	64	49	65	50
rect	64	52	65	53
rect	64	55	65	56
rect	64	58	65	59
rect	64	61	65	62
rect	64	64	65	65
rect	64	67	65	68
rect	64	70	65	71
rect	64	73	65	74
rect	64	76	65	77
rect	64	79	65	80
rect	64	82	65	83
rect	64	85	65	86
rect	64	88	65	89
rect	64	91	65	92
rect	64	94	65	95
rect	64	97	65	98
rect	64	100	65	101
rect	64	103	65	104
rect	64	106	65	107
rect	64	109	65	110
rect	64	112	65	113
rect	64	115	65	116
rect	64	118	65	119
rect	64	121	65	122
rect	64	124	65	125
rect	64	127	65	128
rect	64	130	65	131
rect	64	133	65	134
rect	64	136	65	137
rect	64	139	65	140
rect	64	142	65	143
rect	64	145	65	146
rect	64	148	65	149
rect	64	151	65	152
rect	64	154	65	155
rect	64	157	65	158
rect	64	160	65	161
rect	64	163	65	164
rect	64	166	65	167
rect	64	169	65	170
rect	64	172	65	173
rect	64	175	65	176
rect	64	178	65	179
rect	64	181	65	182
rect	64	184	65	185
rect	64	187	65	188
rect	64	190	65	191
rect	64	193	65	194
rect	64	196	65	197
rect	64	199	65	200
rect	64	202	65	203
rect	64	205	65	206
rect	64	208	65	209
rect	64	211	65	212
rect	64	214	65	215
rect	64	217	65	218
rect	64	220	65	221
rect	64	223	65	224
rect	64	226	65	227
rect	64	229	65	230
rect	64	232	65	233
rect	64	235	65	236
rect	64	238	65	239
rect	64	241	65	242
rect	64	244	65	245
rect	64	247	65	248
rect	64	250	65	251
rect	64	253	65	254
rect	64	256	65	257
rect	64	259	65	260
rect	64	262	65	263
rect	64	265	65	266
rect	64	268	65	269
rect	64	271	65	272
rect	64	274	65	275
rect	64	277	65	278
rect	64	280	65	281
rect	64	283	65	284
rect	64	286	65	287
rect	64	289	65	290
rect	64	292	65	293
rect	64	295	65	296
rect	64	298	65	299
rect	64	301	65	302
rect	64	304	65	305
rect	64	307	65	308
rect	64	310	65	311
rect	64	313	65	314
rect	64	316	65	317
rect	64	319	65	320
rect	64	322	65	323
rect	64	325	65	326
rect	64	328	65	329
rect	64	331	65	332
rect	64	334	65	335
rect	64	337	65	338
rect	64	340	65	341
rect	64	343	65	344
rect	64	346	65	347
rect	64	349	65	350
rect	64	352	65	353
rect	64	355	65	356
rect	64	358	65	359
rect	64	361	65	362
rect	64	364	65	365
rect	64	367	65	368
rect	64	373	65	374
rect	64	376	65	377
rect	64	379	65	380
rect	64	385	65	386
rect	65	1	66	2
rect	65	4	66	5
rect	65	7	66	8
rect	65	10	66	11
rect	65	13	66	14
rect	65	16	66	17
rect	65	19	66	20
rect	65	22	66	23
rect	65	25	66	26
rect	65	28	66	29
rect	65	31	66	32
rect	65	34	66	35
rect	65	37	66	38
rect	65	40	66	41
rect	65	43	66	44
rect	65	46	66	47
rect	65	49	66	50
rect	65	52	66	53
rect	65	55	66	56
rect	65	58	66	59
rect	65	61	66	62
rect	65	64	66	65
rect	65	67	66	68
rect	65	70	66	71
rect	65	73	66	74
rect	65	76	66	77
rect	65	79	66	80
rect	65	82	66	83
rect	65	85	66	86
rect	65	88	66	89
rect	65	91	66	92
rect	65	94	66	95
rect	65	97	66	98
rect	65	100	66	101
rect	65	103	66	104
rect	65	106	66	107
rect	65	109	66	110
rect	65	112	66	113
rect	65	115	66	116
rect	65	118	66	119
rect	65	121	66	122
rect	65	124	66	125
rect	65	127	66	128
rect	65	130	66	131
rect	65	133	66	134
rect	65	136	66	137
rect	65	139	66	140
rect	65	142	66	143
rect	65	145	66	146
rect	65	148	66	149
rect	65	151	66	152
rect	65	154	66	155
rect	65	157	66	158
rect	65	160	66	161
rect	65	163	66	164
rect	65	166	66	167
rect	65	169	66	170
rect	65	172	66	173
rect	65	175	66	176
rect	65	178	66	179
rect	65	181	66	182
rect	65	184	66	185
rect	65	187	66	188
rect	65	190	66	191
rect	65	193	66	194
rect	65	196	66	197
rect	65	199	66	200
rect	65	202	66	203
rect	65	205	66	206
rect	65	208	66	209
rect	65	211	66	212
rect	65	214	66	215
rect	65	217	66	218
rect	65	220	66	221
rect	65	223	66	224
rect	65	226	66	227
rect	65	229	66	230
rect	65	232	66	233
rect	65	235	66	236
rect	65	238	66	239
rect	65	241	66	242
rect	65	244	66	245
rect	65	247	66	248
rect	65	250	66	251
rect	65	253	66	254
rect	65	256	66	257
rect	65	259	66	260
rect	65	262	66	263
rect	65	265	66	266
rect	65	268	66	269
rect	65	271	66	272
rect	65	274	66	275
rect	65	277	66	278
rect	65	280	66	281
rect	65	283	66	284
rect	65	286	66	287
rect	65	289	66	290
rect	65	292	66	293
rect	65	295	66	296
rect	65	298	66	299
rect	65	301	66	302
rect	65	304	66	305
rect	65	307	66	308
rect	65	310	66	311
rect	65	313	66	314
rect	65	316	66	317
rect	65	319	66	320
rect	65	322	66	323
rect	65	325	66	326
rect	65	328	66	329
rect	65	331	66	332
rect	65	334	66	335
rect	65	337	66	338
rect	65	340	66	341
rect	65	343	66	344
rect	65	346	66	347
rect	65	349	66	350
rect	65	352	66	353
rect	65	355	66	356
rect	65	358	66	359
rect	65	361	66	362
rect	65	364	66	365
rect	65	367	66	368
rect	65	373	66	374
rect	65	376	66	377
rect	65	379	66	380
rect	65	385	66	386
rect	66	1	67	2
rect	66	4	67	5
rect	66	7	67	8
rect	66	10	67	11
rect	66	13	67	14
rect	66	16	67	17
rect	66	19	67	20
rect	66	22	67	23
rect	66	25	67	26
rect	66	28	67	29
rect	66	31	67	32
rect	66	34	67	35
rect	66	37	67	38
rect	66	40	67	41
rect	66	43	67	44
rect	66	46	67	47
rect	66	49	67	50
rect	66	52	67	53
rect	66	55	67	56
rect	66	58	67	59
rect	66	61	67	62
rect	66	64	67	65
rect	66	67	67	68
rect	66	70	67	71
rect	66	73	67	74
rect	66	76	67	77
rect	66	79	67	80
rect	66	82	67	83
rect	66	85	67	86
rect	66	88	67	89
rect	66	91	67	92
rect	66	94	67	95
rect	66	97	67	98
rect	66	100	67	101
rect	66	103	67	104
rect	66	106	67	107
rect	66	109	67	110
rect	66	112	67	113
rect	66	115	67	116
rect	66	118	67	119
rect	66	121	67	122
rect	66	124	67	125
rect	66	127	67	128
rect	66	130	67	131
rect	66	133	67	134
rect	66	136	67	137
rect	66	139	67	140
rect	66	142	67	143
rect	66	145	67	146
rect	66	148	67	149
rect	66	151	67	152
rect	66	154	67	155
rect	66	157	67	158
rect	66	160	67	161
rect	66	163	67	164
rect	66	166	67	167
rect	66	169	67	170
rect	66	172	67	173
rect	66	175	67	176
rect	66	178	67	179
rect	66	181	67	182
rect	66	184	67	185
rect	66	187	67	188
rect	66	190	67	191
rect	66	193	67	194
rect	66	196	67	197
rect	66	199	67	200
rect	66	202	67	203
rect	66	205	67	206
rect	66	208	67	209
rect	66	211	67	212
rect	66	214	67	215
rect	66	217	67	218
rect	66	220	67	221
rect	66	223	67	224
rect	66	226	67	227
rect	66	229	67	230
rect	66	232	67	233
rect	66	235	67	236
rect	66	238	67	239
rect	66	241	67	242
rect	66	244	67	245
rect	66	247	67	248
rect	66	250	67	251
rect	66	253	67	254
rect	66	256	67	257
rect	66	259	67	260
rect	66	262	67	263
rect	66	265	67	266
rect	66	268	67	269
rect	66	271	67	272
rect	66	274	67	275
rect	66	277	67	278
rect	66	280	67	281
rect	66	283	67	284
rect	66	286	67	287
rect	66	289	67	290
rect	66	292	67	293
rect	66	295	67	296
rect	66	298	67	299
rect	66	301	67	302
rect	66	304	67	305
rect	66	307	67	308
rect	66	310	67	311
rect	66	313	67	314
rect	66	316	67	317
rect	66	319	67	320
rect	66	322	67	323
rect	66	325	67	326
rect	66	328	67	329
rect	66	331	67	332
rect	66	334	67	335
rect	66	337	67	338
rect	66	340	67	341
rect	66	343	67	344
rect	66	346	67	347
rect	66	349	67	350
rect	66	352	67	353
rect	66	355	67	356
rect	66	358	67	359
rect	66	361	67	362
rect	66	364	67	365
rect	66	367	67	368
rect	66	373	67	374
rect	66	376	67	377
rect	66	379	67	380
rect	66	385	67	386
rect	67	1	68	2
rect	67	4	68	5
rect	67	7	68	8
rect	67	10	68	11
rect	67	13	68	14
rect	67	16	68	17
rect	67	19	68	20
rect	67	22	68	23
rect	67	25	68	26
rect	67	28	68	29
rect	67	31	68	32
rect	67	34	68	35
rect	67	37	68	38
rect	67	40	68	41
rect	67	43	68	44
rect	67	46	68	47
rect	67	49	68	50
rect	67	52	68	53
rect	67	55	68	56
rect	67	58	68	59
rect	67	61	68	62
rect	67	64	68	65
rect	67	67	68	68
rect	67	70	68	71
rect	67	73	68	74
rect	67	76	68	77
rect	67	79	68	80
rect	67	82	68	83
rect	67	85	68	86
rect	67	88	68	89
rect	67	91	68	92
rect	67	94	68	95
rect	67	97	68	98
rect	67	100	68	101
rect	67	103	68	104
rect	67	106	68	107
rect	67	109	68	110
rect	67	112	68	113
rect	67	115	68	116
rect	67	118	68	119
rect	67	121	68	122
rect	67	124	68	125
rect	67	127	68	128
rect	67	130	68	131
rect	67	133	68	134
rect	67	136	68	137
rect	67	139	68	140
rect	67	142	68	143
rect	67	145	68	146
rect	67	148	68	149
rect	67	151	68	152
rect	67	154	68	155
rect	67	157	68	158
rect	67	160	68	161
rect	67	163	68	164
rect	67	166	68	167
rect	67	169	68	170
rect	67	172	68	173
rect	67	175	68	176
rect	67	178	68	179
rect	67	181	68	182
rect	67	184	68	185
rect	67	187	68	188
rect	67	190	68	191
rect	67	193	68	194
rect	67	196	68	197
rect	67	199	68	200
rect	67	202	68	203
rect	67	205	68	206
rect	67	208	68	209
rect	67	211	68	212
rect	67	214	68	215
rect	67	217	68	218
rect	67	220	68	221
rect	67	223	68	224
rect	67	226	68	227
rect	67	229	68	230
rect	67	232	68	233
rect	67	235	68	236
rect	67	238	68	239
rect	67	241	68	242
rect	67	244	68	245
rect	67	247	68	248
rect	67	250	68	251
rect	67	253	68	254
rect	67	256	68	257
rect	67	259	68	260
rect	67	262	68	263
rect	67	265	68	266
rect	67	268	68	269
rect	67	271	68	272
rect	67	274	68	275
rect	67	277	68	278
rect	67	280	68	281
rect	67	283	68	284
rect	67	286	68	287
rect	67	289	68	290
rect	67	292	68	293
rect	67	295	68	296
rect	67	298	68	299
rect	67	301	68	302
rect	67	304	68	305
rect	67	307	68	308
rect	67	310	68	311
rect	67	313	68	314
rect	67	316	68	317
rect	67	319	68	320
rect	67	322	68	323
rect	67	325	68	326
rect	67	328	68	329
rect	67	331	68	332
rect	67	334	68	335
rect	67	337	68	338
rect	67	340	68	341
rect	67	343	68	344
rect	67	346	68	347
rect	67	349	68	350
rect	67	352	68	353
rect	67	355	68	356
rect	67	358	68	359
rect	67	361	68	362
rect	67	364	68	365
rect	67	367	68	368
rect	67	373	68	374
rect	67	376	68	377
rect	67	379	68	380
rect	67	385	68	386
rect	68	1	69	2
rect	68	4	69	5
rect	68	7	69	8
rect	68	10	69	11
rect	68	13	69	14
rect	68	16	69	17
rect	68	19	69	20
rect	68	22	69	23
rect	68	25	69	26
rect	68	28	69	29
rect	68	31	69	32
rect	68	34	69	35
rect	68	37	69	38
rect	68	40	69	41
rect	68	43	69	44
rect	68	46	69	47
rect	68	49	69	50
rect	68	52	69	53
rect	68	55	69	56
rect	68	58	69	59
rect	68	61	69	62
rect	68	64	69	65
rect	68	67	69	68
rect	68	70	69	71
rect	68	73	69	74
rect	68	76	69	77
rect	68	79	69	80
rect	68	82	69	83
rect	68	85	69	86
rect	68	88	69	89
rect	68	91	69	92
rect	68	94	69	95
rect	68	97	69	98
rect	68	100	69	101
rect	68	103	69	104
rect	68	106	69	107
rect	68	109	69	110
rect	68	112	69	113
rect	68	115	69	116
rect	68	118	69	119
rect	68	121	69	122
rect	68	124	69	125
rect	68	127	69	128
rect	68	130	69	131
rect	68	133	69	134
rect	68	136	69	137
rect	68	139	69	140
rect	68	142	69	143
rect	68	145	69	146
rect	68	148	69	149
rect	68	151	69	152
rect	68	154	69	155
rect	68	157	69	158
rect	68	160	69	161
rect	68	163	69	164
rect	68	166	69	167
rect	68	169	69	170
rect	68	172	69	173
rect	68	175	69	176
rect	68	178	69	179
rect	68	181	69	182
rect	68	184	69	185
rect	68	187	69	188
rect	68	190	69	191
rect	68	193	69	194
rect	68	196	69	197
rect	68	199	69	200
rect	68	202	69	203
rect	68	205	69	206
rect	68	208	69	209
rect	68	211	69	212
rect	68	214	69	215
rect	68	217	69	218
rect	68	220	69	221
rect	68	223	69	224
rect	68	226	69	227
rect	68	229	69	230
rect	68	232	69	233
rect	68	235	69	236
rect	68	238	69	239
rect	68	241	69	242
rect	68	244	69	245
rect	68	247	69	248
rect	68	250	69	251
rect	68	253	69	254
rect	68	256	69	257
rect	68	259	69	260
rect	68	262	69	263
rect	68	265	69	266
rect	68	268	69	269
rect	68	271	69	272
rect	68	274	69	275
rect	68	277	69	278
rect	68	280	69	281
rect	68	283	69	284
rect	68	286	69	287
rect	68	289	69	290
rect	68	292	69	293
rect	68	295	69	296
rect	68	298	69	299
rect	68	301	69	302
rect	68	304	69	305
rect	68	307	69	308
rect	68	310	69	311
rect	68	313	69	314
rect	68	316	69	317
rect	68	319	69	320
rect	68	322	69	323
rect	68	325	69	326
rect	68	328	69	329
rect	68	331	69	332
rect	68	334	69	335
rect	68	337	69	338
rect	68	340	69	341
rect	68	343	69	344
rect	68	346	69	347
rect	68	349	69	350
rect	68	352	69	353
rect	68	355	69	356
rect	68	358	69	359
rect	68	361	69	362
rect	68	364	69	365
rect	68	367	69	368
rect	68	373	69	374
rect	68	376	69	377
rect	68	379	69	380
rect	68	385	69	386
rect	69	1	70	2
rect	69	4	70	5
rect	69	7	70	8
rect	69	10	70	11
rect	69	13	70	14
rect	69	16	70	17
rect	69	19	70	20
rect	69	22	70	23
rect	69	25	70	26
rect	69	28	70	29
rect	69	31	70	32
rect	69	34	70	35
rect	69	37	70	38
rect	69	40	70	41
rect	69	43	70	44
rect	69	46	70	47
rect	69	49	70	50
rect	69	52	70	53
rect	69	55	70	56
rect	69	58	70	59
rect	69	61	70	62
rect	69	64	70	65
rect	69	67	70	68
rect	69	70	70	71
rect	69	73	70	74
rect	69	76	70	77
rect	69	79	70	80
rect	69	82	70	83
rect	69	85	70	86
rect	69	88	70	89
rect	69	91	70	92
rect	69	94	70	95
rect	69	97	70	98
rect	69	100	70	101
rect	69	103	70	104
rect	69	106	70	107
rect	69	109	70	110
rect	69	112	70	113
rect	69	115	70	116
rect	69	118	70	119
rect	69	121	70	122
rect	69	124	70	125
rect	69	127	70	128
rect	69	130	70	131
rect	69	133	70	134
rect	69	136	70	137
rect	69	139	70	140
rect	69	142	70	143
rect	69	145	70	146
rect	69	148	70	149
rect	69	151	70	152
rect	69	154	70	155
rect	69	157	70	158
rect	69	160	70	161
rect	69	163	70	164
rect	69	166	70	167
rect	69	169	70	170
rect	69	172	70	173
rect	69	175	70	176
rect	69	178	70	179
rect	69	181	70	182
rect	69	184	70	185
rect	69	187	70	188
rect	69	190	70	191
rect	69	193	70	194
rect	69	196	70	197
rect	69	199	70	200
rect	69	202	70	203
rect	69	205	70	206
rect	69	208	70	209
rect	69	211	70	212
rect	69	214	70	215
rect	69	217	70	218
rect	69	220	70	221
rect	69	223	70	224
rect	69	226	70	227
rect	69	229	70	230
rect	69	232	70	233
rect	69	235	70	236
rect	69	238	70	239
rect	69	241	70	242
rect	69	244	70	245
rect	69	247	70	248
rect	69	250	70	251
rect	69	253	70	254
rect	69	256	70	257
rect	69	259	70	260
rect	69	262	70	263
rect	69	265	70	266
rect	69	268	70	269
rect	69	271	70	272
rect	69	274	70	275
rect	69	277	70	278
rect	69	280	70	281
rect	69	283	70	284
rect	69	286	70	287
rect	69	289	70	290
rect	69	292	70	293
rect	69	295	70	296
rect	69	298	70	299
rect	69	301	70	302
rect	69	304	70	305
rect	69	307	70	308
rect	69	310	70	311
rect	69	313	70	314
rect	69	316	70	317
rect	69	319	70	320
rect	69	322	70	323
rect	69	325	70	326
rect	69	328	70	329
rect	69	331	70	332
rect	69	334	70	335
rect	69	337	70	338
rect	69	340	70	341
rect	69	343	70	344
rect	69	346	70	347
rect	69	349	70	350
rect	69	352	70	353
rect	69	355	70	356
rect	69	358	70	359
rect	69	361	70	362
rect	69	364	70	365
rect	69	367	70	368
rect	69	373	70	374
rect	69	376	70	377
rect	69	379	70	380
rect	69	385	70	386
rect	70	1	71	2
rect	70	4	71	5
rect	70	7	71	8
rect	70	10	71	11
rect	70	13	71	14
rect	70	16	71	17
rect	70	19	71	20
rect	70	22	71	23
rect	70	25	71	26
rect	70	28	71	29
rect	70	31	71	32
rect	70	34	71	35
rect	70	37	71	38
rect	70	40	71	41
rect	70	43	71	44
rect	70	46	71	47
rect	70	49	71	50
rect	70	52	71	53
rect	70	55	71	56
rect	70	58	71	59
rect	70	61	71	62
rect	70	64	71	65
rect	70	67	71	68
rect	70	70	71	71
rect	70	73	71	74
rect	70	76	71	77
rect	70	79	71	80
rect	70	82	71	83
rect	70	85	71	86
rect	70	88	71	89
rect	70	91	71	92
rect	70	94	71	95
rect	70	97	71	98
rect	70	100	71	101
rect	70	103	71	104
rect	70	106	71	107
rect	70	109	71	110
rect	70	112	71	113
rect	70	115	71	116
rect	70	118	71	119
rect	70	121	71	122
rect	70	124	71	125
rect	70	127	71	128
rect	70	130	71	131
rect	70	133	71	134
rect	70	136	71	137
rect	70	139	71	140
rect	70	142	71	143
rect	70	145	71	146
rect	70	148	71	149
rect	70	151	71	152
rect	70	154	71	155
rect	70	157	71	158
rect	70	160	71	161
rect	70	163	71	164
rect	70	166	71	167
rect	70	169	71	170
rect	70	172	71	173
rect	70	175	71	176
rect	70	178	71	179
rect	70	181	71	182
rect	70	184	71	185
rect	70	187	71	188
rect	70	190	71	191
rect	70	193	71	194
rect	70	196	71	197
rect	70	199	71	200
rect	70	202	71	203
rect	70	205	71	206
rect	70	208	71	209
rect	70	211	71	212
rect	70	214	71	215
rect	70	217	71	218
rect	70	220	71	221
rect	70	223	71	224
rect	70	226	71	227
rect	70	229	71	230
rect	70	232	71	233
rect	70	235	71	236
rect	70	238	71	239
rect	70	241	71	242
rect	70	244	71	245
rect	70	247	71	248
rect	70	250	71	251
rect	70	253	71	254
rect	70	256	71	257
rect	70	259	71	260
rect	70	262	71	263
rect	70	265	71	266
rect	70	268	71	269
rect	70	271	71	272
rect	70	274	71	275
rect	70	277	71	278
rect	70	280	71	281
rect	70	283	71	284
rect	70	286	71	287
rect	70	289	71	290
rect	70	292	71	293
rect	70	295	71	296
rect	70	298	71	299
rect	70	301	71	302
rect	70	304	71	305
rect	70	307	71	308
rect	70	310	71	311
rect	70	313	71	314
rect	70	316	71	317
rect	70	319	71	320
rect	70	322	71	323
rect	70	325	71	326
rect	70	328	71	329
rect	70	331	71	332
rect	70	334	71	335
rect	70	337	71	338
rect	70	340	71	341
rect	70	343	71	344
rect	70	346	71	347
rect	70	349	71	350
rect	70	352	71	353
rect	70	355	71	356
rect	70	358	71	359
rect	70	361	71	362
rect	70	364	71	365
rect	70	367	71	368
rect	70	373	71	374
rect	70	376	71	377
rect	70	379	71	380
rect	70	385	71	386
rect	71	1	72	2
rect	71	4	72	5
rect	71	7	72	8
rect	71	10	72	11
rect	71	13	72	14
rect	71	16	72	17
rect	71	19	72	20
rect	71	22	72	23
rect	71	25	72	26
rect	71	28	72	29
rect	71	31	72	32
rect	71	34	72	35
rect	71	37	72	38
rect	71	40	72	41
rect	71	43	72	44
rect	71	46	72	47
rect	71	49	72	50
rect	71	52	72	53
rect	71	55	72	56
rect	71	58	72	59
rect	71	61	72	62
rect	71	64	72	65
rect	71	67	72	68
rect	71	70	72	71
rect	71	73	72	74
rect	71	76	72	77
rect	71	79	72	80
rect	71	82	72	83
rect	71	85	72	86
rect	71	88	72	89
rect	71	91	72	92
rect	71	94	72	95
rect	71	97	72	98
rect	71	100	72	101
rect	71	103	72	104
rect	71	106	72	107
rect	71	109	72	110
rect	71	112	72	113
rect	71	115	72	116
rect	71	118	72	119
rect	71	121	72	122
rect	71	124	72	125
rect	71	127	72	128
rect	71	130	72	131
rect	71	133	72	134
rect	71	136	72	137
rect	71	139	72	140
rect	71	142	72	143
rect	71	145	72	146
rect	71	148	72	149
rect	71	151	72	152
rect	71	154	72	155
rect	71	157	72	158
rect	71	160	72	161
rect	71	163	72	164
rect	71	166	72	167
rect	71	169	72	170
rect	71	172	72	173
rect	71	175	72	176
rect	71	178	72	179
rect	71	181	72	182
rect	71	184	72	185
rect	71	187	72	188
rect	71	190	72	191
rect	71	193	72	194
rect	71	196	72	197
rect	71	199	72	200
rect	71	202	72	203
rect	71	205	72	206
rect	71	208	72	209
rect	71	211	72	212
rect	71	214	72	215
rect	71	217	72	218
rect	71	220	72	221
rect	71	223	72	224
rect	71	226	72	227
rect	71	229	72	230
rect	71	232	72	233
rect	71	235	72	236
rect	71	238	72	239
rect	71	241	72	242
rect	71	244	72	245
rect	71	247	72	248
rect	71	250	72	251
rect	71	253	72	254
rect	71	256	72	257
rect	71	259	72	260
rect	71	262	72	263
rect	71	265	72	266
rect	71	268	72	269
rect	71	271	72	272
rect	71	274	72	275
rect	71	277	72	278
rect	71	280	72	281
rect	71	283	72	284
rect	71	286	72	287
rect	71	289	72	290
rect	71	292	72	293
rect	71	295	72	296
rect	71	298	72	299
rect	71	301	72	302
rect	71	304	72	305
rect	71	307	72	308
rect	71	310	72	311
rect	71	313	72	314
rect	71	316	72	317
rect	71	319	72	320
rect	71	322	72	323
rect	71	325	72	326
rect	71	328	72	329
rect	71	331	72	332
rect	71	334	72	335
rect	71	337	72	338
rect	71	340	72	341
rect	71	343	72	344
rect	71	346	72	347
rect	71	349	72	350
rect	71	352	72	353
rect	71	355	72	356
rect	71	358	72	359
rect	71	361	72	362
rect	71	364	72	365
rect	71	367	72	368
rect	71	373	72	374
rect	71	376	72	377
rect	71	379	72	380
rect	71	385	72	386
rect	72	1	73	2
rect	72	4	73	5
rect	72	7	73	8
rect	72	10	73	11
rect	72	13	73	14
rect	72	16	73	17
rect	72	19	73	20
rect	72	22	73	23
rect	72	25	73	26
rect	72	28	73	29
rect	72	31	73	32
rect	72	34	73	35
rect	72	37	73	38
rect	72	40	73	41
rect	72	43	73	44
rect	72	46	73	47
rect	72	49	73	50
rect	72	52	73	53
rect	72	55	73	56
rect	72	58	73	59
rect	72	61	73	62
rect	72	64	73	65
rect	72	67	73	68
rect	72	70	73	71
rect	72	73	73	74
rect	72	76	73	77
rect	72	79	73	80
rect	72	82	73	83
rect	72	85	73	86
rect	72	88	73	89
rect	72	91	73	92
rect	72	97	73	98
rect	72	100	73	101
rect	72	103	73	104
rect	72	106	73	107
rect	72	109	73	110
rect	72	112	73	113
rect	72	115	73	116
rect	72	118	73	119
rect	72	121	73	122
rect	72	124	73	125
rect	72	127	73	128
rect	72	130	73	131
rect	72	133	73	134
rect	72	136	73	137
rect	72	139	73	140
rect	72	142	73	143
rect	72	145	73	146
rect	72	148	73	149
rect	72	151	73	152
rect	72	154	73	155
rect	72	157	73	158
rect	72	160	73	161
rect	72	163	73	164
rect	72	166	73	167
rect	72	169	73	170
rect	72	172	73	173
rect	72	175	73	176
rect	72	178	73	179
rect	72	181	73	182
rect	72	184	73	185
rect	72	187	73	188
rect	72	190	73	191
rect	72	193	73	194
rect	72	196	73	197
rect	72	199	73	200
rect	72	202	73	203
rect	72	205	73	206
rect	72	208	73	209
rect	72	211	73	212
rect	72	214	73	215
rect	72	217	73	218
rect	72	220	73	221
rect	72	223	73	224
rect	72	226	73	227
rect	72	229	73	230
rect	72	232	73	233
rect	72	235	73	236
rect	72	238	73	239
rect	72	241	73	242
rect	72	244	73	245
rect	72	247	73	248
rect	72	250	73	251
rect	72	253	73	254
rect	72	256	73	257
rect	72	259	73	260
rect	72	262	73	263
rect	72	265	73	266
rect	72	268	73	269
rect	72	271	73	272
rect	72	274	73	275
rect	72	277	73	278
rect	72	280	73	281
rect	72	283	73	284
rect	72	286	73	287
rect	72	289	73	290
rect	72	292	73	293
rect	72	295	73	296
rect	72	298	73	299
rect	72	301	73	302
rect	72	304	73	305
rect	72	310	73	311
rect	72	313	73	314
rect	72	316	73	317
rect	72	319	73	320
rect	72	322	73	323
rect	72	325	73	326
rect	72	328	73	329
rect	72	331	73	332
rect	72	334	73	335
rect	72	337	73	338
rect	72	340	73	341
rect	72	343	73	344
rect	72	346	73	347
rect	72	349	73	350
rect	72	352	73	353
rect	72	355	73	356
rect	72	358	73	359
rect	72	361	73	362
rect	72	364	73	365
rect	72	367	73	368
rect	72	373	73	374
rect	72	376	73	377
rect	72	379	73	380
rect	72	385	73	386
rect	73	1	74	2
rect	73	4	74	5
rect	73	7	74	8
rect	73	10	74	11
rect	73	13	74	14
rect	73	16	74	17
rect	73	19	74	20
rect	73	22	74	23
rect	73	25	74	26
rect	73	28	74	29
rect	73	31	74	32
rect	73	34	74	35
rect	73	37	74	38
rect	73	40	74	41
rect	73	43	74	44
rect	73	46	74	47
rect	73	49	74	50
rect	73	52	74	53
rect	73	55	74	56
rect	73	58	74	59
rect	73	61	74	62
rect	73	64	74	65
rect	73	67	74	68
rect	73	70	74	71
rect	73	73	74	74
rect	73	76	74	77
rect	73	79	74	80
rect	73	82	74	83
rect	73	85	74	86
rect	73	88	74	89
rect	73	91	74	92
rect	73	94	74	95
rect	73	97	74	98
rect	73	100	74	101
rect	73	103	74	104
rect	73	106	74	107
rect	73	109	74	110
rect	73	112	74	113
rect	73	115	74	116
rect	73	118	74	119
rect	73	121	74	122
rect	73	124	74	125
rect	73	127	74	128
rect	73	130	74	131
rect	73	133	74	134
rect	73	136	74	137
rect	73	139	74	140
rect	73	142	74	143
rect	73	145	74	146
rect	73	148	74	149
rect	73	151	74	152
rect	73	154	74	155
rect	73	157	74	158
rect	73	160	74	161
rect	73	163	74	164
rect	73	166	74	167
rect	73	169	74	170
rect	73	172	74	173
rect	73	175	74	176
rect	73	178	74	179
rect	73	181	74	182
rect	73	184	74	185
rect	73	187	74	188
rect	73	190	74	191
rect	73	193	74	194
rect	73	196	74	197
rect	73	199	74	200
rect	73	202	74	203
rect	73	205	74	206
rect	73	208	74	209
rect	73	211	74	212
rect	73	214	74	215
rect	73	217	74	218
rect	73	220	74	221
rect	73	223	74	224
rect	73	226	74	227
rect	73	229	74	230
rect	73	232	74	233
rect	73	235	74	236
rect	73	238	74	239
rect	73	241	74	242
rect	73	244	74	245
rect	73	247	74	248
rect	73	250	74	251
rect	73	253	74	254
rect	73	256	74	257
rect	73	259	74	260
rect	73	262	74	263
rect	73	265	74	266
rect	73	268	74	269
rect	73	271	74	272
rect	73	274	74	275
rect	73	277	74	278
rect	73	280	74	281
rect	73	283	74	284
rect	73	286	74	287
rect	73	289	74	290
rect	73	292	74	293
rect	73	295	74	296
rect	73	298	74	299
rect	73	301	74	302
rect	73	304	74	305
rect	73	307	74	308
rect	73	310	74	311
rect	73	313	74	314
rect	73	316	74	317
rect	73	319	74	320
rect	73	322	74	323
rect	73	325	74	326
rect	73	328	74	329
rect	73	331	74	332
rect	73	334	74	335
rect	73	337	74	338
rect	73	340	74	341
rect	73	343	74	344
rect	73	346	74	347
rect	73	349	74	350
rect	73	352	74	353
rect	73	355	74	356
rect	73	358	74	359
rect	73	361	74	362
rect	73	364	74	365
rect	73	367	74	368
rect	73	373	74	374
rect	73	376	74	377
rect	73	379	74	380
rect	73	385	74	386
rect	74	1	75	2
rect	74	4	75	5
rect	74	7	75	8
rect	74	10	75	11
rect	74	13	75	14
rect	74	16	75	17
rect	74	19	75	20
rect	74	22	75	23
rect	74	25	75	26
rect	74	28	75	29
rect	74	31	75	32
rect	74	34	75	35
rect	74	37	75	38
rect	74	40	75	41
rect	74	43	75	44
rect	74	46	75	47
rect	74	49	75	50
rect	74	52	75	53
rect	74	55	75	56
rect	74	58	75	59
rect	74	61	75	62
rect	74	64	75	65
rect	74	67	75	68
rect	74	70	75	71
rect	74	73	75	74
rect	74	76	75	77
rect	74	79	75	80
rect	74	82	75	83
rect	74	85	75	86
rect	74	88	75	89
rect	74	91	75	92
rect	74	94	75	95
rect	74	97	75	98
rect	74	100	75	101
rect	74	103	75	104
rect	74	106	75	107
rect	74	109	75	110
rect	74	112	75	113
rect	74	115	75	116
rect	74	118	75	119
rect	74	121	75	122
rect	74	124	75	125
rect	74	127	75	128
rect	74	130	75	131
rect	74	133	75	134
rect	74	136	75	137
rect	74	139	75	140
rect	74	142	75	143
rect	74	145	75	146
rect	74	148	75	149
rect	74	151	75	152
rect	74	154	75	155
rect	74	157	75	158
rect	74	160	75	161
rect	74	163	75	164
rect	74	166	75	167
rect	74	169	75	170
rect	74	172	75	173
rect	74	175	75	176
rect	74	178	75	179
rect	74	181	75	182
rect	74	184	75	185
rect	74	187	75	188
rect	74	190	75	191
rect	74	193	75	194
rect	74	196	75	197
rect	74	199	75	200
rect	74	202	75	203
rect	74	205	75	206
rect	74	208	75	209
rect	74	211	75	212
rect	74	214	75	215
rect	74	217	75	218
rect	74	220	75	221
rect	74	223	75	224
rect	74	226	75	227
rect	74	229	75	230
rect	74	232	75	233
rect	74	235	75	236
rect	74	238	75	239
rect	74	241	75	242
rect	74	244	75	245
rect	74	247	75	248
rect	74	250	75	251
rect	74	253	75	254
rect	74	256	75	257
rect	74	259	75	260
rect	74	262	75	263
rect	74	265	75	266
rect	74	268	75	269
rect	74	271	75	272
rect	74	274	75	275
rect	74	277	75	278
rect	74	280	75	281
rect	74	283	75	284
rect	74	286	75	287
rect	74	289	75	290
rect	74	292	75	293
rect	74	295	75	296
rect	74	298	75	299
rect	74	301	75	302
rect	74	304	75	305
rect	74	307	75	308
rect	74	310	75	311
rect	74	313	75	314
rect	74	316	75	317
rect	74	319	75	320
rect	74	322	75	323
rect	74	325	75	326
rect	74	328	75	329
rect	74	331	75	332
rect	74	334	75	335
rect	74	337	75	338
rect	74	340	75	341
rect	74	343	75	344
rect	74	346	75	347
rect	74	349	75	350
rect	74	352	75	353
rect	74	355	75	356
rect	74	358	75	359
rect	74	361	75	362
rect	74	364	75	365
rect	74	367	75	368
rect	74	373	75	374
rect	74	376	75	377
rect	74	379	75	380
rect	74	385	75	386
rect	75	1	76	2
rect	75	4	76	5
rect	75	7	76	8
rect	75	10	76	11
rect	75	13	76	14
rect	75	16	76	17
rect	75	19	76	20
rect	75	22	76	23
rect	75	25	76	26
rect	75	28	76	29
rect	75	31	76	32
rect	75	34	76	35
rect	75	37	76	38
rect	75	40	76	41
rect	75	43	76	44
rect	75	46	76	47
rect	75	49	76	50
rect	75	52	76	53
rect	75	55	76	56
rect	75	58	76	59
rect	75	61	76	62
rect	75	64	76	65
rect	75	67	76	68
rect	75	70	76	71
rect	75	73	76	74
rect	75	76	76	77
rect	75	79	76	80
rect	75	82	76	83
rect	75	85	76	86
rect	75	88	76	89
rect	75	91	76	92
rect	75	94	76	95
rect	75	97	76	98
rect	75	100	76	101
rect	75	103	76	104
rect	75	106	76	107
rect	75	109	76	110
rect	75	112	76	113
rect	75	115	76	116
rect	75	118	76	119
rect	75	121	76	122
rect	75	124	76	125
rect	75	127	76	128
rect	75	130	76	131
rect	75	133	76	134
rect	75	136	76	137
rect	75	139	76	140
rect	75	142	76	143
rect	75	145	76	146
rect	75	148	76	149
rect	75	151	76	152
rect	75	154	76	155
rect	75	157	76	158
rect	75	160	76	161
rect	75	163	76	164
rect	75	166	76	167
rect	75	169	76	170
rect	75	172	76	173
rect	75	175	76	176
rect	75	178	76	179
rect	75	181	76	182
rect	75	184	76	185
rect	75	187	76	188
rect	75	190	76	191
rect	75	193	76	194
rect	75	196	76	197
rect	75	199	76	200
rect	75	202	76	203
rect	75	205	76	206
rect	75	208	76	209
rect	75	211	76	212
rect	75	214	76	215
rect	75	217	76	218
rect	75	220	76	221
rect	75	223	76	224
rect	75	226	76	227
rect	75	229	76	230
rect	75	232	76	233
rect	75	235	76	236
rect	75	238	76	239
rect	75	241	76	242
rect	75	244	76	245
rect	75	247	76	248
rect	75	250	76	251
rect	75	253	76	254
rect	75	256	76	257
rect	75	259	76	260
rect	75	262	76	263
rect	75	265	76	266
rect	75	268	76	269
rect	75	271	76	272
rect	75	274	76	275
rect	75	277	76	278
rect	75	280	76	281
rect	75	283	76	284
rect	75	286	76	287
rect	75	289	76	290
rect	75	292	76	293
rect	75	295	76	296
rect	75	298	76	299
rect	75	301	76	302
rect	75	304	76	305
rect	75	307	76	308
rect	75	310	76	311
rect	75	313	76	314
rect	75	316	76	317
rect	75	319	76	320
rect	75	322	76	323
rect	75	325	76	326
rect	75	328	76	329
rect	75	331	76	332
rect	75	334	76	335
rect	75	337	76	338
rect	75	340	76	341
rect	75	343	76	344
rect	75	346	76	347
rect	75	349	76	350
rect	75	352	76	353
rect	75	355	76	356
rect	75	358	76	359
rect	75	361	76	362
rect	75	364	76	365
rect	75	367	76	368
rect	75	373	76	374
rect	75	376	76	377
rect	75	379	76	380
rect	75	385	76	386
rect	76	1	77	2
rect	76	4	77	5
rect	76	7	77	8
rect	76	10	77	11
rect	76	13	77	14
rect	76	16	77	17
rect	76	19	77	20
rect	76	22	77	23
rect	76	25	77	26
rect	76	28	77	29
rect	76	31	77	32
rect	76	34	77	35
rect	76	37	77	38
rect	76	40	77	41
rect	76	43	77	44
rect	76	46	77	47
rect	76	49	77	50
rect	76	52	77	53
rect	76	55	77	56
rect	76	58	77	59
rect	76	61	77	62
rect	76	64	77	65
rect	76	67	77	68
rect	76	70	77	71
rect	76	73	77	74
rect	76	76	77	77
rect	76	79	77	80
rect	76	82	77	83
rect	76	85	77	86
rect	76	88	77	89
rect	76	91	77	92
rect	76	94	77	95
rect	76	97	77	98
rect	76	100	77	101
rect	76	103	77	104
rect	76	106	77	107
rect	76	109	77	110
rect	76	112	77	113
rect	76	115	77	116
rect	76	118	77	119
rect	76	121	77	122
rect	76	124	77	125
rect	76	127	77	128
rect	76	130	77	131
rect	76	133	77	134
rect	76	136	77	137
rect	76	139	77	140
rect	76	142	77	143
rect	76	145	77	146
rect	76	148	77	149
rect	76	151	77	152
rect	76	154	77	155
rect	76	157	77	158
rect	76	160	77	161
rect	76	163	77	164
rect	76	166	77	167
rect	76	169	77	170
rect	76	172	77	173
rect	76	175	77	176
rect	76	178	77	179
rect	76	181	77	182
rect	76	184	77	185
rect	76	187	77	188
rect	76	190	77	191
rect	76	193	77	194
rect	76	196	77	197
rect	76	199	77	200
rect	76	202	77	203
rect	76	205	77	206
rect	76	208	77	209
rect	76	211	77	212
rect	76	214	77	215
rect	76	217	77	218
rect	76	220	77	221
rect	76	223	77	224
rect	76	226	77	227
rect	76	229	77	230
rect	76	232	77	233
rect	76	235	77	236
rect	76	238	77	239
rect	76	241	77	242
rect	76	244	77	245
rect	76	247	77	248
rect	76	250	77	251
rect	76	253	77	254
rect	76	256	77	257
rect	76	259	77	260
rect	76	262	77	263
rect	76	265	77	266
rect	76	268	77	269
rect	76	271	77	272
rect	76	274	77	275
rect	76	277	77	278
rect	76	280	77	281
rect	76	283	77	284
rect	76	286	77	287
rect	76	289	77	290
rect	76	292	77	293
rect	76	295	77	296
rect	76	298	77	299
rect	76	301	77	302
rect	76	304	77	305
rect	76	307	77	308
rect	76	310	77	311
rect	76	313	77	314
rect	76	316	77	317
rect	76	319	77	320
rect	76	322	77	323
rect	76	325	77	326
rect	76	328	77	329
rect	76	331	77	332
rect	76	334	77	335
rect	76	337	77	338
rect	76	340	77	341
rect	76	343	77	344
rect	76	346	77	347
rect	76	349	77	350
rect	76	352	77	353
rect	76	355	77	356
rect	76	358	77	359
rect	76	361	77	362
rect	76	364	77	365
rect	76	367	77	368
rect	76	373	77	374
rect	76	376	77	377
rect	76	379	77	380
rect	76	385	77	386
rect	77	1	78	2
rect	77	4	78	5
rect	77	7	78	8
rect	77	10	78	11
rect	77	13	78	14
rect	77	16	78	17
rect	77	19	78	20
rect	77	22	78	23
rect	77	25	78	26
rect	77	28	78	29
rect	77	31	78	32
rect	77	34	78	35
rect	77	37	78	38
rect	77	40	78	41
rect	77	43	78	44
rect	77	46	78	47
rect	77	49	78	50
rect	77	52	78	53
rect	77	55	78	56
rect	77	58	78	59
rect	77	61	78	62
rect	77	64	78	65
rect	77	67	78	68
rect	77	70	78	71
rect	77	73	78	74
rect	77	76	78	77
rect	77	79	78	80
rect	77	82	78	83
rect	77	85	78	86
rect	77	88	78	89
rect	77	91	78	92
rect	77	94	78	95
rect	77	97	78	98
rect	77	100	78	101
rect	77	103	78	104
rect	77	106	78	107
rect	77	109	78	110
rect	77	112	78	113
rect	77	115	78	116
rect	77	118	78	119
rect	77	121	78	122
rect	77	124	78	125
rect	77	127	78	128
rect	77	130	78	131
rect	77	133	78	134
rect	77	136	78	137
rect	77	139	78	140
rect	77	142	78	143
rect	77	145	78	146
rect	77	148	78	149
rect	77	151	78	152
rect	77	154	78	155
rect	77	157	78	158
rect	77	160	78	161
rect	77	163	78	164
rect	77	166	78	167
rect	77	169	78	170
rect	77	172	78	173
rect	77	175	78	176
rect	77	178	78	179
rect	77	181	78	182
rect	77	184	78	185
rect	77	187	78	188
rect	77	190	78	191
rect	77	193	78	194
rect	77	196	78	197
rect	77	199	78	200
rect	77	202	78	203
rect	77	205	78	206
rect	77	208	78	209
rect	77	211	78	212
rect	77	214	78	215
rect	77	217	78	218
rect	77	220	78	221
rect	77	223	78	224
rect	77	226	78	227
rect	77	229	78	230
rect	77	232	78	233
rect	77	235	78	236
rect	77	238	78	239
rect	77	241	78	242
rect	77	244	78	245
rect	77	247	78	248
rect	77	250	78	251
rect	77	253	78	254
rect	77	256	78	257
rect	77	259	78	260
rect	77	262	78	263
rect	77	265	78	266
rect	77	268	78	269
rect	77	271	78	272
rect	77	274	78	275
rect	77	277	78	278
rect	77	280	78	281
rect	77	283	78	284
rect	77	286	78	287
rect	77	289	78	290
rect	77	292	78	293
rect	77	295	78	296
rect	77	298	78	299
rect	77	301	78	302
rect	77	304	78	305
rect	77	307	78	308
rect	77	310	78	311
rect	77	313	78	314
rect	77	316	78	317
rect	77	319	78	320
rect	77	322	78	323
rect	77	325	78	326
rect	77	328	78	329
rect	77	331	78	332
rect	77	334	78	335
rect	77	337	78	338
rect	77	340	78	341
rect	77	343	78	344
rect	77	346	78	347
rect	77	349	78	350
rect	77	352	78	353
rect	77	355	78	356
rect	77	358	78	359
rect	77	361	78	362
rect	77	364	78	365
rect	77	367	78	368
rect	77	373	78	374
rect	77	376	78	377
rect	77	379	78	380
rect	77	385	78	386
rect	78	1	79	2
rect	78	4	79	5
rect	78	7	79	8
rect	78	10	79	11
rect	78	13	79	14
rect	78	16	79	17
rect	78	19	79	20
rect	78	22	79	23
rect	78	25	79	26
rect	78	28	79	29
rect	78	31	79	32
rect	78	34	79	35
rect	78	37	79	38
rect	78	40	79	41
rect	78	43	79	44
rect	78	46	79	47
rect	78	49	79	50
rect	78	52	79	53
rect	78	55	79	56
rect	78	58	79	59
rect	78	61	79	62
rect	78	64	79	65
rect	78	67	79	68
rect	78	70	79	71
rect	78	73	79	74
rect	78	76	79	77
rect	78	79	79	80
rect	78	82	79	83
rect	78	85	79	86
rect	78	88	79	89
rect	78	91	79	92
rect	78	94	79	95
rect	78	97	79	98
rect	78	100	79	101
rect	78	103	79	104
rect	78	106	79	107
rect	78	109	79	110
rect	78	112	79	113
rect	78	115	79	116
rect	78	118	79	119
rect	78	121	79	122
rect	78	124	79	125
rect	78	127	79	128
rect	78	130	79	131
rect	78	133	79	134
rect	78	136	79	137
rect	78	139	79	140
rect	78	142	79	143
rect	78	145	79	146
rect	78	148	79	149
rect	78	151	79	152
rect	78	154	79	155
rect	78	157	79	158
rect	78	160	79	161
rect	78	163	79	164
rect	78	166	79	167
rect	78	169	79	170
rect	78	172	79	173
rect	78	175	79	176
rect	78	178	79	179
rect	78	181	79	182
rect	78	184	79	185
rect	78	187	79	188
rect	78	190	79	191
rect	78	193	79	194
rect	78	196	79	197
rect	78	199	79	200
rect	78	202	79	203
rect	78	205	79	206
rect	78	208	79	209
rect	78	211	79	212
rect	78	214	79	215
rect	78	217	79	218
rect	78	220	79	221
rect	78	223	79	224
rect	78	226	79	227
rect	78	229	79	230
rect	78	232	79	233
rect	78	235	79	236
rect	78	238	79	239
rect	78	241	79	242
rect	78	244	79	245
rect	78	247	79	248
rect	78	250	79	251
rect	78	253	79	254
rect	78	256	79	257
rect	78	259	79	260
rect	78	262	79	263
rect	78	265	79	266
rect	78	268	79	269
rect	78	271	79	272
rect	78	274	79	275
rect	78	277	79	278
rect	78	280	79	281
rect	78	283	79	284
rect	78	286	79	287
rect	78	289	79	290
rect	78	292	79	293
rect	78	295	79	296
rect	78	298	79	299
rect	78	301	79	302
rect	78	304	79	305
rect	78	307	79	308
rect	78	310	79	311
rect	78	313	79	314
rect	78	316	79	317
rect	78	319	79	320
rect	78	322	79	323
rect	78	325	79	326
rect	78	328	79	329
rect	78	331	79	332
rect	78	334	79	335
rect	78	337	79	338
rect	78	340	79	341
rect	78	343	79	344
rect	78	346	79	347
rect	78	349	79	350
rect	78	352	79	353
rect	78	355	79	356
rect	78	358	79	359
rect	78	361	79	362
rect	78	364	79	365
rect	78	367	79	368
rect	78	373	79	374
rect	78	376	79	377
rect	78	379	79	380
rect	78	385	79	386
rect	79	1	80	2
rect	79	4	80	5
rect	79	7	80	8
rect	79	10	80	11
rect	79	13	80	14
rect	79	16	80	17
rect	79	19	80	20
rect	79	22	80	23
rect	79	25	80	26
rect	79	28	80	29
rect	79	31	80	32
rect	79	34	80	35
rect	79	37	80	38
rect	79	40	80	41
rect	79	43	80	44
rect	79	46	80	47
rect	79	49	80	50
rect	79	52	80	53
rect	79	55	80	56
rect	79	58	80	59
rect	79	61	80	62
rect	79	64	80	65
rect	79	67	80	68
rect	79	70	80	71
rect	79	73	80	74
rect	79	76	80	77
rect	79	79	80	80
rect	79	82	80	83
rect	79	85	80	86
rect	79	88	80	89
rect	79	91	80	92
rect	79	94	80	95
rect	79	97	80	98
rect	79	100	80	101
rect	79	103	80	104
rect	79	106	80	107
rect	79	109	80	110
rect	79	112	80	113
rect	79	115	80	116
rect	79	118	80	119
rect	79	121	80	122
rect	79	124	80	125
rect	79	127	80	128
rect	79	130	80	131
rect	79	133	80	134
rect	79	136	80	137
rect	79	139	80	140
rect	79	142	80	143
rect	79	145	80	146
rect	79	148	80	149
rect	79	151	80	152
rect	79	154	80	155
rect	79	157	80	158
rect	79	160	80	161
rect	79	163	80	164
rect	79	166	80	167
rect	79	169	80	170
rect	79	172	80	173
rect	79	175	80	176
rect	79	178	80	179
rect	79	181	80	182
rect	79	184	80	185
rect	79	187	80	188
rect	79	190	80	191
rect	79	193	80	194
rect	79	196	80	197
rect	79	199	80	200
rect	79	202	80	203
rect	79	205	80	206
rect	79	208	80	209
rect	79	211	80	212
rect	79	214	80	215
rect	79	217	80	218
rect	79	220	80	221
rect	79	223	80	224
rect	79	226	80	227
rect	79	229	80	230
rect	79	232	80	233
rect	79	235	80	236
rect	79	238	80	239
rect	79	241	80	242
rect	79	244	80	245
rect	79	247	80	248
rect	79	250	80	251
rect	79	253	80	254
rect	79	256	80	257
rect	79	259	80	260
rect	79	262	80	263
rect	79	265	80	266
rect	79	268	80	269
rect	79	271	80	272
rect	79	274	80	275
rect	79	277	80	278
rect	79	280	80	281
rect	79	283	80	284
rect	79	286	80	287
rect	79	289	80	290
rect	79	292	80	293
rect	79	295	80	296
rect	79	298	80	299
rect	79	301	80	302
rect	79	304	80	305
rect	79	307	80	308
rect	79	310	80	311
rect	79	313	80	314
rect	79	316	80	317
rect	79	319	80	320
rect	79	322	80	323
rect	79	325	80	326
rect	79	328	80	329
rect	79	331	80	332
rect	79	334	80	335
rect	79	337	80	338
rect	79	340	80	341
rect	79	343	80	344
rect	79	346	80	347
rect	79	349	80	350
rect	79	352	80	353
rect	79	355	80	356
rect	79	358	80	359
rect	79	361	80	362
rect	79	364	80	365
rect	79	367	80	368
rect	79	373	80	374
rect	79	376	80	377
rect	79	379	80	380
rect	79	385	80	386
rect	80	1	81	2
rect	80	4	81	5
rect	80	7	81	8
rect	80	10	81	11
rect	80	13	81	14
rect	80	16	81	17
rect	80	19	81	20
rect	80	22	81	23
rect	80	25	81	26
rect	80	28	81	29
rect	80	31	81	32
rect	80	34	81	35
rect	80	37	81	38
rect	80	40	81	41
rect	80	43	81	44
rect	80	46	81	47
rect	80	49	81	50
rect	80	52	81	53
rect	80	55	81	56
rect	80	58	81	59
rect	80	61	81	62
rect	80	64	81	65
rect	80	67	81	68
rect	80	70	81	71
rect	80	73	81	74
rect	80	76	81	77
rect	80	79	81	80
rect	80	82	81	83
rect	80	85	81	86
rect	80	88	81	89
rect	80	91	81	92
rect	80	94	81	95
rect	80	97	81	98
rect	80	100	81	101
rect	80	103	81	104
rect	80	106	81	107
rect	80	109	81	110
rect	80	112	81	113
rect	80	115	81	116
rect	80	118	81	119
rect	80	121	81	122
rect	80	124	81	125
rect	80	127	81	128
rect	80	130	81	131
rect	80	133	81	134
rect	80	136	81	137
rect	80	139	81	140
rect	80	142	81	143
rect	80	145	81	146
rect	80	148	81	149
rect	80	151	81	152
rect	80	154	81	155
rect	80	157	81	158
rect	80	160	81	161
rect	80	163	81	164
rect	80	166	81	167
rect	80	169	81	170
rect	80	172	81	173
rect	80	175	81	176
rect	80	178	81	179
rect	80	181	81	182
rect	80	184	81	185
rect	80	187	81	188
rect	80	190	81	191
rect	80	193	81	194
rect	80	196	81	197
rect	80	199	81	200
rect	80	202	81	203
rect	80	205	81	206
rect	80	208	81	209
rect	80	211	81	212
rect	80	214	81	215
rect	80	217	81	218
rect	80	220	81	221
rect	80	223	81	224
rect	80	226	81	227
rect	80	229	81	230
rect	80	232	81	233
rect	80	235	81	236
rect	80	238	81	239
rect	80	241	81	242
rect	80	244	81	245
rect	80	247	81	248
rect	80	250	81	251
rect	80	253	81	254
rect	80	256	81	257
rect	80	259	81	260
rect	80	262	81	263
rect	80	265	81	266
rect	80	268	81	269
rect	80	271	81	272
rect	80	274	81	275
rect	80	277	81	278
rect	80	280	81	281
rect	80	283	81	284
rect	80	286	81	287
rect	80	289	81	290
rect	80	292	81	293
rect	80	295	81	296
rect	80	298	81	299
rect	80	301	81	302
rect	80	304	81	305
rect	80	307	81	308
rect	80	310	81	311
rect	80	313	81	314
rect	80	316	81	317
rect	80	319	81	320
rect	80	322	81	323
rect	80	325	81	326
rect	80	328	81	329
rect	80	331	81	332
rect	80	334	81	335
rect	80	337	81	338
rect	80	340	81	341
rect	80	343	81	344
rect	80	346	81	347
rect	80	349	81	350
rect	80	352	81	353
rect	80	355	81	356
rect	80	358	81	359
rect	80	361	81	362
rect	80	364	81	365
rect	80	367	81	368
rect	80	373	81	374
rect	80	376	81	377
rect	80	379	81	380
rect	80	385	81	386
rect	81	1	82	2
rect	81	4	82	5
rect	81	7	82	8
rect	81	10	82	11
rect	81	13	82	14
rect	81	16	82	17
rect	81	19	82	20
rect	81	22	82	23
rect	81	25	82	26
rect	81	28	82	29
rect	81	31	82	32
rect	81	34	82	35
rect	81	37	82	38
rect	81	40	82	41
rect	81	43	82	44
rect	81	46	82	47
rect	81	49	82	50
rect	81	52	82	53
rect	81	55	82	56
rect	81	58	82	59
rect	81	61	82	62
rect	81	64	82	65
rect	81	67	82	68
rect	81	70	82	71
rect	81	73	82	74
rect	81	76	82	77
rect	81	79	82	80
rect	81	82	82	83
rect	81	85	82	86
rect	81	88	82	89
rect	81	91	82	92
rect	81	94	82	95
rect	81	97	82	98
rect	81	100	82	101
rect	81	103	82	104
rect	81	106	82	107
rect	81	109	82	110
rect	81	112	82	113
rect	81	115	82	116
rect	81	118	82	119
rect	81	121	82	122
rect	81	124	82	125
rect	81	127	82	128
rect	81	130	82	131
rect	81	133	82	134
rect	81	136	82	137
rect	81	139	82	140
rect	81	142	82	143
rect	81	145	82	146
rect	81	148	82	149
rect	81	151	82	152
rect	81	154	82	155
rect	81	157	82	158
rect	81	160	82	161
rect	81	163	82	164
rect	81	166	82	167
rect	81	169	82	170
rect	81	172	82	173
rect	81	175	82	176
rect	81	178	82	179
rect	81	181	82	182
rect	81	184	82	185
rect	81	187	82	188
rect	81	190	82	191
rect	81	193	82	194
rect	81	196	82	197
rect	81	199	82	200
rect	81	202	82	203
rect	81	205	82	206
rect	81	208	82	209
rect	81	211	82	212
rect	81	214	82	215
rect	81	217	82	218
rect	81	220	82	221
rect	81	223	82	224
rect	81	226	82	227
rect	81	229	82	230
rect	81	232	82	233
rect	81	235	82	236
rect	81	238	82	239
rect	81	241	82	242
rect	81	244	82	245
rect	81	247	82	248
rect	81	250	82	251
rect	81	253	82	254
rect	81	256	82	257
rect	81	259	82	260
rect	81	262	82	263
rect	81	265	82	266
rect	81	268	82	269
rect	81	271	82	272
rect	81	274	82	275
rect	81	277	82	278
rect	81	280	82	281
rect	81	283	82	284
rect	81	286	82	287
rect	81	289	82	290
rect	81	292	82	293
rect	81	295	82	296
rect	81	298	82	299
rect	81	301	82	302
rect	81	304	82	305
rect	81	307	82	308
rect	81	310	82	311
rect	81	313	82	314
rect	81	316	82	317
rect	81	319	82	320
rect	81	322	82	323
rect	81	325	82	326
rect	81	328	82	329
rect	81	331	82	332
rect	81	334	82	335
rect	81	337	82	338
rect	81	340	82	341
rect	81	343	82	344
rect	81	346	82	347
rect	81	349	82	350
rect	81	352	82	353
rect	81	355	82	356
rect	81	358	82	359
rect	81	361	82	362
rect	81	364	82	365
rect	81	367	82	368
rect	81	373	82	374
rect	81	376	82	377
rect	81	379	82	380
rect	81	385	82	386
rect	82	1	83	2
rect	82	4	83	5
rect	82	7	83	8
rect	82	10	83	11
rect	82	13	83	14
rect	82	16	83	17
rect	82	19	83	20
rect	82	22	83	23
rect	82	25	83	26
rect	82	28	83	29
rect	82	31	83	32
rect	82	34	83	35
rect	82	37	83	38
rect	82	40	83	41
rect	82	43	83	44
rect	82	46	83	47
rect	82	49	83	50
rect	82	52	83	53
rect	82	55	83	56
rect	82	58	83	59
rect	82	61	83	62
rect	82	64	83	65
rect	82	67	83	68
rect	82	70	83	71
rect	82	73	83	74
rect	82	76	83	77
rect	82	79	83	80
rect	82	82	83	83
rect	82	85	83	86
rect	82	88	83	89
rect	82	91	83	92
rect	82	94	83	95
rect	82	97	83	98
rect	82	100	83	101
rect	82	103	83	104
rect	82	106	83	107
rect	82	109	83	110
rect	82	112	83	113
rect	82	115	83	116
rect	82	118	83	119
rect	82	121	83	122
rect	82	124	83	125
rect	82	127	83	128
rect	82	130	83	131
rect	82	133	83	134
rect	82	136	83	137
rect	82	139	83	140
rect	82	142	83	143
rect	82	145	83	146
rect	82	148	83	149
rect	82	151	83	152
rect	82	154	83	155
rect	82	157	83	158
rect	82	160	83	161
rect	82	163	83	164
rect	82	166	83	167
rect	82	169	83	170
rect	82	172	83	173
rect	82	175	83	176
rect	82	178	83	179
rect	82	181	83	182
rect	82	184	83	185
rect	82	187	83	188
rect	82	190	83	191
rect	82	193	83	194
rect	82	196	83	197
rect	82	199	83	200
rect	82	202	83	203
rect	82	205	83	206
rect	82	208	83	209
rect	82	211	83	212
rect	82	214	83	215
rect	82	217	83	218
rect	82	220	83	221
rect	82	223	83	224
rect	82	226	83	227
rect	82	229	83	230
rect	82	232	83	233
rect	82	235	83	236
rect	82	238	83	239
rect	82	241	83	242
rect	82	244	83	245
rect	82	247	83	248
rect	82	250	83	251
rect	82	253	83	254
rect	82	256	83	257
rect	82	259	83	260
rect	82	262	83	263
rect	82	265	83	266
rect	82	268	83	269
rect	82	271	83	272
rect	82	274	83	275
rect	82	277	83	278
rect	82	280	83	281
rect	82	283	83	284
rect	82	286	83	287
rect	82	289	83	290
rect	82	292	83	293
rect	82	295	83	296
rect	82	298	83	299
rect	82	301	83	302
rect	82	304	83	305
rect	82	307	83	308
rect	82	310	83	311
rect	82	313	83	314
rect	82	316	83	317
rect	82	319	83	320
rect	82	322	83	323
rect	82	325	83	326
rect	82	328	83	329
rect	82	331	83	332
rect	82	334	83	335
rect	82	337	83	338
rect	82	340	83	341
rect	82	343	83	344
rect	82	346	83	347
rect	82	349	83	350
rect	82	352	83	353
rect	82	355	83	356
rect	82	358	83	359
rect	82	361	83	362
rect	82	364	83	365
rect	82	367	83	368
rect	82	373	83	374
rect	82	376	83	377
rect	82	379	83	380
rect	82	385	83	386
rect	83	1	84	2
rect	83	4	84	5
rect	83	7	84	8
rect	83	10	84	11
rect	83	13	84	14
rect	83	16	84	17
rect	83	19	84	20
rect	83	22	84	23
rect	83	25	84	26
rect	83	28	84	29
rect	83	31	84	32
rect	83	34	84	35
rect	83	37	84	38
rect	83	40	84	41
rect	83	43	84	44
rect	83	46	84	47
rect	83	49	84	50
rect	83	52	84	53
rect	83	55	84	56
rect	83	58	84	59
rect	83	61	84	62
rect	83	64	84	65
rect	83	67	84	68
rect	83	70	84	71
rect	83	73	84	74
rect	83	76	84	77
rect	83	79	84	80
rect	83	82	84	83
rect	83	85	84	86
rect	83	88	84	89
rect	83	91	84	92
rect	83	94	84	95
rect	83	97	84	98
rect	83	100	84	101
rect	83	103	84	104
rect	83	106	84	107
rect	83	109	84	110
rect	83	112	84	113
rect	83	115	84	116
rect	83	118	84	119
rect	83	121	84	122
rect	83	124	84	125
rect	83	127	84	128
rect	83	130	84	131
rect	83	133	84	134
rect	83	136	84	137
rect	83	139	84	140
rect	83	142	84	143
rect	83	145	84	146
rect	83	148	84	149
rect	83	151	84	152
rect	83	154	84	155
rect	83	157	84	158
rect	83	160	84	161
rect	83	163	84	164
rect	83	166	84	167
rect	83	169	84	170
rect	83	172	84	173
rect	83	175	84	176
rect	83	178	84	179
rect	83	181	84	182
rect	83	184	84	185
rect	83	187	84	188
rect	83	190	84	191
rect	83	193	84	194
rect	83	196	84	197
rect	83	199	84	200
rect	83	202	84	203
rect	83	205	84	206
rect	83	208	84	209
rect	83	211	84	212
rect	83	214	84	215
rect	83	217	84	218
rect	83	220	84	221
rect	83	223	84	224
rect	83	226	84	227
rect	83	229	84	230
rect	83	232	84	233
rect	83	235	84	236
rect	83	238	84	239
rect	83	241	84	242
rect	83	244	84	245
rect	83	247	84	248
rect	83	250	84	251
rect	83	253	84	254
rect	83	256	84	257
rect	83	259	84	260
rect	83	262	84	263
rect	83	265	84	266
rect	83	268	84	269
rect	83	271	84	272
rect	83	274	84	275
rect	83	277	84	278
rect	83	280	84	281
rect	83	283	84	284
rect	83	286	84	287
rect	83	289	84	290
rect	83	292	84	293
rect	83	295	84	296
rect	83	298	84	299
rect	83	301	84	302
rect	83	304	84	305
rect	83	307	84	308
rect	83	310	84	311
rect	83	313	84	314
rect	83	316	84	317
rect	83	319	84	320
rect	83	322	84	323
rect	83	325	84	326
rect	83	328	84	329
rect	83	331	84	332
rect	83	334	84	335
rect	83	337	84	338
rect	83	340	84	341
rect	83	343	84	344
rect	83	346	84	347
rect	83	349	84	350
rect	83	352	84	353
rect	83	355	84	356
rect	83	358	84	359
rect	83	361	84	362
rect	83	364	84	365
rect	83	367	84	368
rect	83	373	84	374
rect	83	376	84	377
rect	83	379	84	380
rect	83	385	84	386
rect	84	1	85	2
rect	84	4	85	5
rect	84	7	85	8
rect	84	10	85	11
rect	84	13	85	14
rect	84	16	85	17
rect	84	19	85	20
rect	84	22	85	23
rect	84	25	85	26
rect	84	28	85	29
rect	84	31	85	32
rect	84	34	85	35
rect	84	37	85	38
rect	84	40	85	41
rect	84	43	85	44
rect	84	46	85	47
rect	84	49	85	50
rect	84	52	85	53
rect	84	55	85	56
rect	84	58	85	59
rect	84	61	85	62
rect	84	64	85	65
rect	84	67	85	68
rect	84	70	85	71
rect	84	73	85	74
rect	84	76	85	77
rect	84	79	85	80
rect	84	82	85	83
rect	84	85	85	86
rect	84	88	85	89
rect	84	91	85	92
rect	84	94	85	95
rect	84	97	85	98
rect	84	100	85	101
rect	84	103	85	104
rect	84	106	85	107
rect	84	109	85	110
rect	84	112	85	113
rect	84	115	85	116
rect	84	118	85	119
rect	84	121	85	122
rect	84	124	85	125
rect	84	127	85	128
rect	84	130	85	131
rect	84	133	85	134
rect	84	136	85	137
rect	84	139	85	140
rect	84	142	85	143
rect	84	145	85	146
rect	84	148	85	149
rect	84	151	85	152
rect	84	154	85	155
rect	84	157	85	158
rect	84	160	85	161
rect	84	163	85	164
rect	84	166	85	167
rect	84	169	85	170
rect	84	172	85	173
rect	84	175	85	176
rect	84	178	85	179
rect	84	181	85	182
rect	84	184	85	185
rect	84	187	85	188
rect	84	190	85	191
rect	84	193	85	194
rect	84	196	85	197
rect	84	199	85	200
rect	84	202	85	203
rect	84	205	85	206
rect	84	208	85	209
rect	84	211	85	212
rect	84	214	85	215
rect	84	217	85	218
rect	84	220	85	221
rect	84	223	85	224
rect	84	226	85	227
rect	84	229	85	230
rect	84	232	85	233
rect	84	235	85	236
rect	84	238	85	239
rect	84	241	85	242
rect	84	244	85	245
rect	84	247	85	248
rect	84	250	85	251
rect	84	253	85	254
rect	84	256	85	257
rect	84	259	85	260
rect	84	262	85	263
rect	84	265	85	266
rect	84	268	85	269
rect	84	271	85	272
rect	84	274	85	275
rect	84	277	85	278
rect	84	280	85	281
rect	84	283	85	284
rect	84	286	85	287
rect	84	289	85	290
rect	84	292	85	293
rect	84	295	85	296
rect	84	298	85	299
rect	84	301	85	302
rect	84	304	85	305
rect	84	307	85	308
rect	84	310	85	311
rect	84	313	85	314
rect	84	316	85	317
rect	84	319	85	320
rect	84	322	85	323
rect	84	325	85	326
rect	84	328	85	329
rect	84	331	85	332
rect	84	334	85	335
rect	84	337	85	338
rect	84	340	85	341
rect	84	343	85	344
rect	84	346	85	347
rect	84	349	85	350
rect	84	352	85	353
rect	84	355	85	356
rect	84	358	85	359
rect	84	361	85	362
rect	84	364	85	365
rect	84	367	85	368
rect	84	373	85	374
rect	84	376	85	377
rect	84	379	85	380
rect	84	385	85	386
rect	85	1	86	2
rect	85	4	86	5
rect	85	7	86	8
rect	85	10	86	11
rect	85	13	86	14
rect	85	16	86	17
rect	85	19	86	20
rect	85	22	86	23
rect	85	25	86	26
rect	85	28	86	29
rect	85	31	86	32
rect	85	34	86	35
rect	85	37	86	38
rect	85	40	86	41
rect	85	43	86	44
rect	85	46	86	47
rect	85	49	86	50
rect	85	52	86	53
rect	85	55	86	56
rect	85	58	86	59
rect	85	61	86	62
rect	85	64	86	65
rect	85	67	86	68
rect	85	70	86	71
rect	85	73	86	74
rect	85	76	86	77
rect	85	79	86	80
rect	85	82	86	83
rect	85	85	86	86
rect	85	88	86	89
rect	85	91	86	92
rect	85	94	86	95
rect	85	97	86	98
rect	85	100	86	101
rect	85	103	86	104
rect	85	106	86	107
rect	85	109	86	110
rect	85	112	86	113
rect	85	115	86	116
rect	85	118	86	119
rect	85	121	86	122
rect	85	124	86	125
rect	85	127	86	128
rect	85	130	86	131
rect	85	133	86	134
rect	85	136	86	137
rect	85	139	86	140
rect	85	142	86	143
rect	85	145	86	146
rect	85	148	86	149
rect	85	151	86	152
rect	85	154	86	155
rect	85	157	86	158
rect	85	160	86	161
rect	85	163	86	164
rect	85	166	86	167
rect	85	169	86	170
rect	85	172	86	173
rect	85	175	86	176
rect	85	178	86	179
rect	85	181	86	182
rect	85	184	86	185
rect	85	187	86	188
rect	85	190	86	191
rect	85	193	86	194
rect	85	196	86	197
rect	85	199	86	200
rect	85	202	86	203
rect	85	205	86	206
rect	85	208	86	209
rect	85	211	86	212
rect	85	214	86	215
rect	85	217	86	218
rect	85	220	86	221
rect	85	223	86	224
rect	85	226	86	227
rect	85	229	86	230
rect	85	232	86	233
rect	85	235	86	236
rect	85	238	86	239
rect	85	241	86	242
rect	85	244	86	245
rect	85	247	86	248
rect	85	250	86	251
rect	85	253	86	254
rect	85	256	86	257
rect	85	259	86	260
rect	85	262	86	263
rect	85	265	86	266
rect	85	268	86	269
rect	85	271	86	272
rect	85	274	86	275
rect	85	277	86	278
rect	85	280	86	281
rect	85	283	86	284
rect	85	286	86	287
rect	85	289	86	290
rect	85	292	86	293
rect	85	295	86	296
rect	85	298	86	299
rect	85	301	86	302
rect	85	304	86	305
rect	85	307	86	308
rect	85	310	86	311
rect	85	313	86	314
rect	85	316	86	317
rect	85	319	86	320
rect	85	322	86	323
rect	85	325	86	326
rect	85	328	86	329
rect	85	331	86	332
rect	85	334	86	335
rect	85	337	86	338
rect	85	340	86	341
rect	85	343	86	344
rect	85	346	86	347
rect	85	349	86	350
rect	85	352	86	353
rect	85	355	86	356
rect	85	358	86	359
rect	85	361	86	362
rect	85	364	86	365
rect	85	367	86	368
rect	85	373	86	374
rect	85	376	86	377
rect	85	379	86	380
rect	85	385	86	386
rect	86	1	87	2
rect	86	4	87	5
rect	86	7	87	8
rect	86	10	87	11
rect	86	13	87	14
rect	86	16	87	17
rect	86	19	87	20
rect	86	22	87	23
rect	86	25	87	26
rect	86	28	87	29
rect	86	31	87	32
rect	86	34	87	35
rect	86	37	87	38
rect	86	40	87	41
rect	86	43	87	44
rect	86	46	87	47
rect	86	49	87	50
rect	86	52	87	53
rect	86	55	87	56
rect	86	58	87	59
rect	86	61	87	62
rect	86	64	87	65
rect	86	67	87	68
rect	86	70	87	71
rect	86	73	87	74
rect	86	76	87	77
rect	86	79	87	80
rect	86	82	87	83
rect	86	85	87	86
rect	86	88	87	89
rect	86	91	87	92
rect	86	94	87	95
rect	86	97	87	98
rect	86	100	87	101
rect	86	103	87	104
rect	86	106	87	107
rect	86	109	87	110
rect	86	112	87	113
rect	86	115	87	116
rect	86	118	87	119
rect	86	121	87	122
rect	86	124	87	125
rect	86	127	87	128
rect	86	130	87	131
rect	86	133	87	134
rect	86	136	87	137
rect	86	139	87	140
rect	86	142	87	143
rect	86	145	87	146
rect	86	148	87	149
rect	86	151	87	152
rect	86	154	87	155
rect	86	157	87	158
rect	86	160	87	161
rect	86	163	87	164
rect	86	166	87	167
rect	86	169	87	170
rect	86	172	87	173
rect	86	175	87	176
rect	86	178	87	179
rect	86	181	87	182
rect	86	184	87	185
rect	86	187	87	188
rect	86	190	87	191
rect	86	193	87	194
rect	86	196	87	197
rect	86	199	87	200
rect	86	202	87	203
rect	86	205	87	206
rect	86	208	87	209
rect	86	211	87	212
rect	86	214	87	215
rect	86	217	87	218
rect	86	220	87	221
rect	86	223	87	224
rect	86	226	87	227
rect	86	229	87	230
rect	86	232	87	233
rect	86	235	87	236
rect	86	238	87	239
rect	86	241	87	242
rect	86	244	87	245
rect	86	247	87	248
rect	86	250	87	251
rect	86	253	87	254
rect	86	256	87	257
rect	86	259	87	260
rect	86	262	87	263
rect	86	265	87	266
rect	86	268	87	269
rect	86	271	87	272
rect	86	274	87	275
rect	86	277	87	278
rect	86	280	87	281
rect	86	283	87	284
rect	86	286	87	287
rect	86	289	87	290
rect	86	292	87	293
rect	86	295	87	296
rect	86	298	87	299
rect	86	301	87	302
rect	86	304	87	305
rect	86	307	87	308
rect	86	310	87	311
rect	86	313	87	314
rect	86	316	87	317
rect	86	319	87	320
rect	86	322	87	323
rect	86	325	87	326
rect	86	328	87	329
rect	86	331	87	332
rect	86	334	87	335
rect	86	337	87	338
rect	86	340	87	341
rect	86	343	87	344
rect	86	346	87	347
rect	86	349	87	350
rect	86	352	87	353
rect	86	355	87	356
rect	86	358	87	359
rect	86	361	87	362
rect	86	364	87	365
rect	86	367	87	368
rect	86	373	87	374
rect	86	376	87	377
rect	86	379	87	380
rect	86	385	87	386
rect	87	1	88	2
rect	87	4	88	5
rect	87	7	88	8
rect	87	10	88	11
rect	87	13	88	14
rect	87	16	88	17
rect	87	19	88	20
rect	87	22	88	23
rect	87	25	88	26
rect	87	28	88	29
rect	87	31	88	32
rect	87	34	88	35
rect	87	37	88	38
rect	87	40	88	41
rect	87	43	88	44
rect	87	46	88	47
rect	87	49	88	50
rect	87	52	88	53
rect	87	55	88	56
rect	87	58	88	59
rect	87	61	88	62
rect	87	64	88	65
rect	87	67	88	68
rect	87	70	88	71
rect	87	73	88	74
rect	87	76	88	77
rect	87	79	88	80
rect	87	82	88	83
rect	87	85	88	86
rect	87	88	88	89
rect	87	91	88	92
rect	87	94	88	95
rect	87	97	88	98
rect	87	100	88	101
rect	87	103	88	104
rect	87	106	88	107
rect	87	109	88	110
rect	87	115	88	116
rect	87	118	88	119
rect	87	121	88	122
rect	87	124	88	125
rect	87	127	88	128
rect	87	130	88	131
rect	87	133	88	134
rect	87	136	88	137
rect	87	139	88	140
rect	87	142	88	143
rect	87	145	88	146
rect	87	148	88	149
rect	87	151	88	152
rect	87	154	88	155
rect	87	157	88	158
rect	87	160	88	161
rect	87	163	88	164
rect	87	166	88	167
rect	87	169	88	170
rect	87	172	88	173
rect	87	175	88	176
rect	87	178	88	179
rect	87	181	88	182
rect	87	184	88	185
rect	87	187	88	188
rect	87	190	88	191
rect	87	193	88	194
rect	87	196	88	197
rect	87	199	88	200
rect	87	202	88	203
rect	87	205	88	206
rect	87	208	88	209
rect	87	211	88	212
rect	87	214	88	215
rect	87	217	88	218
rect	87	220	88	221
rect	87	223	88	224
rect	87	226	88	227
rect	87	229	88	230
rect	87	232	88	233
rect	87	235	88	236
rect	87	238	88	239
rect	87	241	88	242
rect	87	244	88	245
rect	87	247	88	248
rect	87	250	88	251
rect	87	253	88	254
rect	87	256	88	257
rect	87	259	88	260
rect	87	262	88	263
rect	87	265	88	266
rect	87	268	88	269
rect	87	271	88	272
rect	87	274	88	275
rect	87	277	88	278
rect	87	280	88	281
rect	87	283	88	284
rect	87	286	88	287
rect	87	289	88	290
rect	87	292	88	293
rect	87	295	88	296
rect	87	298	88	299
rect	87	301	88	302
rect	87	304	88	305
rect	87	307	88	308
rect	87	310	88	311
rect	87	313	88	314
rect	87	316	88	317
rect	87	319	88	320
rect	87	322	88	323
rect	87	325	88	326
rect	87	328	88	329
rect	87	331	88	332
rect	87	334	88	335
rect	87	337	88	338
rect	87	340	88	341
rect	87	343	88	344
rect	87	346	88	347
rect	87	349	88	350
rect	87	352	88	353
rect	87	355	88	356
rect	87	358	88	359
rect	87	361	88	362
rect	87	364	88	365
rect	87	367	88	368
rect	87	373	88	374
rect	87	376	88	377
rect	87	379	88	380
rect	87	385	88	386
rect	88	1	89	2
rect	88	4	89	5
rect	88	7	89	8
rect	88	10	89	11
rect	88	13	89	14
rect	88	16	89	17
rect	88	19	89	20
rect	88	22	89	23
rect	88	25	89	26
rect	88	28	89	29
rect	88	31	89	32
rect	88	34	89	35
rect	88	37	89	38
rect	88	40	89	41
rect	88	43	89	44
rect	88	46	89	47
rect	88	49	89	50
rect	88	52	89	53
rect	88	55	89	56
rect	88	58	89	59
rect	88	61	89	62
rect	88	64	89	65
rect	88	67	89	68
rect	88	70	89	71
rect	88	73	89	74
rect	88	76	89	77
rect	88	79	89	80
rect	88	82	89	83
rect	88	85	89	86
rect	88	88	89	89
rect	88	91	89	92
rect	88	94	89	95
rect	88	97	89	98
rect	88	100	89	101
rect	88	103	89	104
rect	88	106	89	107
rect	88	109	89	110
rect	88	112	89	113
rect	88	115	89	116
rect	88	118	89	119
rect	88	121	89	122
rect	88	124	89	125
rect	88	127	89	128
rect	88	130	89	131
rect	88	133	89	134
rect	88	136	89	137
rect	88	139	89	140
rect	88	142	89	143
rect	88	145	89	146
rect	88	148	89	149
rect	88	151	89	152
rect	88	154	89	155
rect	88	157	89	158
rect	88	160	89	161
rect	88	163	89	164
rect	88	166	89	167
rect	88	169	89	170
rect	88	172	89	173
rect	88	175	89	176
rect	88	178	89	179
rect	88	181	89	182
rect	88	184	89	185
rect	88	187	89	188
rect	88	190	89	191
rect	88	193	89	194
rect	88	196	89	197
rect	88	199	89	200
rect	88	202	89	203
rect	88	205	89	206
rect	88	208	89	209
rect	88	211	89	212
rect	88	214	89	215
rect	88	217	89	218
rect	88	220	89	221
rect	88	223	89	224
rect	88	226	89	227
rect	88	229	89	230
rect	88	232	89	233
rect	88	235	89	236
rect	88	238	89	239
rect	88	241	89	242
rect	88	244	89	245
rect	88	247	89	248
rect	88	250	89	251
rect	88	253	89	254
rect	88	256	89	257
rect	88	259	89	260
rect	88	262	89	263
rect	88	265	89	266
rect	88	268	89	269
rect	88	271	89	272
rect	88	274	89	275
rect	88	277	89	278
rect	88	280	89	281
rect	88	283	89	284
rect	88	286	89	287
rect	88	289	89	290
rect	88	292	89	293
rect	88	295	89	296
rect	88	298	89	299
rect	88	301	89	302
rect	88	304	89	305
rect	88	307	89	308
rect	88	310	89	311
rect	88	313	89	314
rect	88	316	89	317
rect	88	319	89	320
rect	88	322	89	323
rect	88	325	89	326
rect	88	328	89	329
rect	88	331	89	332
rect	88	334	89	335
rect	88	337	89	338
rect	88	340	89	341
rect	88	343	89	344
rect	88	346	89	347
rect	88	349	89	350
rect	88	352	89	353
rect	88	355	89	356
rect	88	358	89	359
rect	88	361	89	362
rect	88	364	89	365
rect	88	367	89	368
rect	88	373	89	374
rect	88	376	89	377
rect	88	379	89	380
rect	88	385	89	386
rect	89	1	90	2
rect	89	4	90	5
rect	89	7	90	8
rect	89	10	90	11
rect	89	13	90	14
rect	89	16	90	17
rect	89	19	90	20
rect	89	22	90	23
rect	89	25	90	26
rect	89	28	90	29
rect	89	31	90	32
rect	89	37	90	38
rect	89	40	90	41
rect	89	43	90	44
rect	89	46	90	47
rect	89	49	90	50
rect	89	52	90	53
rect	89	55	90	56
rect	89	58	90	59
rect	89	61	90	62
rect	89	64	90	65
rect	89	67	90	68
rect	89	70	90	71
rect	89	73	90	74
rect	89	76	90	77
rect	89	79	90	80
rect	89	82	90	83
rect	89	85	90	86
rect	89	88	90	89
rect	89	91	90	92
rect	89	94	90	95
rect	89	97	90	98
rect	89	100	90	101
rect	89	103	90	104
rect	89	106	90	107
rect	89	109	90	110
rect	89	112	90	113
rect	89	115	90	116
rect	89	118	90	119
rect	89	121	90	122
rect	89	124	90	125
rect	89	127	90	128
rect	89	130	90	131
rect	89	133	90	134
rect	89	136	90	137
rect	89	139	90	140
rect	89	142	90	143
rect	89	145	90	146
rect	89	148	90	149
rect	89	151	90	152
rect	89	154	90	155
rect	89	157	90	158
rect	89	160	90	161
rect	89	166	90	167
rect	89	169	90	170
rect	89	172	90	173
rect	89	175	90	176
rect	89	178	90	179
rect	89	181	90	182
rect	89	184	90	185
rect	89	187	90	188
rect	89	190	90	191
rect	89	193	90	194
rect	89	196	90	197
rect	89	199	90	200
rect	89	202	90	203
rect	89	205	90	206
rect	89	208	90	209
rect	89	211	90	212
rect	89	214	90	215
rect	89	217	90	218
rect	89	220	90	221
rect	89	223	90	224
rect	89	226	90	227
rect	89	229	90	230
rect	89	232	90	233
rect	89	235	90	236
rect	89	238	90	239
rect	89	241	90	242
rect	89	244	90	245
rect	89	247	90	248
rect	89	250	90	251
rect	89	253	90	254
rect	89	256	90	257
rect	89	259	90	260
rect	89	262	90	263
rect	89	265	90	266
rect	89	268	90	269
rect	89	271	90	272
rect	89	274	90	275
rect	89	277	90	278
rect	89	280	90	281
rect	89	283	90	284
rect	89	286	90	287
rect	89	289	90	290
rect	89	292	90	293
rect	89	295	90	296
rect	89	298	90	299
rect	89	301	90	302
rect	89	304	90	305
rect	89	307	90	308
rect	89	310	90	311
rect	89	313	90	314
rect	89	316	90	317
rect	89	319	90	320
rect	89	322	90	323
rect	89	325	90	326
rect	89	328	90	329
rect	89	331	90	332
rect	89	334	90	335
rect	89	337	90	338
rect	89	340	90	341
rect	89	343	90	344
rect	89	346	90	347
rect	89	349	90	350
rect	89	352	90	353
rect	89	355	90	356
rect	89	358	90	359
rect	89	361	90	362
rect	89	364	90	365
rect	89	367	90	368
rect	89	373	90	374
rect	89	376	90	377
rect	89	379	90	380
rect	89	385	90	386
rect	90	1	91	2
rect	90	4	91	5
rect	90	7	91	8
rect	90	10	91	11
rect	90	13	91	14
rect	90	16	91	17
rect	90	19	91	20
rect	90	22	91	23
rect	90	25	91	26
rect	90	28	91	29
rect	90	31	91	32
rect	90	34	91	35
rect	90	37	91	38
rect	90	40	91	41
rect	90	43	91	44
rect	90	46	91	47
rect	90	49	91	50
rect	90	52	91	53
rect	90	55	91	56
rect	90	58	91	59
rect	90	61	91	62
rect	90	64	91	65
rect	90	67	91	68
rect	90	70	91	71
rect	90	73	91	74
rect	90	76	91	77
rect	90	79	91	80
rect	90	82	91	83
rect	90	85	91	86
rect	90	88	91	89
rect	90	91	91	92
rect	90	94	91	95
rect	90	97	91	98
rect	90	100	91	101
rect	90	103	91	104
rect	90	106	91	107
rect	90	109	91	110
rect	90	112	91	113
rect	90	115	91	116
rect	90	118	91	119
rect	90	121	91	122
rect	90	124	91	125
rect	90	127	91	128
rect	90	130	91	131
rect	90	133	91	134
rect	90	136	91	137
rect	90	139	91	140
rect	90	142	91	143
rect	90	145	91	146
rect	90	148	91	149
rect	90	151	91	152
rect	90	154	91	155
rect	90	157	91	158
rect	90	160	91	161
rect	90	163	91	164
rect	90	166	91	167
rect	90	169	91	170
rect	90	172	91	173
rect	90	175	91	176
rect	90	178	91	179
rect	90	181	91	182
rect	90	184	91	185
rect	90	187	91	188
rect	90	190	91	191
rect	90	193	91	194
rect	90	196	91	197
rect	90	199	91	200
rect	90	202	91	203
rect	90	205	91	206
rect	90	208	91	209
rect	90	211	91	212
rect	90	214	91	215
rect	90	217	91	218
rect	90	220	91	221
rect	90	223	91	224
rect	90	226	91	227
rect	90	229	91	230
rect	90	232	91	233
rect	90	235	91	236
rect	90	238	91	239
rect	90	241	91	242
rect	90	244	91	245
rect	90	247	91	248
rect	90	250	91	251
rect	90	253	91	254
rect	90	256	91	257
rect	90	259	91	260
rect	90	262	91	263
rect	90	265	91	266
rect	90	268	91	269
rect	90	271	91	272
rect	90	274	91	275
rect	90	277	91	278
rect	90	280	91	281
rect	90	283	91	284
rect	90	286	91	287
rect	90	289	91	290
rect	90	292	91	293
rect	90	295	91	296
rect	90	298	91	299
rect	90	301	91	302
rect	90	304	91	305
rect	90	307	91	308
rect	90	310	91	311
rect	90	313	91	314
rect	90	316	91	317
rect	90	319	91	320
rect	90	322	91	323
rect	90	325	91	326
rect	90	328	91	329
rect	90	331	91	332
rect	90	334	91	335
rect	90	337	91	338
rect	90	340	91	341
rect	90	343	91	344
rect	90	346	91	347
rect	90	349	91	350
rect	90	352	91	353
rect	90	355	91	356
rect	90	358	91	359
rect	90	361	91	362
rect	90	364	91	365
rect	90	367	91	368
rect	90	373	91	374
rect	90	376	91	377
rect	90	379	91	380
rect	90	385	91	386
rect	91	1	92	2
rect	91	4	92	5
rect	91	7	92	8
rect	91	10	92	11
rect	91	13	92	14
rect	91	16	92	17
rect	91	19	92	20
rect	91	22	92	23
rect	91	25	92	26
rect	91	28	92	29
rect	91	31	92	32
rect	91	34	92	35
rect	91	37	92	38
rect	91	40	92	41
rect	91	43	92	44
rect	91	46	92	47
rect	91	49	92	50
rect	91	52	92	53
rect	91	55	92	56
rect	91	58	92	59
rect	91	61	92	62
rect	91	64	92	65
rect	91	67	92	68
rect	91	70	92	71
rect	91	73	92	74
rect	91	76	92	77
rect	91	79	92	80
rect	91	82	92	83
rect	91	85	92	86
rect	91	88	92	89
rect	91	91	92	92
rect	91	94	92	95
rect	91	97	92	98
rect	91	100	92	101
rect	91	103	92	104
rect	91	106	92	107
rect	91	109	92	110
rect	91	112	92	113
rect	91	115	92	116
rect	91	118	92	119
rect	91	121	92	122
rect	91	124	92	125
rect	91	127	92	128
rect	91	130	92	131
rect	91	133	92	134
rect	91	136	92	137
rect	91	139	92	140
rect	91	142	92	143
rect	91	145	92	146
rect	91	148	92	149
rect	91	151	92	152
rect	91	154	92	155
rect	91	157	92	158
rect	91	160	92	161
rect	91	163	92	164
rect	91	166	92	167
rect	91	169	92	170
rect	91	172	92	173
rect	91	175	92	176
rect	91	178	92	179
rect	91	181	92	182
rect	91	184	92	185
rect	91	187	92	188
rect	91	190	92	191
rect	91	193	92	194
rect	91	196	92	197
rect	91	199	92	200
rect	91	202	92	203
rect	91	205	92	206
rect	91	208	92	209
rect	91	211	92	212
rect	91	214	92	215
rect	91	217	92	218
rect	91	220	92	221
rect	91	223	92	224
rect	91	226	92	227
rect	91	229	92	230
rect	91	232	92	233
rect	91	235	92	236
rect	91	238	92	239
rect	91	241	92	242
rect	91	244	92	245
rect	91	247	92	248
rect	91	250	92	251
rect	91	253	92	254
rect	91	256	92	257
rect	91	259	92	260
rect	91	262	92	263
rect	91	265	92	266
rect	91	268	92	269
rect	91	271	92	272
rect	91	274	92	275
rect	91	277	92	278
rect	91	280	92	281
rect	91	283	92	284
rect	91	286	92	287
rect	91	289	92	290
rect	91	292	92	293
rect	91	295	92	296
rect	91	298	92	299
rect	91	301	92	302
rect	91	304	92	305
rect	91	310	92	311
rect	91	316	92	317
rect	91	319	92	320
rect	91	322	92	323
rect	91	325	92	326
rect	91	328	92	329
rect	91	331	92	332
rect	91	334	92	335
rect	91	337	92	338
rect	91	340	92	341
rect	91	343	92	344
rect	91	346	92	347
rect	91	349	92	350
rect	91	352	92	353
rect	91	355	92	356
rect	91	358	92	359
rect	91	361	92	362
rect	91	364	92	365
rect	91	367	92	368
rect	91	373	92	374
rect	91	376	92	377
rect	91	379	92	380
rect	91	385	92	386
rect	92	1	93	2
rect	92	4	93	5
rect	92	7	93	8
rect	92	10	93	11
rect	92	13	93	14
rect	92	16	93	17
rect	92	19	93	20
rect	92	22	93	23
rect	92	25	93	26
rect	92	28	93	29
rect	92	31	93	32
rect	92	34	93	35
rect	92	37	93	38
rect	92	40	93	41
rect	92	43	93	44
rect	92	46	93	47
rect	92	49	93	50
rect	92	52	93	53
rect	92	55	93	56
rect	92	58	93	59
rect	92	61	93	62
rect	92	64	93	65
rect	92	67	93	68
rect	92	70	93	71
rect	92	73	93	74
rect	92	76	93	77
rect	92	79	93	80
rect	92	82	93	83
rect	92	85	93	86
rect	92	88	93	89
rect	92	91	93	92
rect	92	94	93	95
rect	92	97	93	98
rect	92	100	93	101
rect	92	103	93	104
rect	92	106	93	107
rect	92	109	93	110
rect	92	112	93	113
rect	92	115	93	116
rect	92	118	93	119
rect	92	121	93	122
rect	92	124	93	125
rect	92	127	93	128
rect	92	130	93	131
rect	92	133	93	134
rect	92	136	93	137
rect	92	139	93	140
rect	92	142	93	143
rect	92	145	93	146
rect	92	148	93	149
rect	92	151	93	152
rect	92	154	93	155
rect	92	157	93	158
rect	92	160	93	161
rect	92	163	93	164
rect	92	166	93	167
rect	92	169	93	170
rect	92	172	93	173
rect	92	175	93	176
rect	92	178	93	179
rect	92	181	93	182
rect	92	184	93	185
rect	92	187	93	188
rect	92	190	93	191
rect	92	193	93	194
rect	92	196	93	197
rect	92	199	93	200
rect	92	202	93	203
rect	92	205	93	206
rect	92	208	93	209
rect	92	211	93	212
rect	92	214	93	215
rect	92	217	93	218
rect	92	220	93	221
rect	92	223	93	224
rect	92	226	93	227
rect	92	229	93	230
rect	92	232	93	233
rect	92	235	93	236
rect	92	238	93	239
rect	92	241	93	242
rect	92	244	93	245
rect	92	247	93	248
rect	92	250	93	251
rect	92	253	93	254
rect	92	256	93	257
rect	92	259	93	260
rect	92	262	93	263
rect	92	265	93	266
rect	92	268	93	269
rect	92	271	93	272
rect	92	274	93	275
rect	92	277	93	278
rect	92	280	93	281
rect	92	283	93	284
rect	92	286	93	287
rect	92	289	93	290
rect	92	292	93	293
rect	92	295	93	296
rect	92	298	93	299
rect	92	301	93	302
rect	92	304	93	305
rect	92	307	93	308
rect	92	310	93	311
rect	92	313	93	314
rect	92	316	93	317
rect	92	319	93	320
rect	92	322	93	323
rect	92	325	93	326
rect	92	328	93	329
rect	92	331	93	332
rect	92	334	93	335
rect	92	337	93	338
rect	92	340	93	341
rect	92	343	93	344
rect	92	346	93	347
rect	92	349	93	350
rect	92	352	93	353
rect	92	355	93	356
rect	92	358	93	359
rect	92	361	93	362
rect	92	364	93	365
rect	92	367	93	368
rect	92	373	93	374
rect	92	376	93	377
rect	92	379	93	380
rect	92	385	93	386
rect	93	1	94	2
rect	93	4	94	5
rect	93	7	94	8
rect	93	10	94	11
rect	93	13	94	14
rect	93	16	94	17
rect	93	19	94	20
rect	93	22	94	23
rect	93	25	94	26
rect	93	28	94	29
rect	93	31	94	32
rect	93	34	94	35
rect	93	37	94	38
rect	93	40	94	41
rect	93	43	94	44
rect	93	46	94	47
rect	93	49	94	50
rect	93	52	94	53
rect	93	55	94	56
rect	93	58	94	59
rect	93	61	94	62
rect	93	64	94	65
rect	93	67	94	68
rect	93	70	94	71
rect	93	73	94	74
rect	93	76	94	77
rect	93	79	94	80
rect	93	82	94	83
rect	93	85	94	86
rect	93	88	94	89
rect	93	91	94	92
rect	93	94	94	95
rect	93	97	94	98
rect	93	100	94	101
rect	93	103	94	104
rect	93	106	94	107
rect	93	109	94	110
rect	93	112	94	113
rect	93	115	94	116
rect	93	118	94	119
rect	93	121	94	122
rect	93	124	94	125
rect	93	127	94	128
rect	93	130	94	131
rect	93	133	94	134
rect	93	136	94	137
rect	93	139	94	140
rect	93	142	94	143
rect	93	145	94	146
rect	93	148	94	149
rect	93	151	94	152
rect	93	154	94	155
rect	93	157	94	158
rect	93	160	94	161
rect	93	163	94	164
rect	93	166	94	167
rect	93	169	94	170
rect	93	172	94	173
rect	93	175	94	176
rect	93	178	94	179
rect	93	181	94	182
rect	93	184	94	185
rect	93	187	94	188
rect	93	190	94	191
rect	93	193	94	194
rect	93	196	94	197
rect	93	199	94	200
rect	93	202	94	203
rect	93	205	94	206
rect	93	208	94	209
rect	93	211	94	212
rect	93	214	94	215
rect	93	217	94	218
rect	93	220	94	221
rect	93	223	94	224
rect	93	226	94	227
rect	93	229	94	230
rect	93	232	94	233
rect	93	235	94	236
rect	93	238	94	239
rect	93	241	94	242
rect	93	244	94	245
rect	93	247	94	248
rect	93	250	94	251
rect	93	253	94	254
rect	93	256	94	257
rect	93	259	94	260
rect	93	262	94	263
rect	93	265	94	266
rect	93	268	94	269
rect	93	271	94	272
rect	93	274	94	275
rect	93	277	94	278
rect	93	280	94	281
rect	93	283	94	284
rect	93	286	94	287
rect	93	289	94	290
rect	93	292	94	293
rect	93	295	94	296
rect	93	298	94	299
rect	93	301	94	302
rect	93	304	94	305
rect	93	307	94	308
rect	93	310	94	311
rect	93	313	94	314
rect	93	316	94	317
rect	93	319	94	320
rect	93	322	94	323
rect	93	325	94	326
rect	93	328	94	329
rect	93	331	94	332
rect	93	334	94	335
rect	93	337	94	338
rect	93	340	94	341
rect	93	343	94	344
rect	93	346	94	347
rect	93	349	94	350
rect	93	352	94	353
rect	93	355	94	356
rect	93	358	94	359
rect	93	361	94	362
rect	93	364	94	365
rect	93	367	94	368
rect	93	373	94	374
rect	93	376	94	377
rect	93	379	94	380
rect	93	385	94	386
rect	94	1	95	2
rect	94	4	95	5
rect	94	7	95	8
rect	94	10	95	11
rect	94	13	95	14
rect	94	16	95	17
rect	94	19	95	20
rect	94	22	95	23
rect	94	25	95	26
rect	94	28	95	29
rect	94	31	95	32
rect	94	34	95	35
rect	94	37	95	38
rect	94	40	95	41
rect	94	43	95	44
rect	94	46	95	47
rect	94	49	95	50
rect	94	52	95	53
rect	94	55	95	56
rect	94	58	95	59
rect	94	61	95	62
rect	94	64	95	65
rect	94	67	95	68
rect	94	70	95	71
rect	94	73	95	74
rect	94	76	95	77
rect	94	79	95	80
rect	94	82	95	83
rect	94	85	95	86
rect	94	88	95	89
rect	94	91	95	92
rect	94	94	95	95
rect	94	97	95	98
rect	94	100	95	101
rect	94	103	95	104
rect	94	106	95	107
rect	94	109	95	110
rect	94	112	95	113
rect	94	115	95	116
rect	94	118	95	119
rect	94	121	95	122
rect	94	124	95	125
rect	94	127	95	128
rect	94	130	95	131
rect	94	133	95	134
rect	94	136	95	137
rect	94	139	95	140
rect	94	142	95	143
rect	94	145	95	146
rect	94	148	95	149
rect	94	151	95	152
rect	94	154	95	155
rect	94	157	95	158
rect	94	160	95	161
rect	94	163	95	164
rect	94	166	95	167
rect	94	169	95	170
rect	94	172	95	173
rect	94	175	95	176
rect	94	178	95	179
rect	94	181	95	182
rect	94	184	95	185
rect	94	187	95	188
rect	94	190	95	191
rect	94	193	95	194
rect	94	196	95	197
rect	94	199	95	200
rect	94	202	95	203
rect	94	205	95	206
rect	94	208	95	209
rect	94	211	95	212
rect	94	214	95	215
rect	94	217	95	218
rect	94	220	95	221
rect	94	223	95	224
rect	94	226	95	227
rect	94	229	95	230
rect	94	232	95	233
rect	94	235	95	236
rect	94	238	95	239
rect	94	241	95	242
rect	94	244	95	245
rect	94	247	95	248
rect	94	250	95	251
rect	94	253	95	254
rect	94	256	95	257
rect	94	259	95	260
rect	94	262	95	263
rect	94	265	95	266
rect	94	268	95	269
rect	94	271	95	272
rect	94	274	95	275
rect	94	277	95	278
rect	94	280	95	281
rect	94	283	95	284
rect	94	286	95	287
rect	94	289	95	290
rect	94	292	95	293
rect	94	295	95	296
rect	94	298	95	299
rect	94	301	95	302
rect	94	304	95	305
rect	94	307	95	308
rect	94	310	95	311
rect	94	313	95	314
rect	94	316	95	317
rect	94	319	95	320
rect	94	322	95	323
rect	94	325	95	326
rect	94	328	95	329
rect	94	331	95	332
rect	94	334	95	335
rect	94	337	95	338
rect	94	340	95	341
rect	94	343	95	344
rect	94	346	95	347
rect	94	349	95	350
rect	94	352	95	353
rect	94	355	95	356
rect	94	358	95	359
rect	94	361	95	362
rect	94	364	95	365
rect	94	367	95	368
rect	94	373	95	374
rect	94	376	95	377
rect	94	379	95	380
rect	94	385	95	386
rect	95	1	96	2
rect	95	4	96	5
rect	95	7	96	8
rect	95	10	96	11
rect	95	13	96	14
rect	95	16	96	17
rect	95	19	96	20
rect	95	22	96	23
rect	95	25	96	26
rect	95	28	96	29
rect	95	31	96	32
rect	95	34	96	35
rect	95	37	96	38
rect	95	40	96	41
rect	95	43	96	44
rect	95	46	96	47
rect	95	49	96	50
rect	95	52	96	53
rect	95	55	96	56
rect	95	58	96	59
rect	95	61	96	62
rect	95	64	96	65
rect	95	67	96	68
rect	95	70	96	71
rect	95	73	96	74
rect	95	76	96	77
rect	95	79	96	80
rect	95	82	96	83
rect	95	85	96	86
rect	95	88	96	89
rect	95	91	96	92
rect	95	94	96	95
rect	95	97	96	98
rect	95	100	96	101
rect	95	103	96	104
rect	95	106	96	107
rect	95	109	96	110
rect	95	112	96	113
rect	95	115	96	116
rect	95	118	96	119
rect	95	121	96	122
rect	95	124	96	125
rect	95	127	96	128
rect	95	130	96	131
rect	95	133	96	134
rect	95	136	96	137
rect	95	139	96	140
rect	95	142	96	143
rect	95	145	96	146
rect	95	148	96	149
rect	95	151	96	152
rect	95	154	96	155
rect	95	157	96	158
rect	95	160	96	161
rect	95	163	96	164
rect	95	166	96	167
rect	95	169	96	170
rect	95	172	96	173
rect	95	175	96	176
rect	95	178	96	179
rect	95	181	96	182
rect	95	184	96	185
rect	95	187	96	188
rect	95	190	96	191
rect	95	193	96	194
rect	95	196	96	197
rect	95	199	96	200
rect	95	202	96	203
rect	95	205	96	206
rect	95	208	96	209
rect	95	211	96	212
rect	95	214	96	215
rect	95	217	96	218
rect	95	220	96	221
rect	95	223	96	224
rect	95	226	96	227
rect	95	229	96	230
rect	95	232	96	233
rect	95	235	96	236
rect	95	238	96	239
rect	95	241	96	242
rect	95	244	96	245
rect	95	247	96	248
rect	95	250	96	251
rect	95	253	96	254
rect	95	256	96	257
rect	95	259	96	260
rect	95	262	96	263
rect	95	265	96	266
rect	95	268	96	269
rect	95	271	96	272
rect	95	274	96	275
rect	95	277	96	278
rect	95	280	96	281
rect	95	283	96	284
rect	95	286	96	287
rect	95	289	96	290
rect	95	292	96	293
rect	95	295	96	296
rect	95	298	96	299
rect	95	301	96	302
rect	95	304	96	305
rect	95	307	96	308
rect	95	310	96	311
rect	95	313	96	314
rect	95	316	96	317
rect	95	319	96	320
rect	95	322	96	323
rect	95	325	96	326
rect	95	328	96	329
rect	95	331	96	332
rect	95	334	96	335
rect	95	337	96	338
rect	95	340	96	341
rect	95	343	96	344
rect	95	346	96	347
rect	95	349	96	350
rect	95	352	96	353
rect	95	355	96	356
rect	95	358	96	359
rect	95	361	96	362
rect	95	364	96	365
rect	95	367	96	368
rect	95	373	96	374
rect	95	376	96	377
rect	95	379	96	380
rect	95	385	96	386
rect	96	1	97	2
rect	96	4	97	5
rect	96	7	97	8
rect	96	10	97	11
rect	96	13	97	14
rect	96	16	97	17
rect	96	19	97	20
rect	96	22	97	23
rect	96	25	97	26
rect	96	28	97	29
rect	96	31	97	32
rect	96	34	97	35
rect	96	37	97	38
rect	96	40	97	41
rect	96	43	97	44
rect	96	46	97	47
rect	96	49	97	50
rect	96	52	97	53
rect	96	55	97	56
rect	96	58	97	59
rect	96	61	97	62
rect	96	64	97	65
rect	96	67	97	68
rect	96	70	97	71
rect	96	73	97	74
rect	96	76	97	77
rect	96	79	97	80
rect	96	82	97	83
rect	96	85	97	86
rect	96	88	97	89
rect	96	91	97	92
rect	96	94	97	95
rect	96	97	97	98
rect	96	100	97	101
rect	96	103	97	104
rect	96	106	97	107
rect	96	109	97	110
rect	96	112	97	113
rect	96	115	97	116
rect	96	118	97	119
rect	96	121	97	122
rect	96	124	97	125
rect	96	127	97	128
rect	96	130	97	131
rect	96	133	97	134
rect	96	136	97	137
rect	96	139	97	140
rect	96	142	97	143
rect	96	145	97	146
rect	96	148	97	149
rect	96	151	97	152
rect	96	154	97	155
rect	96	157	97	158
rect	96	160	97	161
rect	96	163	97	164
rect	96	166	97	167
rect	96	169	97	170
rect	96	172	97	173
rect	96	175	97	176
rect	96	178	97	179
rect	96	181	97	182
rect	96	184	97	185
rect	96	187	97	188
rect	96	190	97	191
rect	96	193	97	194
rect	96	196	97	197
rect	96	199	97	200
rect	96	202	97	203
rect	96	205	97	206
rect	96	208	97	209
rect	96	211	97	212
rect	96	214	97	215
rect	96	217	97	218
rect	96	220	97	221
rect	96	223	97	224
rect	96	226	97	227
rect	96	229	97	230
rect	96	232	97	233
rect	96	235	97	236
rect	96	238	97	239
rect	96	241	97	242
rect	96	244	97	245
rect	96	247	97	248
rect	96	250	97	251
rect	96	253	97	254
rect	96	256	97	257
rect	96	259	97	260
rect	96	262	97	263
rect	96	265	97	266
rect	96	268	97	269
rect	96	271	97	272
rect	96	274	97	275
rect	96	277	97	278
rect	96	280	97	281
rect	96	283	97	284
rect	96	286	97	287
rect	96	289	97	290
rect	96	292	97	293
rect	96	295	97	296
rect	96	298	97	299
rect	96	301	97	302
rect	96	304	97	305
rect	96	307	97	308
rect	96	310	97	311
rect	96	313	97	314
rect	96	316	97	317
rect	96	319	97	320
rect	96	322	97	323
rect	96	325	97	326
rect	96	328	97	329
rect	96	331	97	332
rect	96	334	97	335
rect	96	337	97	338
rect	96	340	97	341
rect	96	343	97	344
rect	96	346	97	347
rect	96	349	97	350
rect	96	352	97	353
rect	96	355	97	356
rect	96	358	97	359
rect	96	361	97	362
rect	96	364	97	365
rect	96	367	97	368
rect	96	373	97	374
rect	96	376	97	377
rect	96	379	97	380
rect	96	385	97	386
rect	97	1	98	2
rect	97	4	98	5
rect	97	7	98	8
rect	97	10	98	11
rect	97	13	98	14
rect	97	16	98	17
rect	97	19	98	20
rect	97	22	98	23
rect	97	25	98	26
rect	97	28	98	29
rect	97	31	98	32
rect	97	34	98	35
rect	97	37	98	38
rect	97	40	98	41
rect	97	43	98	44
rect	97	46	98	47
rect	97	49	98	50
rect	97	52	98	53
rect	97	55	98	56
rect	97	58	98	59
rect	97	61	98	62
rect	97	64	98	65
rect	97	67	98	68
rect	97	70	98	71
rect	97	73	98	74
rect	97	76	98	77
rect	97	79	98	80
rect	97	82	98	83
rect	97	85	98	86
rect	97	88	98	89
rect	97	91	98	92
rect	97	94	98	95
rect	97	97	98	98
rect	97	100	98	101
rect	97	103	98	104
rect	97	106	98	107
rect	97	109	98	110
rect	97	112	98	113
rect	97	115	98	116
rect	97	118	98	119
rect	97	121	98	122
rect	97	124	98	125
rect	97	127	98	128
rect	97	130	98	131
rect	97	133	98	134
rect	97	136	98	137
rect	97	139	98	140
rect	97	142	98	143
rect	97	145	98	146
rect	97	148	98	149
rect	97	151	98	152
rect	97	154	98	155
rect	97	157	98	158
rect	97	160	98	161
rect	97	163	98	164
rect	97	166	98	167
rect	97	169	98	170
rect	97	172	98	173
rect	97	175	98	176
rect	97	178	98	179
rect	97	181	98	182
rect	97	184	98	185
rect	97	187	98	188
rect	97	190	98	191
rect	97	193	98	194
rect	97	196	98	197
rect	97	199	98	200
rect	97	202	98	203
rect	97	205	98	206
rect	97	208	98	209
rect	97	211	98	212
rect	97	214	98	215
rect	97	217	98	218
rect	97	220	98	221
rect	97	223	98	224
rect	97	226	98	227
rect	97	229	98	230
rect	97	232	98	233
rect	97	235	98	236
rect	97	238	98	239
rect	97	241	98	242
rect	97	244	98	245
rect	97	247	98	248
rect	97	250	98	251
rect	97	253	98	254
rect	97	256	98	257
rect	97	259	98	260
rect	97	262	98	263
rect	97	265	98	266
rect	97	268	98	269
rect	97	271	98	272
rect	97	274	98	275
rect	97	277	98	278
rect	97	280	98	281
rect	97	283	98	284
rect	97	286	98	287
rect	97	289	98	290
rect	97	292	98	293
rect	97	295	98	296
rect	97	298	98	299
rect	97	301	98	302
rect	97	304	98	305
rect	97	307	98	308
rect	97	310	98	311
rect	97	313	98	314
rect	97	316	98	317
rect	97	319	98	320
rect	97	322	98	323
rect	97	325	98	326
rect	97	328	98	329
rect	97	331	98	332
rect	97	334	98	335
rect	97	337	98	338
rect	97	340	98	341
rect	97	343	98	344
rect	97	346	98	347
rect	97	349	98	350
rect	97	352	98	353
rect	97	355	98	356
rect	97	358	98	359
rect	97	361	98	362
rect	97	364	98	365
rect	97	367	98	368
rect	97	373	98	374
rect	97	376	98	377
rect	97	379	98	380
rect	97	385	98	386
rect	98	1	99	2
rect	98	4	99	5
rect	98	7	99	8
rect	98	10	99	11
rect	98	13	99	14
rect	98	16	99	17
rect	98	19	99	20
rect	98	22	99	23
rect	98	25	99	26
rect	98	28	99	29
rect	98	31	99	32
rect	98	34	99	35
rect	98	37	99	38
rect	98	40	99	41
rect	98	43	99	44
rect	98	46	99	47
rect	98	49	99	50
rect	98	52	99	53
rect	98	55	99	56
rect	98	58	99	59
rect	98	61	99	62
rect	98	64	99	65
rect	98	67	99	68
rect	98	70	99	71
rect	98	73	99	74
rect	98	76	99	77
rect	98	79	99	80
rect	98	82	99	83
rect	98	85	99	86
rect	98	88	99	89
rect	98	91	99	92
rect	98	94	99	95
rect	98	97	99	98
rect	98	100	99	101
rect	98	103	99	104
rect	98	106	99	107
rect	98	109	99	110
rect	98	112	99	113
rect	98	115	99	116
rect	98	118	99	119
rect	98	121	99	122
rect	98	124	99	125
rect	98	127	99	128
rect	98	130	99	131
rect	98	133	99	134
rect	98	136	99	137
rect	98	139	99	140
rect	98	142	99	143
rect	98	145	99	146
rect	98	148	99	149
rect	98	151	99	152
rect	98	154	99	155
rect	98	157	99	158
rect	98	160	99	161
rect	98	163	99	164
rect	98	166	99	167
rect	98	169	99	170
rect	98	172	99	173
rect	98	175	99	176
rect	98	178	99	179
rect	98	181	99	182
rect	98	184	99	185
rect	98	187	99	188
rect	98	190	99	191
rect	98	193	99	194
rect	98	196	99	197
rect	98	199	99	200
rect	98	202	99	203
rect	98	205	99	206
rect	98	208	99	209
rect	98	211	99	212
rect	98	214	99	215
rect	98	217	99	218
rect	98	220	99	221
rect	98	223	99	224
rect	98	226	99	227
rect	98	229	99	230
rect	98	232	99	233
rect	98	235	99	236
rect	98	238	99	239
rect	98	241	99	242
rect	98	244	99	245
rect	98	247	99	248
rect	98	250	99	251
rect	98	253	99	254
rect	98	256	99	257
rect	98	259	99	260
rect	98	262	99	263
rect	98	265	99	266
rect	98	268	99	269
rect	98	271	99	272
rect	98	274	99	275
rect	98	277	99	278
rect	98	280	99	281
rect	98	283	99	284
rect	98	286	99	287
rect	98	289	99	290
rect	98	292	99	293
rect	98	295	99	296
rect	98	298	99	299
rect	98	301	99	302
rect	98	304	99	305
rect	98	307	99	308
rect	98	310	99	311
rect	98	313	99	314
rect	98	316	99	317
rect	98	319	99	320
rect	98	322	99	323
rect	98	325	99	326
rect	98	328	99	329
rect	98	331	99	332
rect	98	334	99	335
rect	98	337	99	338
rect	98	340	99	341
rect	98	343	99	344
rect	98	346	99	347
rect	98	349	99	350
rect	98	352	99	353
rect	98	355	99	356
rect	98	358	99	359
rect	98	361	99	362
rect	98	364	99	365
rect	98	367	99	368
rect	98	373	99	374
rect	98	376	99	377
rect	98	379	99	380
rect	98	385	99	386
rect	99	1	100	2
rect	99	4	100	5
rect	99	7	100	8
rect	99	10	100	11
rect	99	13	100	14
rect	99	16	100	17
rect	99	19	100	20
rect	99	22	100	23
rect	99	25	100	26
rect	99	28	100	29
rect	99	31	100	32
rect	99	34	100	35
rect	99	37	100	38
rect	99	40	100	41
rect	99	43	100	44
rect	99	46	100	47
rect	99	49	100	50
rect	99	52	100	53
rect	99	55	100	56
rect	99	58	100	59
rect	99	61	100	62
rect	99	64	100	65
rect	99	67	100	68
rect	99	70	100	71
rect	99	73	100	74
rect	99	76	100	77
rect	99	79	100	80
rect	99	82	100	83
rect	99	85	100	86
rect	99	88	100	89
rect	99	91	100	92
rect	99	94	100	95
rect	99	97	100	98
rect	99	100	100	101
rect	99	103	100	104
rect	99	106	100	107
rect	99	109	100	110
rect	99	112	100	113
rect	99	115	100	116
rect	99	118	100	119
rect	99	121	100	122
rect	99	124	100	125
rect	99	127	100	128
rect	99	130	100	131
rect	99	133	100	134
rect	99	136	100	137
rect	99	139	100	140
rect	99	142	100	143
rect	99	145	100	146
rect	99	148	100	149
rect	99	151	100	152
rect	99	154	100	155
rect	99	157	100	158
rect	99	160	100	161
rect	99	163	100	164
rect	99	166	100	167
rect	99	169	100	170
rect	99	172	100	173
rect	99	175	100	176
rect	99	178	100	179
rect	99	181	100	182
rect	99	184	100	185
rect	99	187	100	188
rect	99	190	100	191
rect	99	193	100	194
rect	99	196	100	197
rect	99	199	100	200
rect	99	202	100	203
rect	99	205	100	206
rect	99	208	100	209
rect	99	211	100	212
rect	99	214	100	215
rect	99	217	100	218
rect	99	220	100	221
rect	99	223	100	224
rect	99	226	100	227
rect	99	229	100	230
rect	99	232	100	233
rect	99	235	100	236
rect	99	238	100	239
rect	99	241	100	242
rect	99	244	100	245
rect	99	247	100	248
rect	99	250	100	251
rect	99	253	100	254
rect	99	256	100	257
rect	99	259	100	260
rect	99	262	100	263
rect	99	265	100	266
rect	99	268	100	269
rect	99	271	100	272
rect	99	274	100	275
rect	99	277	100	278
rect	99	280	100	281
rect	99	283	100	284
rect	99	286	100	287
rect	99	289	100	290
rect	99	292	100	293
rect	99	295	100	296
rect	99	298	100	299
rect	99	301	100	302
rect	99	304	100	305
rect	99	307	100	308
rect	99	310	100	311
rect	99	313	100	314
rect	99	316	100	317
rect	99	319	100	320
rect	99	322	100	323
rect	99	325	100	326
rect	99	328	100	329
rect	99	331	100	332
rect	99	334	100	335
rect	99	337	100	338
rect	99	340	100	341
rect	99	343	100	344
rect	99	346	100	347
rect	99	349	100	350
rect	99	352	100	353
rect	99	355	100	356
rect	99	358	100	359
rect	99	361	100	362
rect	99	364	100	365
rect	99	367	100	368
rect	99	373	100	374
rect	99	376	100	377
rect	99	379	100	380
rect	99	385	100	386
rect	100	1	101	2
rect	100	4	101	5
rect	100	7	101	8
rect	100	10	101	11
rect	100	13	101	14
rect	100	16	101	17
rect	100	19	101	20
rect	100	22	101	23
rect	100	25	101	26
rect	100	28	101	29
rect	100	31	101	32
rect	100	34	101	35
rect	100	37	101	38
rect	100	40	101	41
rect	100	43	101	44
rect	100	46	101	47
rect	100	49	101	50
rect	100	52	101	53
rect	100	55	101	56
rect	100	58	101	59
rect	100	61	101	62
rect	100	64	101	65
rect	100	67	101	68
rect	100	70	101	71
rect	100	73	101	74
rect	100	76	101	77
rect	100	79	101	80
rect	100	82	101	83
rect	100	85	101	86
rect	100	88	101	89
rect	100	91	101	92
rect	100	94	101	95
rect	100	97	101	98
rect	100	100	101	101
rect	100	103	101	104
rect	100	106	101	107
rect	100	109	101	110
rect	100	112	101	113
rect	100	115	101	116
rect	100	118	101	119
rect	100	121	101	122
rect	100	124	101	125
rect	100	127	101	128
rect	100	130	101	131
rect	100	133	101	134
rect	100	136	101	137
rect	100	139	101	140
rect	100	142	101	143
rect	100	145	101	146
rect	100	148	101	149
rect	100	151	101	152
rect	100	154	101	155
rect	100	157	101	158
rect	100	160	101	161
rect	100	163	101	164
rect	100	166	101	167
rect	100	169	101	170
rect	100	172	101	173
rect	100	175	101	176
rect	100	178	101	179
rect	100	181	101	182
rect	100	184	101	185
rect	100	187	101	188
rect	100	190	101	191
rect	100	193	101	194
rect	100	196	101	197
rect	100	199	101	200
rect	100	202	101	203
rect	100	205	101	206
rect	100	208	101	209
rect	100	211	101	212
rect	100	214	101	215
rect	100	217	101	218
rect	100	220	101	221
rect	100	223	101	224
rect	100	226	101	227
rect	100	229	101	230
rect	100	232	101	233
rect	100	235	101	236
rect	100	238	101	239
rect	100	241	101	242
rect	100	244	101	245
rect	100	247	101	248
rect	100	250	101	251
rect	100	253	101	254
rect	100	256	101	257
rect	100	259	101	260
rect	100	262	101	263
rect	100	265	101	266
rect	100	268	101	269
rect	100	271	101	272
rect	100	274	101	275
rect	100	277	101	278
rect	100	280	101	281
rect	100	283	101	284
rect	100	286	101	287
rect	100	289	101	290
rect	100	292	101	293
rect	100	295	101	296
rect	100	298	101	299
rect	100	301	101	302
rect	100	304	101	305
rect	100	307	101	308
rect	100	310	101	311
rect	100	313	101	314
rect	100	316	101	317
rect	100	319	101	320
rect	100	322	101	323
rect	100	325	101	326
rect	100	328	101	329
rect	100	331	101	332
rect	100	334	101	335
rect	100	337	101	338
rect	100	340	101	341
rect	100	343	101	344
rect	100	346	101	347
rect	100	349	101	350
rect	100	352	101	353
rect	100	355	101	356
rect	100	358	101	359
rect	100	361	101	362
rect	100	364	101	365
rect	100	367	101	368
rect	100	373	101	374
rect	100	376	101	377
rect	100	379	101	380
rect	100	385	101	386
rect	101	1	102	2
rect	101	4	102	5
rect	101	7	102	8
rect	101	10	102	11
rect	101	13	102	14
rect	101	16	102	17
rect	101	19	102	20
rect	101	22	102	23
rect	101	25	102	26
rect	101	28	102	29
rect	101	31	102	32
rect	101	34	102	35
rect	101	37	102	38
rect	101	40	102	41
rect	101	43	102	44
rect	101	46	102	47
rect	101	49	102	50
rect	101	52	102	53
rect	101	55	102	56
rect	101	58	102	59
rect	101	61	102	62
rect	101	64	102	65
rect	101	67	102	68
rect	101	70	102	71
rect	101	73	102	74
rect	101	76	102	77
rect	101	79	102	80
rect	101	82	102	83
rect	101	85	102	86
rect	101	88	102	89
rect	101	91	102	92
rect	101	94	102	95
rect	101	97	102	98
rect	101	100	102	101
rect	101	103	102	104
rect	101	106	102	107
rect	101	109	102	110
rect	101	112	102	113
rect	101	115	102	116
rect	101	118	102	119
rect	101	121	102	122
rect	101	124	102	125
rect	101	127	102	128
rect	101	130	102	131
rect	101	133	102	134
rect	101	136	102	137
rect	101	139	102	140
rect	101	142	102	143
rect	101	145	102	146
rect	101	148	102	149
rect	101	151	102	152
rect	101	154	102	155
rect	101	157	102	158
rect	101	160	102	161
rect	101	163	102	164
rect	101	166	102	167
rect	101	169	102	170
rect	101	172	102	173
rect	101	175	102	176
rect	101	178	102	179
rect	101	181	102	182
rect	101	184	102	185
rect	101	187	102	188
rect	101	190	102	191
rect	101	193	102	194
rect	101	196	102	197
rect	101	199	102	200
rect	101	202	102	203
rect	101	205	102	206
rect	101	208	102	209
rect	101	211	102	212
rect	101	214	102	215
rect	101	217	102	218
rect	101	220	102	221
rect	101	223	102	224
rect	101	226	102	227
rect	101	229	102	230
rect	101	232	102	233
rect	101	235	102	236
rect	101	238	102	239
rect	101	241	102	242
rect	101	244	102	245
rect	101	247	102	248
rect	101	250	102	251
rect	101	253	102	254
rect	101	256	102	257
rect	101	259	102	260
rect	101	262	102	263
rect	101	265	102	266
rect	101	268	102	269
rect	101	271	102	272
rect	101	274	102	275
rect	101	277	102	278
rect	101	280	102	281
rect	101	283	102	284
rect	101	286	102	287
rect	101	289	102	290
rect	101	292	102	293
rect	101	295	102	296
rect	101	298	102	299
rect	101	301	102	302
rect	101	304	102	305
rect	101	307	102	308
rect	101	310	102	311
rect	101	313	102	314
rect	101	316	102	317
rect	101	319	102	320
rect	101	322	102	323
rect	101	325	102	326
rect	101	328	102	329
rect	101	331	102	332
rect	101	334	102	335
rect	101	337	102	338
rect	101	340	102	341
rect	101	343	102	344
rect	101	346	102	347
rect	101	349	102	350
rect	101	352	102	353
rect	101	355	102	356
rect	101	358	102	359
rect	101	361	102	362
rect	101	364	102	365
rect	101	367	102	368
rect	101	373	102	374
rect	101	376	102	377
rect	101	379	102	380
rect	101	385	102	386
rect	102	1	103	2
rect	102	4	103	5
rect	102	7	103	8
rect	102	10	103	11
rect	102	13	103	14
rect	102	16	103	17
rect	102	19	103	20
rect	102	22	103	23
rect	102	25	103	26
rect	102	28	103	29
rect	102	31	103	32
rect	102	34	103	35
rect	102	37	103	38
rect	102	40	103	41
rect	102	43	103	44
rect	102	46	103	47
rect	102	49	103	50
rect	102	52	103	53
rect	102	55	103	56
rect	102	58	103	59
rect	102	61	103	62
rect	102	64	103	65
rect	102	67	103	68
rect	102	70	103	71
rect	102	73	103	74
rect	102	76	103	77
rect	102	79	103	80
rect	102	82	103	83
rect	102	85	103	86
rect	102	88	103	89
rect	102	91	103	92
rect	102	94	103	95
rect	102	97	103	98
rect	102	100	103	101
rect	102	103	103	104
rect	102	106	103	107
rect	102	109	103	110
rect	102	112	103	113
rect	102	115	103	116
rect	102	118	103	119
rect	102	121	103	122
rect	102	124	103	125
rect	102	127	103	128
rect	102	130	103	131
rect	102	133	103	134
rect	102	136	103	137
rect	102	139	103	140
rect	102	142	103	143
rect	102	145	103	146
rect	102	148	103	149
rect	102	151	103	152
rect	102	154	103	155
rect	102	157	103	158
rect	102	160	103	161
rect	102	163	103	164
rect	102	166	103	167
rect	102	169	103	170
rect	102	172	103	173
rect	102	175	103	176
rect	102	178	103	179
rect	102	181	103	182
rect	102	184	103	185
rect	102	187	103	188
rect	102	190	103	191
rect	102	193	103	194
rect	102	196	103	197
rect	102	199	103	200
rect	102	202	103	203
rect	102	205	103	206
rect	102	208	103	209
rect	102	211	103	212
rect	102	214	103	215
rect	102	217	103	218
rect	102	220	103	221
rect	102	223	103	224
rect	102	226	103	227
rect	102	229	103	230
rect	102	232	103	233
rect	102	235	103	236
rect	102	238	103	239
rect	102	241	103	242
rect	102	244	103	245
rect	102	247	103	248
rect	102	250	103	251
rect	102	253	103	254
rect	102	256	103	257
rect	102	259	103	260
rect	102	262	103	263
rect	102	265	103	266
rect	102	268	103	269
rect	102	271	103	272
rect	102	274	103	275
rect	102	277	103	278
rect	102	280	103	281
rect	102	283	103	284
rect	102	286	103	287
rect	102	289	103	290
rect	102	292	103	293
rect	102	295	103	296
rect	102	298	103	299
rect	102	301	103	302
rect	102	304	103	305
rect	102	307	103	308
rect	102	310	103	311
rect	102	313	103	314
rect	102	316	103	317
rect	102	319	103	320
rect	102	322	103	323
rect	102	325	103	326
rect	102	328	103	329
rect	102	331	103	332
rect	102	334	103	335
rect	102	337	103	338
rect	102	340	103	341
rect	102	343	103	344
rect	102	346	103	347
rect	102	349	103	350
rect	102	352	103	353
rect	102	355	103	356
rect	102	358	103	359
rect	102	361	103	362
rect	102	364	103	365
rect	102	367	103	368
rect	102	373	103	374
rect	102	376	103	377
rect	102	379	103	380
rect	102	385	103	386
rect	103	1	104	2
rect	103	4	104	5
rect	103	7	104	8
rect	103	10	104	11
rect	103	13	104	14
rect	103	16	104	17
rect	103	19	104	20
rect	103	22	104	23
rect	103	25	104	26
rect	103	28	104	29
rect	103	31	104	32
rect	103	34	104	35
rect	103	37	104	38
rect	103	40	104	41
rect	103	43	104	44
rect	103	46	104	47
rect	103	49	104	50
rect	103	52	104	53
rect	103	55	104	56
rect	103	58	104	59
rect	103	61	104	62
rect	103	64	104	65
rect	103	67	104	68
rect	103	70	104	71
rect	103	73	104	74
rect	103	76	104	77
rect	103	79	104	80
rect	103	82	104	83
rect	103	85	104	86
rect	103	88	104	89
rect	103	91	104	92
rect	103	94	104	95
rect	103	97	104	98
rect	103	100	104	101
rect	103	103	104	104
rect	103	106	104	107
rect	103	109	104	110
rect	103	112	104	113
rect	103	115	104	116
rect	103	118	104	119
rect	103	121	104	122
rect	103	124	104	125
rect	103	127	104	128
rect	103	130	104	131
rect	103	133	104	134
rect	103	136	104	137
rect	103	139	104	140
rect	103	142	104	143
rect	103	145	104	146
rect	103	148	104	149
rect	103	151	104	152
rect	103	154	104	155
rect	103	157	104	158
rect	103	160	104	161
rect	103	163	104	164
rect	103	166	104	167
rect	103	169	104	170
rect	103	172	104	173
rect	103	175	104	176
rect	103	178	104	179
rect	103	181	104	182
rect	103	184	104	185
rect	103	187	104	188
rect	103	190	104	191
rect	103	193	104	194
rect	103	196	104	197
rect	103	199	104	200
rect	103	202	104	203
rect	103	205	104	206
rect	103	208	104	209
rect	103	211	104	212
rect	103	214	104	215
rect	103	217	104	218
rect	103	220	104	221
rect	103	223	104	224
rect	103	226	104	227
rect	103	229	104	230
rect	103	232	104	233
rect	103	235	104	236
rect	103	238	104	239
rect	103	241	104	242
rect	103	244	104	245
rect	103	247	104	248
rect	103	250	104	251
rect	103	253	104	254
rect	103	256	104	257
rect	103	259	104	260
rect	103	262	104	263
rect	103	265	104	266
rect	103	268	104	269
rect	103	271	104	272
rect	103	274	104	275
rect	103	277	104	278
rect	103	280	104	281
rect	103	283	104	284
rect	103	286	104	287
rect	103	289	104	290
rect	103	292	104	293
rect	103	295	104	296
rect	103	298	104	299
rect	103	301	104	302
rect	103	304	104	305
rect	103	307	104	308
rect	103	310	104	311
rect	103	313	104	314
rect	103	316	104	317
rect	103	319	104	320
rect	103	322	104	323
rect	103	325	104	326
rect	103	328	104	329
rect	103	331	104	332
rect	103	334	104	335
rect	103	337	104	338
rect	103	340	104	341
rect	103	343	104	344
rect	103	346	104	347
rect	103	349	104	350
rect	103	352	104	353
rect	103	355	104	356
rect	103	358	104	359
rect	103	361	104	362
rect	103	364	104	365
rect	103	367	104	368
rect	103	373	104	374
rect	103	376	104	377
rect	103	379	104	380
rect	103	385	104	386
rect	104	1	105	2
rect	104	4	105	5
rect	104	7	105	8
rect	104	10	105	11
rect	104	13	105	14
rect	104	16	105	17
rect	104	19	105	20
rect	104	22	105	23
rect	104	25	105	26
rect	104	28	105	29
rect	104	31	105	32
rect	104	34	105	35
rect	104	37	105	38
rect	104	40	105	41
rect	104	43	105	44
rect	104	46	105	47
rect	104	49	105	50
rect	104	52	105	53
rect	104	55	105	56
rect	104	58	105	59
rect	104	61	105	62
rect	104	64	105	65
rect	104	67	105	68
rect	104	70	105	71
rect	104	73	105	74
rect	104	76	105	77
rect	104	79	105	80
rect	104	82	105	83
rect	104	85	105	86
rect	104	88	105	89
rect	104	91	105	92
rect	104	94	105	95
rect	104	97	105	98
rect	104	100	105	101
rect	104	103	105	104
rect	104	106	105	107
rect	104	109	105	110
rect	104	112	105	113
rect	104	115	105	116
rect	104	118	105	119
rect	104	121	105	122
rect	104	124	105	125
rect	104	127	105	128
rect	104	130	105	131
rect	104	133	105	134
rect	104	136	105	137
rect	104	139	105	140
rect	104	142	105	143
rect	104	145	105	146
rect	104	148	105	149
rect	104	151	105	152
rect	104	154	105	155
rect	104	157	105	158
rect	104	160	105	161
rect	104	163	105	164
rect	104	166	105	167
rect	104	169	105	170
rect	104	172	105	173
rect	104	175	105	176
rect	104	178	105	179
rect	104	181	105	182
rect	104	184	105	185
rect	104	187	105	188
rect	104	190	105	191
rect	104	193	105	194
rect	104	196	105	197
rect	104	199	105	200
rect	104	202	105	203
rect	104	205	105	206
rect	104	208	105	209
rect	104	211	105	212
rect	104	214	105	215
rect	104	217	105	218
rect	104	220	105	221
rect	104	223	105	224
rect	104	226	105	227
rect	104	229	105	230
rect	104	232	105	233
rect	104	235	105	236
rect	104	238	105	239
rect	104	241	105	242
rect	104	244	105	245
rect	104	247	105	248
rect	104	250	105	251
rect	104	253	105	254
rect	104	256	105	257
rect	104	259	105	260
rect	104	262	105	263
rect	104	265	105	266
rect	104	268	105	269
rect	104	271	105	272
rect	104	274	105	275
rect	104	277	105	278
rect	104	280	105	281
rect	104	283	105	284
rect	104	286	105	287
rect	104	289	105	290
rect	104	292	105	293
rect	104	295	105	296
rect	104	298	105	299
rect	104	301	105	302
rect	104	304	105	305
rect	104	307	105	308
rect	104	310	105	311
rect	104	313	105	314
rect	104	316	105	317
rect	104	319	105	320
rect	104	322	105	323
rect	104	325	105	326
rect	104	328	105	329
rect	104	331	105	332
rect	104	334	105	335
rect	104	337	105	338
rect	104	340	105	341
rect	104	343	105	344
rect	104	346	105	347
rect	104	349	105	350
rect	104	352	105	353
rect	104	355	105	356
rect	104	358	105	359
rect	104	361	105	362
rect	104	364	105	365
rect	104	367	105	368
rect	104	373	105	374
rect	104	376	105	377
rect	104	379	105	380
rect	104	385	105	386
rect	105	1	106	2
rect	105	4	106	5
rect	105	7	106	8
rect	105	10	106	11
rect	105	13	106	14
rect	105	16	106	17
rect	105	19	106	20
rect	105	22	106	23
rect	105	25	106	26
rect	105	28	106	29
rect	105	31	106	32
rect	105	34	106	35
rect	105	37	106	38
rect	105	40	106	41
rect	105	43	106	44
rect	105	46	106	47
rect	105	49	106	50
rect	105	52	106	53
rect	105	55	106	56
rect	105	58	106	59
rect	105	61	106	62
rect	105	64	106	65
rect	105	67	106	68
rect	105	70	106	71
rect	105	73	106	74
rect	105	76	106	77
rect	105	79	106	80
rect	105	82	106	83
rect	105	85	106	86
rect	105	88	106	89
rect	105	91	106	92
rect	105	94	106	95
rect	105	97	106	98
rect	105	100	106	101
rect	105	103	106	104
rect	105	106	106	107
rect	105	109	106	110
rect	105	112	106	113
rect	105	115	106	116
rect	105	118	106	119
rect	105	121	106	122
rect	105	124	106	125
rect	105	127	106	128
rect	105	130	106	131
rect	105	133	106	134
rect	105	136	106	137
rect	105	139	106	140
rect	105	142	106	143
rect	105	145	106	146
rect	105	148	106	149
rect	105	151	106	152
rect	105	154	106	155
rect	105	157	106	158
rect	105	160	106	161
rect	105	163	106	164
rect	105	166	106	167
rect	105	169	106	170
rect	105	172	106	173
rect	105	175	106	176
rect	105	178	106	179
rect	105	181	106	182
rect	105	184	106	185
rect	105	187	106	188
rect	105	190	106	191
rect	105	193	106	194
rect	105	196	106	197
rect	105	199	106	200
rect	105	202	106	203
rect	105	205	106	206
rect	105	208	106	209
rect	105	211	106	212
rect	105	214	106	215
rect	105	217	106	218
rect	105	220	106	221
rect	105	223	106	224
rect	105	226	106	227
rect	105	229	106	230
rect	105	232	106	233
rect	105	235	106	236
rect	105	238	106	239
rect	105	241	106	242
rect	105	244	106	245
rect	105	247	106	248
rect	105	250	106	251
rect	105	253	106	254
rect	105	256	106	257
rect	105	259	106	260
rect	105	262	106	263
rect	105	265	106	266
rect	105	268	106	269
rect	105	271	106	272
rect	105	274	106	275
rect	105	277	106	278
rect	105	280	106	281
rect	105	283	106	284
rect	105	286	106	287
rect	105	289	106	290
rect	105	292	106	293
rect	105	295	106	296
rect	105	298	106	299
rect	105	301	106	302
rect	105	304	106	305
rect	105	307	106	308
rect	105	310	106	311
rect	105	313	106	314
rect	105	316	106	317
rect	105	319	106	320
rect	105	322	106	323
rect	105	325	106	326
rect	105	328	106	329
rect	105	331	106	332
rect	105	334	106	335
rect	105	337	106	338
rect	105	340	106	341
rect	105	343	106	344
rect	105	346	106	347
rect	105	349	106	350
rect	105	352	106	353
rect	105	355	106	356
rect	105	358	106	359
rect	105	361	106	362
rect	105	364	106	365
rect	105	367	106	368
rect	105	373	106	374
rect	105	376	106	377
rect	105	379	106	380
rect	105	385	106	386
rect	106	1	107	2
rect	106	4	107	5
rect	106	7	107	8
rect	106	10	107	11
rect	106	13	107	14
rect	106	16	107	17
rect	106	19	107	20
rect	106	22	107	23
rect	106	25	107	26
rect	106	28	107	29
rect	106	31	107	32
rect	106	34	107	35
rect	106	37	107	38
rect	106	40	107	41
rect	106	43	107	44
rect	106	46	107	47
rect	106	49	107	50
rect	106	52	107	53
rect	106	55	107	56
rect	106	58	107	59
rect	106	61	107	62
rect	106	64	107	65
rect	106	67	107	68
rect	106	70	107	71
rect	106	73	107	74
rect	106	76	107	77
rect	106	79	107	80
rect	106	82	107	83
rect	106	85	107	86
rect	106	88	107	89
rect	106	91	107	92
rect	106	94	107	95
rect	106	97	107	98
rect	106	100	107	101
rect	106	103	107	104
rect	106	106	107	107
rect	106	109	107	110
rect	106	112	107	113
rect	106	115	107	116
rect	106	118	107	119
rect	106	121	107	122
rect	106	124	107	125
rect	106	127	107	128
rect	106	130	107	131
rect	106	133	107	134
rect	106	136	107	137
rect	106	139	107	140
rect	106	142	107	143
rect	106	145	107	146
rect	106	148	107	149
rect	106	151	107	152
rect	106	154	107	155
rect	106	157	107	158
rect	106	160	107	161
rect	106	163	107	164
rect	106	166	107	167
rect	106	169	107	170
rect	106	172	107	173
rect	106	175	107	176
rect	106	178	107	179
rect	106	181	107	182
rect	106	184	107	185
rect	106	187	107	188
rect	106	190	107	191
rect	106	193	107	194
rect	106	196	107	197
rect	106	199	107	200
rect	106	202	107	203
rect	106	205	107	206
rect	106	208	107	209
rect	106	211	107	212
rect	106	214	107	215
rect	106	217	107	218
rect	106	220	107	221
rect	106	223	107	224
rect	106	226	107	227
rect	106	229	107	230
rect	106	232	107	233
rect	106	235	107	236
rect	106	238	107	239
rect	106	241	107	242
rect	106	244	107	245
rect	106	247	107	248
rect	106	250	107	251
rect	106	253	107	254
rect	106	256	107	257
rect	106	259	107	260
rect	106	262	107	263
rect	106	265	107	266
rect	106	268	107	269
rect	106	271	107	272
rect	106	274	107	275
rect	106	277	107	278
rect	106	280	107	281
rect	106	283	107	284
rect	106	286	107	287
rect	106	289	107	290
rect	106	292	107	293
rect	106	295	107	296
rect	106	298	107	299
rect	106	301	107	302
rect	106	304	107	305
rect	106	307	107	308
rect	106	310	107	311
rect	106	313	107	314
rect	106	316	107	317
rect	106	319	107	320
rect	106	322	107	323
rect	106	325	107	326
rect	106	328	107	329
rect	106	331	107	332
rect	106	334	107	335
rect	106	337	107	338
rect	106	340	107	341
rect	106	343	107	344
rect	106	346	107	347
rect	106	349	107	350
rect	106	352	107	353
rect	106	355	107	356
rect	106	358	107	359
rect	106	361	107	362
rect	106	364	107	365
rect	106	367	107	368
rect	106	373	107	374
rect	106	376	107	377
rect	106	379	107	380
rect	106	385	107	386
rect	107	1	108	2
rect	107	4	108	5
rect	107	7	108	8
rect	107	10	108	11
rect	107	13	108	14
rect	107	16	108	17
rect	107	19	108	20
rect	107	22	108	23
rect	107	25	108	26
rect	107	28	108	29
rect	107	31	108	32
rect	107	34	108	35
rect	107	37	108	38
rect	107	40	108	41
rect	107	43	108	44
rect	107	46	108	47
rect	107	49	108	50
rect	107	52	108	53
rect	107	55	108	56
rect	107	58	108	59
rect	107	61	108	62
rect	107	64	108	65
rect	107	67	108	68
rect	107	70	108	71
rect	107	73	108	74
rect	107	76	108	77
rect	107	79	108	80
rect	107	82	108	83
rect	107	85	108	86
rect	107	88	108	89
rect	107	91	108	92
rect	107	94	108	95
rect	107	97	108	98
rect	107	100	108	101
rect	107	103	108	104
rect	107	106	108	107
rect	107	109	108	110
rect	107	112	108	113
rect	107	115	108	116
rect	107	118	108	119
rect	107	121	108	122
rect	107	124	108	125
rect	107	127	108	128
rect	107	130	108	131
rect	107	133	108	134
rect	107	136	108	137
rect	107	139	108	140
rect	107	142	108	143
rect	107	145	108	146
rect	107	148	108	149
rect	107	151	108	152
rect	107	154	108	155
rect	107	157	108	158
rect	107	160	108	161
rect	107	163	108	164
rect	107	166	108	167
rect	107	169	108	170
rect	107	172	108	173
rect	107	175	108	176
rect	107	178	108	179
rect	107	181	108	182
rect	107	184	108	185
rect	107	187	108	188
rect	107	190	108	191
rect	107	193	108	194
rect	107	196	108	197
rect	107	199	108	200
rect	107	202	108	203
rect	107	205	108	206
rect	107	208	108	209
rect	107	211	108	212
rect	107	214	108	215
rect	107	217	108	218
rect	107	220	108	221
rect	107	223	108	224
rect	107	226	108	227
rect	107	229	108	230
rect	107	232	108	233
rect	107	235	108	236
rect	107	238	108	239
rect	107	241	108	242
rect	107	244	108	245
rect	107	247	108	248
rect	107	250	108	251
rect	107	253	108	254
rect	107	256	108	257
rect	107	259	108	260
rect	107	262	108	263
rect	107	265	108	266
rect	107	268	108	269
rect	107	271	108	272
rect	107	274	108	275
rect	107	277	108	278
rect	107	280	108	281
rect	107	283	108	284
rect	107	286	108	287
rect	107	289	108	290
rect	107	292	108	293
rect	107	295	108	296
rect	107	298	108	299
rect	107	301	108	302
rect	107	304	108	305
rect	107	307	108	308
rect	107	310	108	311
rect	107	313	108	314
rect	107	316	108	317
rect	107	319	108	320
rect	107	322	108	323
rect	107	325	108	326
rect	107	328	108	329
rect	107	331	108	332
rect	107	334	108	335
rect	107	337	108	338
rect	107	340	108	341
rect	107	343	108	344
rect	107	346	108	347
rect	107	349	108	350
rect	107	352	108	353
rect	107	355	108	356
rect	107	358	108	359
rect	107	361	108	362
rect	107	364	108	365
rect	107	367	108	368
rect	107	373	108	374
rect	107	376	108	377
rect	107	379	108	380
rect	107	385	108	386
rect	108	1	109	2
rect	108	4	109	5
rect	108	7	109	8
rect	108	10	109	11
rect	108	13	109	14
rect	108	16	109	17
rect	108	19	109	20
rect	108	22	109	23
rect	108	25	109	26
rect	108	28	109	29
rect	108	31	109	32
rect	108	34	109	35
rect	108	37	109	38
rect	108	40	109	41
rect	108	43	109	44
rect	108	46	109	47
rect	108	49	109	50
rect	108	52	109	53
rect	108	55	109	56
rect	108	58	109	59
rect	108	61	109	62
rect	108	64	109	65
rect	108	67	109	68
rect	108	70	109	71
rect	108	73	109	74
rect	108	76	109	77
rect	108	79	109	80
rect	108	82	109	83
rect	108	85	109	86
rect	108	88	109	89
rect	108	91	109	92
rect	108	94	109	95
rect	108	97	109	98
rect	108	100	109	101
rect	108	103	109	104
rect	108	106	109	107
rect	108	109	109	110
rect	108	112	109	113
rect	108	115	109	116
rect	108	118	109	119
rect	108	121	109	122
rect	108	124	109	125
rect	108	127	109	128
rect	108	130	109	131
rect	108	133	109	134
rect	108	136	109	137
rect	108	139	109	140
rect	108	142	109	143
rect	108	145	109	146
rect	108	148	109	149
rect	108	151	109	152
rect	108	154	109	155
rect	108	157	109	158
rect	108	160	109	161
rect	108	163	109	164
rect	108	166	109	167
rect	108	169	109	170
rect	108	172	109	173
rect	108	175	109	176
rect	108	178	109	179
rect	108	181	109	182
rect	108	184	109	185
rect	108	187	109	188
rect	108	190	109	191
rect	108	193	109	194
rect	108	196	109	197
rect	108	199	109	200
rect	108	202	109	203
rect	108	205	109	206
rect	108	208	109	209
rect	108	211	109	212
rect	108	214	109	215
rect	108	217	109	218
rect	108	220	109	221
rect	108	223	109	224
rect	108	226	109	227
rect	108	229	109	230
rect	108	232	109	233
rect	108	235	109	236
rect	108	238	109	239
rect	108	241	109	242
rect	108	244	109	245
rect	108	247	109	248
rect	108	250	109	251
rect	108	253	109	254
rect	108	256	109	257
rect	108	259	109	260
rect	108	262	109	263
rect	108	265	109	266
rect	108	268	109	269
rect	108	271	109	272
rect	108	274	109	275
rect	108	277	109	278
rect	108	280	109	281
rect	108	283	109	284
rect	108	286	109	287
rect	108	289	109	290
rect	108	292	109	293
rect	108	295	109	296
rect	108	298	109	299
rect	108	301	109	302
rect	108	304	109	305
rect	108	307	109	308
rect	108	310	109	311
rect	108	313	109	314
rect	108	316	109	317
rect	108	319	109	320
rect	108	322	109	323
rect	108	325	109	326
rect	108	328	109	329
rect	108	331	109	332
rect	108	334	109	335
rect	108	337	109	338
rect	108	340	109	341
rect	108	343	109	344
rect	108	346	109	347
rect	108	349	109	350
rect	108	352	109	353
rect	108	355	109	356
rect	108	358	109	359
rect	108	361	109	362
rect	108	364	109	365
rect	108	367	109	368
rect	108	373	109	374
rect	108	376	109	377
rect	108	379	109	380
rect	108	385	109	386
rect	109	1	110	2
rect	109	4	110	5
rect	109	7	110	8
rect	109	10	110	11
rect	109	13	110	14
rect	109	16	110	17
rect	109	19	110	20
rect	109	22	110	23
rect	109	25	110	26
rect	109	28	110	29
rect	109	31	110	32
rect	109	34	110	35
rect	109	37	110	38
rect	109	40	110	41
rect	109	43	110	44
rect	109	46	110	47
rect	109	49	110	50
rect	109	52	110	53
rect	109	55	110	56
rect	109	58	110	59
rect	109	61	110	62
rect	109	64	110	65
rect	109	67	110	68
rect	109	70	110	71
rect	109	73	110	74
rect	109	76	110	77
rect	109	79	110	80
rect	109	82	110	83
rect	109	85	110	86
rect	109	88	110	89
rect	109	91	110	92
rect	109	94	110	95
rect	109	97	110	98
rect	109	100	110	101
rect	109	103	110	104
rect	109	106	110	107
rect	109	109	110	110
rect	109	112	110	113
rect	109	115	110	116
rect	109	118	110	119
rect	109	121	110	122
rect	109	124	110	125
rect	109	127	110	128
rect	109	130	110	131
rect	109	133	110	134
rect	109	136	110	137
rect	109	139	110	140
rect	109	142	110	143
rect	109	145	110	146
rect	109	148	110	149
rect	109	151	110	152
rect	109	154	110	155
rect	109	157	110	158
rect	109	160	110	161
rect	109	163	110	164
rect	109	166	110	167
rect	109	169	110	170
rect	109	172	110	173
rect	109	175	110	176
rect	109	178	110	179
rect	109	181	110	182
rect	109	184	110	185
rect	109	187	110	188
rect	109	190	110	191
rect	109	193	110	194
rect	109	196	110	197
rect	109	199	110	200
rect	109	202	110	203
rect	109	205	110	206
rect	109	208	110	209
rect	109	211	110	212
rect	109	214	110	215
rect	109	217	110	218
rect	109	220	110	221
rect	109	223	110	224
rect	109	226	110	227
rect	109	229	110	230
rect	109	232	110	233
rect	109	235	110	236
rect	109	238	110	239
rect	109	241	110	242
rect	109	244	110	245
rect	109	247	110	248
rect	109	250	110	251
rect	109	253	110	254
rect	109	256	110	257
rect	109	259	110	260
rect	109	262	110	263
rect	109	265	110	266
rect	109	268	110	269
rect	109	271	110	272
rect	109	274	110	275
rect	109	277	110	278
rect	109	280	110	281
rect	109	283	110	284
rect	109	286	110	287
rect	109	289	110	290
rect	109	292	110	293
rect	109	295	110	296
rect	109	298	110	299
rect	109	301	110	302
rect	109	304	110	305
rect	109	307	110	308
rect	109	310	110	311
rect	109	313	110	314
rect	109	316	110	317
rect	109	319	110	320
rect	109	322	110	323
rect	109	325	110	326
rect	109	328	110	329
rect	109	331	110	332
rect	109	334	110	335
rect	109	337	110	338
rect	109	340	110	341
rect	109	343	110	344
rect	109	346	110	347
rect	109	349	110	350
rect	109	352	110	353
rect	109	355	110	356
rect	109	358	110	359
rect	109	361	110	362
rect	109	364	110	365
rect	109	367	110	368
rect	109	373	110	374
rect	109	376	110	377
rect	109	379	110	380
rect	109	385	110	386
rect	110	1	111	2
rect	110	4	111	5
rect	110	7	111	8
rect	110	10	111	11
rect	110	13	111	14
rect	110	16	111	17
rect	110	19	111	20
rect	110	22	111	23
rect	110	25	111	26
rect	110	28	111	29
rect	110	31	111	32
rect	110	34	111	35
rect	110	37	111	38
rect	110	40	111	41
rect	110	43	111	44
rect	110	46	111	47
rect	110	49	111	50
rect	110	52	111	53
rect	110	55	111	56
rect	110	58	111	59
rect	110	61	111	62
rect	110	64	111	65
rect	110	67	111	68
rect	110	70	111	71
rect	110	73	111	74
rect	110	76	111	77
rect	110	79	111	80
rect	110	82	111	83
rect	110	85	111	86
rect	110	88	111	89
rect	110	91	111	92
rect	110	94	111	95
rect	110	97	111	98
rect	110	100	111	101
rect	110	103	111	104
rect	110	106	111	107
rect	110	109	111	110
rect	110	112	111	113
rect	110	115	111	116
rect	110	118	111	119
rect	110	121	111	122
rect	110	124	111	125
rect	110	127	111	128
rect	110	130	111	131
rect	110	133	111	134
rect	110	136	111	137
rect	110	139	111	140
rect	110	142	111	143
rect	110	145	111	146
rect	110	148	111	149
rect	110	151	111	152
rect	110	154	111	155
rect	110	157	111	158
rect	110	160	111	161
rect	110	163	111	164
rect	110	166	111	167
rect	110	169	111	170
rect	110	172	111	173
rect	110	175	111	176
rect	110	178	111	179
rect	110	181	111	182
rect	110	184	111	185
rect	110	187	111	188
rect	110	190	111	191
rect	110	193	111	194
rect	110	196	111	197
rect	110	199	111	200
rect	110	202	111	203
rect	110	205	111	206
rect	110	208	111	209
rect	110	211	111	212
rect	110	214	111	215
rect	110	217	111	218
rect	110	220	111	221
rect	110	223	111	224
rect	110	226	111	227
rect	110	229	111	230
rect	110	232	111	233
rect	110	235	111	236
rect	110	238	111	239
rect	110	241	111	242
rect	110	244	111	245
rect	110	247	111	248
rect	110	250	111	251
rect	110	253	111	254
rect	110	256	111	257
rect	110	259	111	260
rect	110	262	111	263
rect	110	265	111	266
rect	110	268	111	269
rect	110	271	111	272
rect	110	274	111	275
rect	110	277	111	278
rect	110	280	111	281
rect	110	283	111	284
rect	110	286	111	287
rect	110	289	111	290
rect	110	292	111	293
rect	110	295	111	296
rect	110	298	111	299
rect	110	301	111	302
rect	110	304	111	305
rect	110	307	111	308
rect	110	310	111	311
rect	110	313	111	314
rect	110	316	111	317
rect	110	319	111	320
rect	110	322	111	323
rect	110	325	111	326
rect	110	328	111	329
rect	110	331	111	332
rect	110	334	111	335
rect	110	337	111	338
rect	110	340	111	341
rect	110	343	111	344
rect	110	346	111	347
rect	110	349	111	350
rect	110	352	111	353
rect	110	355	111	356
rect	110	358	111	359
rect	110	361	111	362
rect	110	364	111	365
rect	110	367	111	368
rect	110	373	111	374
rect	110	376	111	377
rect	110	379	111	380
rect	110	385	111	386
rect	111	1	112	2
rect	111	4	112	5
rect	111	7	112	8
rect	111	10	112	11
rect	111	13	112	14
rect	111	16	112	17
rect	111	19	112	20
rect	111	22	112	23
rect	111	25	112	26
rect	111	28	112	29
rect	111	31	112	32
rect	111	34	112	35
rect	111	37	112	38
rect	111	40	112	41
rect	111	43	112	44
rect	111	46	112	47
rect	111	49	112	50
rect	111	52	112	53
rect	111	55	112	56
rect	111	58	112	59
rect	111	61	112	62
rect	111	64	112	65
rect	111	67	112	68
rect	111	70	112	71
rect	111	73	112	74
rect	111	76	112	77
rect	111	79	112	80
rect	111	82	112	83
rect	111	85	112	86
rect	111	88	112	89
rect	111	91	112	92
rect	111	94	112	95
rect	111	97	112	98
rect	111	100	112	101
rect	111	103	112	104
rect	111	106	112	107
rect	111	109	112	110
rect	111	112	112	113
rect	111	115	112	116
rect	111	118	112	119
rect	111	121	112	122
rect	111	124	112	125
rect	111	127	112	128
rect	111	130	112	131
rect	111	133	112	134
rect	111	136	112	137
rect	111	139	112	140
rect	111	142	112	143
rect	111	145	112	146
rect	111	148	112	149
rect	111	151	112	152
rect	111	154	112	155
rect	111	157	112	158
rect	111	160	112	161
rect	111	163	112	164
rect	111	166	112	167
rect	111	169	112	170
rect	111	172	112	173
rect	111	175	112	176
rect	111	178	112	179
rect	111	181	112	182
rect	111	184	112	185
rect	111	187	112	188
rect	111	190	112	191
rect	111	193	112	194
rect	111	196	112	197
rect	111	199	112	200
rect	111	202	112	203
rect	111	205	112	206
rect	111	208	112	209
rect	111	211	112	212
rect	111	214	112	215
rect	111	217	112	218
rect	111	220	112	221
rect	111	223	112	224
rect	111	226	112	227
rect	111	229	112	230
rect	111	232	112	233
rect	111	235	112	236
rect	111	238	112	239
rect	111	241	112	242
rect	111	244	112	245
rect	111	247	112	248
rect	111	250	112	251
rect	111	253	112	254
rect	111	256	112	257
rect	111	259	112	260
rect	111	262	112	263
rect	111	265	112	266
rect	111	268	112	269
rect	111	271	112	272
rect	111	274	112	275
rect	111	277	112	278
rect	111	280	112	281
rect	111	283	112	284
rect	111	286	112	287
rect	111	289	112	290
rect	111	292	112	293
rect	111	295	112	296
rect	111	298	112	299
rect	111	301	112	302
rect	111	304	112	305
rect	111	307	112	308
rect	111	310	112	311
rect	111	313	112	314
rect	111	316	112	317
rect	111	319	112	320
rect	111	322	112	323
rect	111	325	112	326
rect	111	328	112	329
rect	111	331	112	332
rect	111	334	112	335
rect	111	337	112	338
rect	111	340	112	341
rect	111	343	112	344
rect	111	346	112	347
rect	111	349	112	350
rect	111	352	112	353
rect	111	355	112	356
rect	111	358	112	359
rect	111	361	112	362
rect	111	364	112	365
rect	111	367	112	368
rect	111	373	112	374
rect	111	376	112	377
rect	111	379	112	380
rect	111	385	112	386
rect	112	1	113	2
rect	112	4	113	5
rect	112	7	113	8
rect	112	10	113	11
rect	112	13	113	14
rect	112	16	113	17
rect	112	19	113	20
rect	112	22	113	23
rect	112	25	113	26
rect	112	28	113	29
rect	112	31	113	32
rect	112	34	113	35
rect	112	37	113	38
rect	112	40	113	41
rect	112	43	113	44
rect	112	46	113	47
rect	112	49	113	50
rect	112	52	113	53
rect	112	55	113	56
rect	112	58	113	59
rect	112	61	113	62
rect	112	64	113	65
rect	112	67	113	68
rect	112	70	113	71
rect	112	73	113	74
rect	112	76	113	77
rect	112	79	113	80
rect	112	82	113	83
rect	112	85	113	86
rect	112	88	113	89
rect	112	91	113	92
rect	112	94	113	95
rect	112	97	113	98
rect	112	100	113	101
rect	112	103	113	104
rect	112	106	113	107
rect	112	109	113	110
rect	112	112	113	113
rect	112	115	113	116
rect	112	118	113	119
rect	112	121	113	122
rect	112	124	113	125
rect	112	127	113	128
rect	112	130	113	131
rect	112	133	113	134
rect	112	136	113	137
rect	112	139	113	140
rect	112	142	113	143
rect	112	145	113	146
rect	112	148	113	149
rect	112	151	113	152
rect	112	154	113	155
rect	112	157	113	158
rect	112	160	113	161
rect	112	163	113	164
rect	112	166	113	167
rect	112	169	113	170
rect	112	172	113	173
rect	112	175	113	176
rect	112	178	113	179
rect	112	181	113	182
rect	112	184	113	185
rect	112	187	113	188
rect	112	190	113	191
rect	112	193	113	194
rect	112	196	113	197
rect	112	199	113	200
rect	112	202	113	203
rect	112	205	113	206
rect	112	208	113	209
rect	112	211	113	212
rect	112	214	113	215
rect	112	217	113	218
rect	112	220	113	221
rect	112	223	113	224
rect	112	226	113	227
rect	112	229	113	230
rect	112	232	113	233
rect	112	235	113	236
rect	112	238	113	239
rect	112	241	113	242
rect	112	244	113	245
rect	112	247	113	248
rect	112	250	113	251
rect	112	253	113	254
rect	112	256	113	257
rect	112	259	113	260
rect	112	262	113	263
rect	112	265	113	266
rect	112	268	113	269
rect	112	271	113	272
rect	112	274	113	275
rect	112	277	113	278
rect	112	280	113	281
rect	112	283	113	284
rect	112	286	113	287
rect	112	289	113	290
rect	112	292	113	293
rect	112	295	113	296
rect	112	298	113	299
rect	112	301	113	302
rect	112	304	113	305
rect	112	307	113	308
rect	112	310	113	311
rect	112	313	113	314
rect	112	316	113	317
rect	112	319	113	320
rect	112	322	113	323
rect	112	325	113	326
rect	112	328	113	329
rect	112	331	113	332
rect	112	334	113	335
rect	112	337	113	338
rect	112	340	113	341
rect	112	343	113	344
rect	112	346	113	347
rect	112	349	113	350
rect	112	352	113	353
rect	112	355	113	356
rect	112	358	113	359
rect	112	361	113	362
rect	112	364	113	365
rect	112	367	113	368
rect	112	373	113	374
rect	112	376	113	377
rect	112	379	113	380
rect	112	385	113	386
rect	113	1	114	2
rect	113	4	114	5
rect	113	7	114	8
rect	113	10	114	11
rect	113	13	114	14
rect	113	16	114	17
rect	113	19	114	20
rect	113	22	114	23
rect	113	25	114	26
rect	113	28	114	29
rect	113	31	114	32
rect	113	34	114	35
rect	113	37	114	38
rect	113	40	114	41
rect	113	43	114	44
rect	113	46	114	47
rect	113	49	114	50
rect	113	52	114	53
rect	113	55	114	56
rect	113	58	114	59
rect	113	61	114	62
rect	113	64	114	65
rect	113	67	114	68
rect	113	70	114	71
rect	113	73	114	74
rect	113	76	114	77
rect	113	79	114	80
rect	113	82	114	83
rect	113	85	114	86
rect	113	88	114	89
rect	113	91	114	92
rect	113	94	114	95
rect	113	97	114	98
rect	113	100	114	101
rect	113	103	114	104
rect	113	106	114	107
rect	113	109	114	110
rect	113	112	114	113
rect	113	115	114	116
rect	113	118	114	119
rect	113	121	114	122
rect	113	124	114	125
rect	113	127	114	128
rect	113	130	114	131
rect	113	133	114	134
rect	113	136	114	137
rect	113	139	114	140
rect	113	142	114	143
rect	113	145	114	146
rect	113	148	114	149
rect	113	151	114	152
rect	113	154	114	155
rect	113	157	114	158
rect	113	160	114	161
rect	113	163	114	164
rect	113	166	114	167
rect	113	169	114	170
rect	113	172	114	173
rect	113	175	114	176
rect	113	178	114	179
rect	113	181	114	182
rect	113	184	114	185
rect	113	187	114	188
rect	113	190	114	191
rect	113	193	114	194
rect	113	196	114	197
rect	113	199	114	200
rect	113	202	114	203
rect	113	205	114	206
rect	113	208	114	209
rect	113	211	114	212
rect	113	214	114	215
rect	113	217	114	218
rect	113	220	114	221
rect	113	223	114	224
rect	113	226	114	227
rect	113	229	114	230
rect	113	232	114	233
rect	113	235	114	236
rect	113	238	114	239
rect	113	241	114	242
rect	113	244	114	245
rect	113	247	114	248
rect	113	250	114	251
rect	113	253	114	254
rect	113	256	114	257
rect	113	259	114	260
rect	113	262	114	263
rect	113	265	114	266
rect	113	268	114	269
rect	113	271	114	272
rect	113	274	114	275
rect	113	277	114	278
rect	113	280	114	281
rect	113	283	114	284
rect	113	286	114	287
rect	113	289	114	290
rect	113	292	114	293
rect	113	295	114	296
rect	113	298	114	299
rect	113	301	114	302
rect	113	304	114	305
rect	113	307	114	308
rect	113	310	114	311
rect	113	313	114	314
rect	113	316	114	317
rect	113	319	114	320
rect	113	322	114	323
rect	113	325	114	326
rect	113	328	114	329
rect	113	331	114	332
rect	113	334	114	335
rect	113	337	114	338
rect	113	340	114	341
rect	113	343	114	344
rect	113	346	114	347
rect	113	349	114	350
rect	113	352	114	353
rect	113	355	114	356
rect	113	358	114	359
rect	113	361	114	362
rect	113	364	114	365
rect	113	367	114	368
rect	113	373	114	374
rect	113	376	114	377
rect	113	379	114	380
rect	113	385	114	386
rect	114	1	115	2
rect	114	4	115	5
rect	114	7	115	8
rect	114	10	115	11
rect	114	13	115	14
rect	114	16	115	17
rect	114	19	115	20
rect	114	22	115	23
rect	114	25	115	26
rect	114	28	115	29
rect	114	31	115	32
rect	114	34	115	35
rect	114	37	115	38
rect	114	40	115	41
rect	114	43	115	44
rect	114	46	115	47
rect	114	49	115	50
rect	114	52	115	53
rect	114	55	115	56
rect	114	58	115	59
rect	114	61	115	62
rect	114	64	115	65
rect	114	67	115	68
rect	114	70	115	71
rect	114	73	115	74
rect	114	76	115	77
rect	114	79	115	80
rect	114	82	115	83
rect	114	85	115	86
rect	114	88	115	89
rect	114	91	115	92
rect	114	94	115	95
rect	114	97	115	98
rect	114	100	115	101
rect	114	103	115	104
rect	114	106	115	107
rect	114	109	115	110
rect	114	112	115	113
rect	114	115	115	116
rect	114	118	115	119
rect	114	121	115	122
rect	114	124	115	125
rect	114	127	115	128
rect	114	130	115	131
rect	114	133	115	134
rect	114	136	115	137
rect	114	139	115	140
rect	114	142	115	143
rect	114	145	115	146
rect	114	148	115	149
rect	114	151	115	152
rect	114	154	115	155
rect	114	157	115	158
rect	114	160	115	161
rect	114	163	115	164
rect	114	166	115	167
rect	114	169	115	170
rect	114	172	115	173
rect	114	175	115	176
rect	114	178	115	179
rect	114	181	115	182
rect	114	184	115	185
rect	114	187	115	188
rect	114	190	115	191
rect	114	193	115	194
rect	114	196	115	197
rect	114	199	115	200
rect	114	202	115	203
rect	114	205	115	206
rect	114	208	115	209
rect	114	211	115	212
rect	114	214	115	215
rect	114	217	115	218
rect	114	220	115	221
rect	114	223	115	224
rect	114	226	115	227
rect	114	229	115	230
rect	114	232	115	233
rect	114	235	115	236
rect	114	238	115	239
rect	114	241	115	242
rect	114	244	115	245
rect	114	247	115	248
rect	114	250	115	251
rect	114	253	115	254
rect	114	256	115	257
rect	114	259	115	260
rect	114	262	115	263
rect	114	265	115	266
rect	114	268	115	269
rect	114	271	115	272
rect	114	274	115	275
rect	114	277	115	278
rect	114	280	115	281
rect	114	283	115	284
rect	114	286	115	287
rect	114	289	115	290
rect	114	292	115	293
rect	114	295	115	296
rect	114	298	115	299
rect	114	301	115	302
rect	114	304	115	305
rect	114	307	115	308
rect	114	310	115	311
rect	114	313	115	314
rect	114	316	115	317
rect	114	319	115	320
rect	114	322	115	323
rect	114	325	115	326
rect	114	328	115	329
rect	114	331	115	332
rect	114	334	115	335
rect	114	337	115	338
rect	114	340	115	341
rect	114	343	115	344
rect	114	346	115	347
rect	114	349	115	350
rect	114	352	115	353
rect	114	355	115	356
rect	114	358	115	359
rect	114	361	115	362
rect	114	364	115	365
rect	114	367	115	368
rect	114	373	115	374
rect	114	376	115	377
rect	114	379	115	380
rect	114	385	115	386
rect	115	1	116	2
rect	115	4	116	5
rect	115	7	116	8
rect	115	10	116	11
rect	115	13	116	14
rect	115	16	116	17
rect	115	19	116	20
rect	115	22	116	23
rect	115	25	116	26
rect	115	28	116	29
rect	115	31	116	32
rect	115	34	116	35
rect	115	37	116	38
rect	115	40	116	41
rect	115	43	116	44
rect	115	46	116	47
rect	115	49	116	50
rect	115	52	116	53
rect	115	55	116	56
rect	115	58	116	59
rect	115	61	116	62
rect	115	64	116	65
rect	115	67	116	68
rect	115	70	116	71
rect	115	73	116	74
rect	115	76	116	77
rect	115	79	116	80
rect	115	82	116	83
rect	115	85	116	86
rect	115	88	116	89
rect	115	91	116	92
rect	115	94	116	95
rect	115	97	116	98
rect	115	100	116	101
rect	115	103	116	104
rect	115	106	116	107
rect	115	109	116	110
rect	115	112	116	113
rect	115	115	116	116
rect	115	118	116	119
rect	115	121	116	122
rect	115	124	116	125
rect	115	127	116	128
rect	115	130	116	131
rect	115	133	116	134
rect	115	136	116	137
rect	115	139	116	140
rect	115	142	116	143
rect	115	145	116	146
rect	115	148	116	149
rect	115	151	116	152
rect	115	154	116	155
rect	115	157	116	158
rect	115	160	116	161
rect	115	163	116	164
rect	115	166	116	167
rect	115	169	116	170
rect	115	172	116	173
rect	115	175	116	176
rect	115	178	116	179
rect	115	181	116	182
rect	115	184	116	185
rect	115	187	116	188
rect	115	190	116	191
rect	115	193	116	194
rect	115	196	116	197
rect	115	199	116	200
rect	115	202	116	203
rect	115	205	116	206
rect	115	208	116	209
rect	115	211	116	212
rect	115	214	116	215
rect	115	217	116	218
rect	115	220	116	221
rect	115	223	116	224
rect	115	226	116	227
rect	115	229	116	230
rect	115	232	116	233
rect	115	235	116	236
rect	115	238	116	239
rect	115	241	116	242
rect	115	244	116	245
rect	115	247	116	248
rect	115	250	116	251
rect	115	253	116	254
rect	115	256	116	257
rect	115	259	116	260
rect	115	262	116	263
rect	115	265	116	266
rect	115	268	116	269
rect	115	271	116	272
rect	115	274	116	275
rect	115	277	116	278
rect	115	280	116	281
rect	115	283	116	284
rect	115	286	116	287
rect	115	289	116	290
rect	115	292	116	293
rect	115	295	116	296
rect	115	298	116	299
rect	115	301	116	302
rect	115	304	116	305
rect	115	307	116	308
rect	115	310	116	311
rect	115	313	116	314
rect	115	316	116	317
rect	115	319	116	320
rect	115	322	116	323
rect	115	325	116	326
rect	115	328	116	329
rect	115	331	116	332
rect	115	334	116	335
rect	115	337	116	338
rect	115	340	116	341
rect	115	343	116	344
rect	115	346	116	347
rect	115	349	116	350
rect	115	352	116	353
rect	115	355	116	356
rect	115	358	116	359
rect	115	361	116	362
rect	115	364	116	365
rect	115	367	116	368
rect	115	373	116	374
rect	115	376	116	377
rect	115	379	116	380
rect	115	385	116	386
rect	116	1	117	2
rect	116	4	117	5
rect	116	7	117	8
rect	116	10	117	11
rect	116	13	117	14
rect	116	16	117	17
rect	116	19	117	20
rect	116	22	117	23
rect	116	25	117	26
rect	116	28	117	29
rect	116	31	117	32
rect	116	34	117	35
rect	116	37	117	38
rect	116	40	117	41
rect	116	43	117	44
rect	116	46	117	47
rect	116	49	117	50
rect	116	52	117	53
rect	116	55	117	56
rect	116	58	117	59
rect	116	61	117	62
rect	116	64	117	65
rect	116	67	117	68
rect	116	70	117	71
rect	116	73	117	74
rect	116	76	117	77
rect	116	79	117	80
rect	116	82	117	83
rect	116	85	117	86
rect	116	88	117	89
rect	116	91	117	92
rect	116	94	117	95
rect	116	97	117	98
rect	116	100	117	101
rect	116	103	117	104
rect	116	106	117	107
rect	116	109	117	110
rect	116	112	117	113
rect	116	115	117	116
rect	116	118	117	119
rect	116	121	117	122
rect	116	124	117	125
rect	116	127	117	128
rect	116	130	117	131
rect	116	133	117	134
rect	116	136	117	137
rect	116	139	117	140
rect	116	142	117	143
rect	116	145	117	146
rect	116	148	117	149
rect	116	151	117	152
rect	116	154	117	155
rect	116	157	117	158
rect	116	160	117	161
rect	116	163	117	164
rect	116	166	117	167
rect	116	169	117	170
rect	116	172	117	173
rect	116	175	117	176
rect	116	178	117	179
rect	116	181	117	182
rect	116	184	117	185
rect	116	187	117	188
rect	116	190	117	191
rect	116	193	117	194
rect	116	196	117	197
rect	116	199	117	200
rect	116	202	117	203
rect	116	205	117	206
rect	116	208	117	209
rect	116	211	117	212
rect	116	214	117	215
rect	116	217	117	218
rect	116	220	117	221
rect	116	223	117	224
rect	116	226	117	227
rect	116	229	117	230
rect	116	232	117	233
rect	116	235	117	236
rect	116	238	117	239
rect	116	241	117	242
rect	116	244	117	245
rect	116	247	117	248
rect	116	250	117	251
rect	116	253	117	254
rect	116	256	117	257
rect	116	259	117	260
rect	116	262	117	263
rect	116	265	117	266
rect	116	268	117	269
rect	116	271	117	272
rect	116	274	117	275
rect	116	277	117	278
rect	116	280	117	281
rect	116	283	117	284
rect	116	286	117	287
rect	116	289	117	290
rect	116	292	117	293
rect	116	295	117	296
rect	116	298	117	299
rect	116	301	117	302
rect	116	304	117	305
rect	116	307	117	308
rect	116	310	117	311
rect	116	313	117	314
rect	116	316	117	317
rect	116	319	117	320
rect	116	322	117	323
rect	116	325	117	326
rect	116	328	117	329
rect	116	331	117	332
rect	116	334	117	335
rect	116	337	117	338
rect	116	340	117	341
rect	116	343	117	344
rect	116	346	117	347
rect	116	349	117	350
rect	116	352	117	353
rect	116	355	117	356
rect	116	358	117	359
rect	116	361	117	362
rect	116	364	117	365
rect	116	367	117	368
rect	116	373	117	374
rect	116	376	117	377
rect	116	379	117	380
rect	116	385	117	386
rect	117	1	118	2
rect	117	4	118	5
rect	117	7	118	8
rect	117	10	118	11
rect	117	13	118	14
rect	117	16	118	17
rect	117	19	118	20
rect	117	22	118	23
rect	117	25	118	26
rect	117	28	118	29
rect	117	31	118	32
rect	117	34	118	35
rect	117	37	118	38
rect	117	40	118	41
rect	117	43	118	44
rect	117	46	118	47
rect	117	49	118	50
rect	117	52	118	53
rect	117	55	118	56
rect	117	58	118	59
rect	117	61	118	62
rect	117	64	118	65
rect	117	67	118	68
rect	117	70	118	71
rect	117	73	118	74
rect	117	76	118	77
rect	117	79	118	80
rect	117	82	118	83
rect	117	85	118	86
rect	117	88	118	89
rect	117	91	118	92
rect	117	94	118	95
rect	117	97	118	98
rect	117	100	118	101
rect	117	103	118	104
rect	117	106	118	107
rect	117	109	118	110
rect	117	112	118	113
rect	117	115	118	116
rect	117	118	118	119
rect	117	121	118	122
rect	117	124	118	125
rect	117	127	118	128
rect	117	130	118	131
rect	117	133	118	134
rect	117	136	118	137
rect	117	139	118	140
rect	117	142	118	143
rect	117	145	118	146
rect	117	148	118	149
rect	117	151	118	152
rect	117	154	118	155
rect	117	157	118	158
rect	117	160	118	161
rect	117	163	118	164
rect	117	166	118	167
rect	117	169	118	170
rect	117	172	118	173
rect	117	175	118	176
rect	117	178	118	179
rect	117	181	118	182
rect	117	184	118	185
rect	117	187	118	188
rect	117	190	118	191
rect	117	193	118	194
rect	117	196	118	197
rect	117	199	118	200
rect	117	202	118	203
rect	117	205	118	206
rect	117	208	118	209
rect	117	211	118	212
rect	117	214	118	215
rect	117	217	118	218
rect	117	220	118	221
rect	117	223	118	224
rect	117	226	118	227
rect	117	229	118	230
rect	117	232	118	233
rect	117	235	118	236
rect	117	238	118	239
rect	117	241	118	242
rect	117	244	118	245
rect	117	247	118	248
rect	117	250	118	251
rect	117	253	118	254
rect	117	256	118	257
rect	117	259	118	260
rect	117	262	118	263
rect	117	265	118	266
rect	117	268	118	269
rect	117	271	118	272
rect	117	274	118	275
rect	117	277	118	278
rect	117	280	118	281
rect	117	283	118	284
rect	117	286	118	287
rect	117	289	118	290
rect	117	292	118	293
rect	117	295	118	296
rect	117	298	118	299
rect	117	301	118	302
rect	117	304	118	305
rect	117	307	118	308
rect	117	310	118	311
rect	117	313	118	314
rect	117	316	118	317
rect	117	319	118	320
rect	117	322	118	323
rect	117	325	118	326
rect	117	328	118	329
rect	117	331	118	332
rect	117	334	118	335
rect	117	337	118	338
rect	117	340	118	341
rect	117	343	118	344
rect	117	346	118	347
rect	117	349	118	350
rect	117	352	118	353
rect	117	355	118	356
rect	117	358	118	359
rect	117	361	118	362
rect	117	364	118	365
rect	117	367	118	368
rect	117	373	118	374
rect	117	376	118	377
rect	117	379	118	380
rect	117	385	118	386
rect	118	1	119	2
rect	118	4	119	5
rect	118	7	119	8
rect	118	10	119	11
rect	118	13	119	14
rect	118	16	119	17
rect	118	19	119	20
rect	118	22	119	23
rect	118	25	119	26
rect	118	28	119	29
rect	118	31	119	32
rect	118	34	119	35
rect	118	37	119	38
rect	118	40	119	41
rect	118	43	119	44
rect	118	46	119	47
rect	118	49	119	50
rect	118	52	119	53
rect	118	55	119	56
rect	118	58	119	59
rect	118	61	119	62
rect	118	64	119	65
rect	118	67	119	68
rect	118	70	119	71
rect	118	73	119	74
rect	118	76	119	77
rect	118	79	119	80
rect	118	82	119	83
rect	118	85	119	86
rect	118	88	119	89
rect	118	91	119	92
rect	118	94	119	95
rect	118	97	119	98
rect	118	100	119	101
rect	118	103	119	104
rect	118	106	119	107
rect	118	109	119	110
rect	118	112	119	113
rect	118	115	119	116
rect	118	118	119	119
rect	118	121	119	122
rect	118	124	119	125
rect	118	127	119	128
rect	118	130	119	131
rect	118	133	119	134
rect	118	136	119	137
rect	118	139	119	140
rect	118	142	119	143
rect	118	145	119	146
rect	118	148	119	149
rect	118	151	119	152
rect	118	154	119	155
rect	118	157	119	158
rect	118	160	119	161
rect	118	163	119	164
rect	118	166	119	167
rect	118	169	119	170
rect	118	172	119	173
rect	118	175	119	176
rect	118	178	119	179
rect	118	181	119	182
rect	118	184	119	185
rect	118	187	119	188
rect	118	190	119	191
rect	118	193	119	194
rect	118	196	119	197
rect	118	199	119	200
rect	118	202	119	203
rect	118	205	119	206
rect	118	208	119	209
rect	118	211	119	212
rect	118	214	119	215
rect	118	217	119	218
rect	118	220	119	221
rect	118	223	119	224
rect	118	226	119	227
rect	118	229	119	230
rect	118	232	119	233
rect	118	235	119	236
rect	118	238	119	239
rect	118	241	119	242
rect	118	244	119	245
rect	118	247	119	248
rect	118	250	119	251
rect	118	253	119	254
rect	118	256	119	257
rect	118	259	119	260
rect	118	262	119	263
rect	118	265	119	266
rect	118	268	119	269
rect	118	271	119	272
rect	118	274	119	275
rect	118	277	119	278
rect	118	280	119	281
rect	118	283	119	284
rect	118	286	119	287
rect	118	289	119	290
rect	118	292	119	293
rect	118	295	119	296
rect	118	298	119	299
rect	118	301	119	302
rect	118	304	119	305
rect	118	307	119	308
rect	118	310	119	311
rect	118	313	119	314
rect	118	316	119	317
rect	118	319	119	320
rect	118	322	119	323
rect	118	325	119	326
rect	118	328	119	329
rect	118	331	119	332
rect	118	334	119	335
rect	118	337	119	338
rect	118	340	119	341
rect	118	343	119	344
rect	118	346	119	347
rect	118	349	119	350
rect	118	352	119	353
rect	118	355	119	356
rect	118	358	119	359
rect	118	361	119	362
rect	118	364	119	365
rect	118	367	119	368
rect	118	373	119	374
rect	118	376	119	377
rect	118	379	119	380
rect	118	385	119	386
rect	119	1	120	2
rect	119	4	120	5
rect	119	7	120	8
rect	119	10	120	11
rect	119	13	120	14
rect	119	16	120	17
rect	119	19	120	20
rect	119	22	120	23
rect	119	25	120	26
rect	119	28	120	29
rect	119	31	120	32
rect	119	34	120	35
rect	119	37	120	38
rect	119	40	120	41
rect	119	43	120	44
rect	119	46	120	47
rect	119	49	120	50
rect	119	52	120	53
rect	119	55	120	56
rect	119	58	120	59
rect	119	61	120	62
rect	119	64	120	65
rect	119	67	120	68
rect	119	70	120	71
rect	119	73	120	74
rect	119	76	120	77
rect	119	79	120	80
rect	119	82	120	83
rect	119	85	120	86
rect	119	88	120	89
rect	119	91	120	92
rect	119	94	120	95
rect	119	97	120	98
rect	119	100	120	101
rect	119	103	120	104
rect	119	106	120	107
rect	119	109	120	110
rect	119	112	120	113
rect	119	115	120	116
rect	119	118	120	119
rect	119	121	120	122
rect	119	124	120	125
rect	119	127	120	128
rect	119	130	120	131
rect	119	133	120	134
rect	119	136	120	137
rect	119	139	120	140
rect	119	142	120	143
rect	119	145	120	146
rect	119	148	120	149
rect	119	151	120	152
rect	119	154	120	155
rect	119	157	120	158
rect	119	160	120	161
rect	119	163	120	164
rect	119	166	120	167
rect	119	169	120	170
rect	119	172	120	173
rect	119	175	120	176
rect	119	178	120	179
rect	119	181	120	182
rect	119	184	120	185
rect	119	187	120	188
rect	119	190	120	191
rect	119	193	120	194
rect	119	196	120	197
rect	119	199	120	200
rect	119	202	120	203
rect	119	205	120	206
rect	119	208	120	209
rect	119	211	120	212
rect	119	214	120	215
rect	119	217	120	218
rect	119	220	120	221
rect	119	223	120	224
rect	119	226	120	227
rect	119	229	120	230
rect	119	232	120	233
rect	119	235	120	236
rect	119	238	120	239
rect	119	241	120	242
rect	119	244	120	245
rect	119	247	120	248
rect	119	250	120	251
rect	119	253	120	254
rect	119	256	120	257
rect	119	259	120	260
rect	119	262	120	263
rect	119	265	120	266
rect	119	268	120	269
rect	119	271	120	272
rect	119	274	120	275
rect	119	277	120	278
rect	119	280	120	281
rect	119	283	120	284
rect	119	286	120	287
rect	119	289	120	290
rect	119	292	120	293
rect	119	295	120	296
rect	119	298	120	299
rect	119	301	120	302
rect	119	304	120	305
rect	119	307	120	308
rect	119	310	120	311
rect	119	313	120	314
rect	119	316	120	317
rect	119	319	120	320
rect	119	322	120	323
rect	119	325	120	326
rect	119	328	120	329
rect	119	331	120	332
rect	119	334	120	335
rect	119	337	120	338
rect	119	340	120	341
rect	119	343	120	344
rect	119	346	120	347
rect	119	349	120	350
rect	119	352	120	353
rect	119	355	120	356
rect	119	358	120	359
rect	119	361	120	362
rect	119	364	120	365
rect	119	367	120	368
rect	119	373	120	374
rect	119	376	120	377
rect	119	379	120	380
rect	119	385	120	386
rect	120	1	121	2
rect	120	4	121	5
rect	120	7	121	8
rect	120	10	121	11
rect	120	13	121	14
rect	120	16	121	17
rect	120	19	121	20
rect	120	22	121	23
rect	120	25	121	26
rect	120	28	121	29
rect	120	31	121	32
rect	120	34	121	35
rect	120	37	121	38
rect	120	40	121	41
rect	120	43	121	44
rect	120	46	121	47
rect	120	49	121	50
rect	120	52	121	53
rect	120	55	121	56
rect	120	58	121	59
rect	120	61	121	62
rect	120	64	121	65
rect	120	67	121	68
rect	120	70	121	71
rect	120	73	121	74
rect	120	76	121	77
rect	120	79	121	80
rect	120	82	121	83
rect	120	85	121	86
rect	120	88	121	89
rect	120	91	121	92
rect	120	94	121	95
rect	120	97	121	98
rect	120	100	121	101
rect	120	103	121	104
rect	120	106	121	107
rect	120	109	121	110
rect	120	112	121	113
rect	120	115	121	116
rect	120	118	121	119
rect	120	121	121	122
rect	120	124	121	125
rect	120	127	121	128
rect	120	130	121	131
rect	120	133	121	134
rect	120	136	121	137
rect	120	139	121	140
rect	120	142	121	143
rect	120	145	121	146
rect	120	148	121	149
rect	120	151	121	152
rect	120	154	121	155
rect	120	157	121	158
rect	120	160	121	161
rect	120	163	121	164
rect	120	166	121	167
rect	120	169	121	170
rect	120	172	121	173
rect	120	175	121	176
rect	120	178	121	179
rect	120	181	121	182
rect	120	184	121	185
rect	120	187	121	188
rect	120	190	121	191
rect	120	193	121	194
rect	120	196	121	197
rect	120	199	121	200
rect	120	202	121	203
rect	120	205	121	206
rect	120	208	121	209
rect	120	211	121	212
rect	120	214	121	215
rect	120	217	121	218
rect	120	220	121	221
rect	120	223	121	224
rect	120	226	121	227
rect	120	229	121	230
rect	120	232	121	233
rect	120	235	121	236
rect	120	238	121	239
rect	120	241	121	242
rect	120	244	121	245
rect	120	247	121	248
rect	120	250	121	251
rect	120	253	121	254
rect	120	256	121	257
rect	120	259	121	260
rect	120	262	121	263
rect	120	265	121	266
rect	120	268	121	269
rect	120	271	121	272
rect	120	274	121	275
rect	120	277	121	278
rect	120	280	121	281
rect	120	283	121	284
rect	120	286	121	287
rect	120	289	121	290
rect	120	292	121	293
rect	120	295	121	296
rect	120	298	121	299
rect	120	301	121	302
rect	120	304	121	305
rect	120	307	121	308
rect	120	310	121	311
rect	120	313	121	314
rect	120	316	121	317
rect	120	319	121	320
rect	120	322	121	323
rect	120	325	121	326
rect	120	328	121	329
rect	120	331	121	332
rect	120	334	121	335
rect	120	337	121	338
rect	120	340	121	341
rect	120	343	121	344
rect	120	346	121	347
rect	120	349	121	350
rect	120	352	121	353
rect	120	355	121	356
rect	120	358	121	359
rect	120	361	121	362
rect	120	364	121	365
rect	120	367	121	368
rect	120	373	121	374
rect	120	376	121	377
rect	120	379	121	380
rect	120	385	121	386
rect	121	1	122	2
rect	121	4	122	5
rect	121	7	122	8
rect	121	10	122	11
rect	121	13	122	14
rect	121	16	122	17
rect	121	19	122	20
rect	121	22	122	23
rect	121	25	122	26
rect	121	28	122	29
rect	121	31	122	32
rect	121	34	122	35
rect	121	37	122	38
rect	121	40	122	41
rect	121	43	122	44
rect	121	46	122	47
rect	121	49	122	50
rect	121	52	122	53
rect	121	55	122	56
rect	121	58	122	59
rect	121	61	122	62
rect	121	64	122	65
rect	121	67	122	68
rect	121	70	122	71
rect	121	73	122	74
rect	121	76	122	77
rect	121	79	122	80
rect	121	82	122	83
rect	121	85	122	86
rect	121	88	122	89
rect	121	91	122	92
rect	121	94	122	95
rect	121	97	122	98
rect	121	100	122	101
rect	121	103	122	104
rect	121	106	122	107
rect	121	109	122	110
rect	121	112	122	113
rect	121	115	122	116
rect	121	118	122	119
rect	121	121	122	122
rect	121	124	122	125
rect	121	127	122	128
rect	121	130	122	131
rect	121	133	122	134
rect	121	136	122	137
rect	121	139	122	140
rect	121	142	122	143
rect	121	145	122	146
rect	121	148	122	149
rect	121	151	122	152
rect	121	154	122	155
rect	121	157	122	158
rect	121	160	122	161
rect	121	163	122	164
rect	121	166	122	167
rect	121	169	122	170
rect	121	172	122	173
rect	121	175	122	176
rect	121	178	122	179
rect	121	181	122	182
rect	121	184	122	185
rect	121	187	122	188
rect	121	190	122	191
rect	121	193	122	194
rect	121	196	122	197
rect	121	199	122	200
rect	121	202	122	203
rect	121	205	122	206
rect	121	208	122	209
rect	121	211	122	212
rect	121	214	122	215
rect	121	217	122	218
rect	121	220	122	221
rect	121	223	122	224
rect	121	226	122	227
rect	121	229	122	230
rect	121	232	122	233
rect	121	235	122	236
rect	121	238	122	239
rect	121	241	122	242
rect	121	244	122	245
rect	121	247	122	248
rect	121	250	122	251
rect	121	253	122	254
rect	121	256	122	257
rect	121	259	122	260
rect	121	262	122	263
rect	121	265	122	266
rect	121	268	122	269
rect	121	271	122	272
rect	121	274	122	275
rect	121	277	122	278
rect	121	280	122	281
rect	121	283	122	284
rect	121	286	122	287
rect	121	289	122	290
rect	121	292	122	293
rect	121	295	122	296
rect	121	298	122	299
rect	121	301	122	302
rect	121	304	122	305
rect	121	307	122	308
rect	121	310	122	311
rect	121	313	122	314
rect	121	316	122	317
rect	121	319	122	320
rect	121	322	122	323
rect	121	325	122	326
rect	121	328	122	329
rect	121	331	122	332
rect	121	334	122	335
rect	121	337	122	338
rect	121	340	122	341
rect	121	343	122	344
rect	121	346	122	347
rect	121	349	122	350
rect	121	352	122	353
rect	121	355	122	356
rect	121	358	122	359
rect	121	361	122	362
rect	121	364	122	365
rect	121	367	122	368
rect	121	373	122	374
rect	121	376	122	377
rect	121	379	122	380
rect	121	385	122	386
rect	122	1	123	2
rect	122	4	123	5
rect	122	7	123	8
rect	122	10	123	11
rect	122	13	123	14
rect	122	16	123	17
rect	122	19	123	20
rect	122	22	123	23
rect	122	25	123	26
rect	122	28	123	29
rect	122	31	123	32
rect	122	34	123	35
rect	122	37	123	38
rect	122	40	123	41
rect	122	43	123	44
rect	122	46	123	47
rect	122	49	123	50
rect	122	52	123	53
rect	122	55	123	56
rect	122	58	123	59
rect	122	61	123	62
rect	122	64	123	65
rect	122	67	123	68
rect	122	70	123	71
rect	122	73	123	74
rect	122	76	123	77
rect	122	79	123	80
rect	122	82	123	83
rect	122	85	123	86
rect	122	88	123	89
rect	122	91	123	92
rect	122	94	123	95
rect	122	97	123	98
rect	122	100	123	101
rect	122	103	123	104
rect	122	106	123	107
rect	122	109	123	110
rect	122	112	123	113
rect	122	115	123	116
rect	122	118	123	119
rect	122	121	123	122
rect	122	124	123	125
rect	122	127	123	128
rect	122	130	123	131
rect	122	133	123	134
rect	122	136	123	137
rect	122	139	123	140
rect	122	142	123	143
rect	122	145	123	146
rect	122	148	123	149
rect	122	151	123	152
rect	122	154	123	155
rect	122	157	123	158
rect	122	160	123	161
rect	122	163	123	164
rect	122	166	123	167
rect	122	169	123	170
rect	122	172	123	173
rect	122	175	123	176
rect	122	178	123	179
rect	122	181	123	182
rect	122	184	123	185
rect	122	187	123	188
rect	122	190	123	191
rect	122	193	123	194
rect	122	196	123	197
rect	122	199	123	200
rect	122	202	123	203
rect	122	205	123	206
rect	122	208	123	209
rect	122	211	123	212
rect	122	214	123	215
rect	122	217	123	218
rect	122	220	123	221
rect	122	223	123	224
rect	122	226	123	227
rect	122	229	123	230
rect	122	232	123	233
rect	122	235	123	236
rect	122	238	123	239
rect	122	241	123	242
rect	122	244	123	245
rect	122	247	123	248
rect	122	250	123	251
rect	122	253	123	254
rect	122	256	123	257
rect	122	259	123	260
rect	122	262	123	263
rect	122	265	123	266
rect	122	268	123	269
rect	122	271	123	272
rect	122	274	123	275
rect	122	277	123	278
rect	122	280	123	281
rect	122	283	123	284
rect	122	286	123	287
rect	122	289	123	290
rect	122	292	123	293
rect	122	295	123	296
rect	122	298	123	299
rect	122	301	123	302
rect	122	304	123	305
rect	122	307	123	308
rect	122	310	123	311
rect	122	313	123	314
rect	122	316	123	317
rect	122	319	123	320
rect	122	322	123	323
rect	122	325	123	326
rect	122	328	123	329
rect	122	331	123	332
rect	122	334	123	335
rect	122	337	123	338
rect	122	340	123	341
rect	122	343	123	344
rect	122	346	123	347
rect	122	349	123	350
rect	122	352	123	353
rect	122	355	123	356
rect	122	358	123	359
rect	122	361	123	362
rect	122	364	123	365
rect	122	367	123	368
rect	122	373	123	374
rect	122	376	123	377
rect	122	379	123	380
rect	122	385	123	386
rect	123	1	124	2
rect	123	4	124	5
rect	123	7	124	8
rect	123	10	124	11
rect	123	13	124	14
rect	123	16	124	17
rect	123	19	124	20
rect	123	22	124	23
rect	123	25	124	26
rect	123	28	124	29
rect	123	31	124	32
rect	123	34	124	35
rect	123	37	124	38
rect	123	40	124	41
rect	123	43	124	44
rect	123	46	124	47
rect	123	49	124	50
rect	123	52	124	53
rect	123	55	124	56
rect	123	58	124	59
rect	123	61	124	62
rect	123	64	124	65
rect	123	67	124	68
rect	123	70	124	71
rect	123	73	124	74
rect	123	76	124	77
rect	123	79	124	80
rect	123	82	124	83
rect	123	85	124	86
rect	123	88	124	89
rect	123	91	124	92
rect	123	94	124	95
rect	123	97	124	98
rect	123	100	124	101
rect	123	103	124	104
rect	123	106	124	107
rect	123	109	124	110
rect	123	112	124	113
rect	123	115	124	116
rect	123	118	124	119
rect	123	121	124	122
rect	123	124	124	125
rect	123	127	124	128
rect	123	130	124	131
rect	123	133	124	134
rect	123	136	124	137
rect	123	139	124	140
rect	123	142	124	143
rect	123	145	124	146
rect	123	148	124	149
rect	123	151	124	152
rect	123	154	124	155
rect	123	157	124	158
rect	123	160	124	161
rect	123	163	124	164
rect	123	166	124	167
rect	123	169	124	170
rect	123	172	124	173
rect	123	175	124	176
rect	123	178	124	179
rect	123	181	124	182
rect	123	184	124	185
rect	123	187	124	188
rect	123	190	124	191
rect	123	193	124	194
rect	123	196	124	197
rect	123	199	124	200
rect	123	202	124	203
rect	123	205	124	206
rect	123	208	124	209
rect	123	211	124	212
rect	123	214	124	215
rect	123	217	124	218
rect	123	220	124	221
rect	123	223	124	224
rect	123	226	124	227
rect	123	229	124	230
rect	123	232	124	233
rect	123	235	124	236
rect	123	238	124	239
rect	123	241	124	242
rect	123	244	124	245
rect	123	247	124	248
rect	123	250	124	251
rect	123	253	124	254
rect	123	256	124	257
rect	123	259	124	260
rect	123	262	124	263
rect	123	265	124	266
rect	123	268	124	269
rect	123	271	124	272
rect	123	274	124	275
rect	123	277	124	278
rect	123	280	124	281
rect	123	283	124	284
rect	123	286	124	287
rect	123	289	124	290
rect	123	292	124	293
rect	123	295	124	296
rect	123	298	124	299
rect	123	301	124	302
rect	123	304	124	305
rect	123	307	124	308
rect	123	310	124	311
rect	123	313	124	314
rect	123	316	124	317
rect	123	319	124	320
rect	123	322	124	323
rect	123	325	124	326
rect	123	328	124	329
rect	123	331	124	332
rect	123	334	124	335
rect	123	337	124	338
rect	123	340	124	341
rect	123	343	124	344
rect	123	346	124	347
rect	123	349	124	350
rect	123	352	124	353
rect	123	355	124	356
rect	123	358	124	359
rect	123	361	124	362
rect	123	364	124	365
rect	123	367	124	368
rect	123	373	124	374
rect	123	376	124	377
rect	123	379	124	380
rect	123	385	124	386
rect	124	1	125	2
rect	124	4	125	5
rect	124	7	125	8
rect	124	10	125	11
rect	124	13	125	14
rect	124	16	125	17
rect	124	19	125	20
rect	124	22	125	23
rect	124	25	125	26
rect	124	28	125	29
rect	124	31	125	32
rect	124	34	125	35
rect	124	37	125	38
rect	124	40	125	41
rect	124	43	125	44
rect	124	46	125	47
rect	124	49	125	50
rect	124	52	125	53
rect	124	55	125	56
rect	124	58	125	59
rect	124	61	125	62
rect	124	64	125	65
rect	124	67	125	68
rect	124	70	125	71
rect	124	73	125	74
rect	124	76	125	77
rect	124	79	125	80
rect	124	82	125	83
rect	124	85	125	86
rect	124	88	125	89
rect	124	91	125	92
rect	124	94	125	95
rect	124	97	125	98
rect	124	100	125	101
rect	124	103	125	104
rect	124	106	125	107
rect	124	109	125	110
rect	124	112	125	113
rect	124	115	125	116
rect	124	118	125	119
rect	124	121	125	122
rect	124	124	125	125
rect	124	127	125	128
rect	124	130	125	131
rect	124	133	125	134
rect	124	136	125	137
rect	124	139	125	140
rect	124	142	125	143
rect	124	145	125	146
rect	124	148	125	149
rect	124	151	125	152
rect	124	154	125	155
rect	124	157	125	158
rect	124	160	125	161
rect	124	163	125	164
rect	124	166	125	167
rect	124	169	125	170
rect	124	172	125	173
rect	124	175	125	176
rect	124	178	125	179
rect	124	181	125	182
rect	124	184	125	185
rect	124	187	125	188
rect	124	190	125	191
rect	124	193	125	194
rect	124	196	125	197
rect	124	199	125	200
rect	124	202	125	203
rect	124	205	125	206
rect	124	208	125	209
rect	124	211	125	212
rect	124	214	125	215
rect	124	217	125	218
rect	124	220	125	221
rect	124	223	125	224
rect	124	226	125	227
rect	124	229	125	230
rect	124	232	125	233
rect	124	235	125	236
rect	124	238	125	239
rect	124	241	125	242
rect	124	244	125	245
rect	124	247	125	248
rect	124	250	125	251
rect	124	253	125	254
rect	124	256	125	257
rect	124	259	125	260
rect	124	262	125	263
rect	124	265	125	266
rect	124	268	125	269
rect	124	271	125	272
rect	124	274	125	275
rect	124	277	125	278
rect	124	280	125	281
rect	124	283	125	284
rect	124	286	125	287
rect	124	289	125	290
rect	124	292	125	293
rect	124	295	125	296
rect	124	298	125	299
rect	124	301	125	302
rect	124	304	125	305
rect	124	307	125	308
rect	124	310	125	311
rect	124	313	125	314
rect	124	316	125	317
rect	124	319	125	320
rect	124	322	125	323
rect	124	325	125	326
rect	124	328	125	329
rect	124	331	125	332
rect	124	334	125	335
rect	124	337	125	338
rect	124	340	125	341
rect	124	343	125	344
rect	124	346	125	347
rect	124	349	125	350
rect	124	352	125	353
rect	124	355	125	356
rect	124	358	125	359
rect	124	361	125	362
rect	124	364	125	365
rect	124	367	125	368
rect	124	373	125	374
rect	124	376	125	377
rect	124	379	125	380
rect	124	385	125	386
rect	125	1	126	2
rect	125	4	126	5
rect	125	7	126	8
rect	125	10	126	11
rect	125	13	126	14
rect	125	16	126	17
rect	125	19	126	20
rect	125	22	126	23
rect	125	25	126	26
rect	125	28	126	29
rect	125	31	126	32
rect	125	34	126	35
rect	125	37	126	38
rect	125	40	126	41
rect	125	43	126	44
rect	125	46	126	47
rect	125	49	126	50
rect	125	52	126	53
rect	125	55	126	56
rect	125	58	126	59
rect	125	61	126	62
rect	125	64	126	65
rect	125	67	126	68
rect	125	70	126	71
rect	125	73	126	74
rect	125	76	126	77
rect	125	79	126	80
rect	125	82	126	83
rect	125	85	126	86
rect	125	88	126	89
rect	125	91	126	92
rect	125	94	126	95
rect	125	97	126	98
rect	125	100	126	101
rect	125	103	126	104
rect	125	106	126	107
rect	125	109	126	110
rect	125	112	126	113
rect	125	115	126	116
rect	125	118	126	119
rect	125	121	126	122
rect	125	124	126	125
rect	125	127	126	128
rect	125	130	126	131
rect	125	133	126	134
rect	125	136	126	137
rect	125	139	126	140
rect	125	142	126	143
rect	125	145	126	146
rect	125	148	126	149
rect	125	151	126	152
rect	125	154	126	155
rect	125	157	126	158
rect	125	160	126	161
rect	125	163	126	164
rect	125	166	126	167
rect	125	169	126	170
rect	125	172	126	173
rect	125	175	126	176
rect	125	178	126	179
rect	125	181	126	182
rect	125	184	126	185
rect	125	187	126	188
rect	125	190	126	191
rect	125	193	126	194
rect	125	196	126	197
rect	125	199	126	200
rect	125	202	126	203
rect	125	205	126	206
rect	125	208	126	209
rect	125	211	126	212
rect	125	214	126	215
rect	125	217	126	218
rect	125	220	126	221
rect	125	223	126	224
rect	125	226	126	227
rect	125	229	126	230
rect	125	232	126	233
rect	125	235	126	236
rect	125	238	126	239
rect	125	241	126	242
rect	125	244	126	245
rect	125	247	126	248
rect	125	250	126	251
rect	125	253	126	254
rect	125	256	126	257
rect	125	259	126	260
rect	125	262	126	263
rect	125	265	126	266
rect	125	268	126	269
rect	125	271	126	272
rect	125	274	126	275
rect	125	277	126	278
rect	125	280	126	281
rect	125	283	126	284
rect	125	286	126	287
rect	125	289	126	290
rect	125	292	126	293
rect	125	295	126	296
rect	125	298	126	299
rect	125	301	126	302
rect	125	304	126	305
rect	125	307	126	308
rect	125	310	126	311
rect	125	313	126	314
rect	125	316	126	317
rect	125	319	126	320
rect	125	322	126	323
rect	125	325	126	326
rect	125	328	126	329
rect	125	331	126	332
rect	125	334	126	335
rect	125	337	126	338
rect	125	340	126	341
rect	125	343	126	344
rect	125	346	126	347
rect	125	349	126	350
rect	125	352	126	353
rect	125	355	126	356
rect	125	358	126	359
rect	125	361	126	362
rect	125	364	126	365
rect	125	367	126	368
rect	125	373	126	374
rect	125	376	126	377
rect	125	379	126	380
rect	125	385	126	386
rect	126	1	127	2
rect	126	4	127	5
rect	126	7	127	8
rect	126	10	127	11
rect	126	13	127	14
rect	126	16	127	17
rect	126	19	127	20
rect	126	22	127	23
rect	126	25	127	26
rect	126	28	127	29
rect	126	31	127	32
rect	126	34	127	35
rect	126	37	127	38
rect	126	40	127	41
rect	126	43	127	44
rect	126	46	127	47
rect	126	49	127	50
rect	126	52	127	53
rect	126	55	127	56
rect	126	58	127	59
rect	126	61	127	62
rect	126	64	127	65
rect	126	67	127	68
rect	126	70	127	71
rect	126	73	127	74
rect	126	76	127	77
rect	126	79	127	80
rect	126	82	127	83
rect	126	85	127	86
rect	126	88	127	89
rect	126	91	127	92
rect	126	94	127	95
rect	126	97	127	98
rect	126	100	127	101
rect	126	103	127	104
rect	126	106	127	107
rect	126	109	127	110
rect	126	112	127	113
rect	126	115	127	116
rect	126	118	127	119
rect	126	121	127	122
rect	126	124	127	125
rect	126	127	127	128
rect	126	130	127	131
rect	126	133	127	134
rect	126	136	127	137
rect	126	139	127	140
rect	126	142	127	143
rect	126	145	127	146
rect	126	148	127	149
rect	126	151	127	152
rect	126	154	127	155
rect	126	157	127	158
rect	126	160	127	161
rect	126	163	127	164
rect	126	166	127	167
rect	126	169	127	170
rect	126	172	127	173
rect	126	175	127	176
rect	126	178	127	179
rect	126	181	127	182
rect	126	184	127	185
rect	126	187	127	188
rect	126	190	127	191
rect	126	193	127	194
rect	126	196	127	197
rect	126	199	127	200
rect	126	202	127	203
rect	126	205	127	206
rect	126	208	127	209
rect	126	211	127	212
rect	126	214	127	215
rect	126	217	127	218
rect	126	220	127	221
rect	126	223	127	224
rect	126	226	127	227
rect	126	229	127	230
rect	126	232	127	233
rect	126	235	127	236
rect	126	238	127	239
rect	126	241	127	242
rect	126	244	127	245
rect	126	247	127	248
rect	126	250	127	251
rect	126	253	127	254
rect	126	256	127	257
rect	126	259	127	260
rect	126	262	127	263
rect	126	265	127	266
rect	126	268	127	269
rect	126	271	127	272
rect	126	274	127	275
rect	126	277	127	278
rect	126	280	127	281
rect	126	283	127	284
rect	126	286	127	287
rect	126	289	127	290
rect	126	292	127	293
rect	126	295	127	296
rect	126	298	127	299
rect	126	301	127	302
rect	126	304	127	305
rect	126	307	127	308
rect	126	310	127	311
rect	126	313	127	314
rect	126	316	127	317
rect	126	319	127	320
rect	126	322	127	323
rect	126	325	127	326
rect	126	328	127	329
rect	126	331	127	332
rect	126	334	127	335
rect	126	337	127	338
rect	126	340	127	341
rect	126	343	127	344
rect	126	346	127	347
rect	126	349	127	350
rect	126	352	127	353
rect	126	355	127	356
rect	126	358	127	359
rect	126	361	127	362
rect	126	364	127	365
rect	126	367	127	368
rect	126	373	127	374
rect	126	376	127	377
rect	126	379	127	380
rect	126	385	127	386
rect	127	1	128	2
rect	127	4	128	5
rect	127	7	128	8
rect	127	10	128	11
rect	127	13	128	14
rect	127	16	128	17
rect	127	19	128	20
rect	127	22	128	23
rect	127	25	128	26
rect	127	28	128	29
rect	127	31	128	32
rect	127	34	128	35
rect	127	37	128	38
rect	127	40	128	41
rect	127	43	128	44
rect	127	46	128	47
rect	127	49	128	50
rect	127	52	128	53
rect	127	55	128	56
rect	127	58	128	59
rect	127	61	128	62
rect	127	64	128	65
rect	127	67	128	68
rect	127	70	128	71
rect	127	73	128	74
rect	127	76	128	77
rect	127	79	128	80
rect	127	82	128	83
rect	127	85	128	86
rect	127	88	128	89
rect	127	91	128	92
rect	127	94	128	95
rect	127	97	128	98
rect	127	100	128	101
rect	127	103	128	104
rect	127	106	128	107
rect	127	109	128	110
rect	127	112	128	113
rect	127	115	128	116
rect	127	118	128	119
rect	127	121	128	122
rect	127	124	128	125
rect	127	127	128	128
rect	127	130	128	131
rect	127	133	128	134
rect	127	136	128	137
rect	127	139	128	140
rect	127	142	128	143
rect	127	145	128	146
rect	127	148	128	149
rect	127	151	128	152
rect	127	154	128	155
rect	127	157	128	158
rect	127	160	128	161
rect	127	163	128	164
rect	127	166	128	167
rect	127	169	128	170
rect	127	172	128	173
rect	127	175	128	176
rect	127	178	128	179
rect	127	181	128	182
rect	127	184	128	185
rect	127	187	128	188
rect	127	190	128	191
rect	127	193	128	194
rect	127	196	128	197
rect	127	199	128	200
rect	127	202	128	203
rect	127	205	128	206
rect	127	208	128	209
rect	127	211	128	212
rect	127	214	128	215
rect	127	217	128	218
rect	127	220	128	221
rect	127	223	128	224
rect	127	226	128	227
rect	127	229	128	230
rect	127	232	128	233
rect	127	235	128	236
rect	127	238	128	239
rect	127	241	128	242
rect	127	244	128	245
rect	127	247	128	248
rect	127	250	128	251
rect	127	253	128	254
rect	127	256	128	257
rect	127	259	128	260
rect	127	262	128	263
rect	127	265	128	266
rect	127	268	128	269
rect	127	271	128	272
rect	127	274	128	275
rect	127	277	128	278
rect	127	280	128	281
rect	127	283	128	284
rect	127	286	128	287
rect	127	289	128	290
rect	127	292	128	293
rect	127	295	128	296
rect	127	298	128	299
rect	127	301	128	302
rect	127	304	128	305
rect	127	307	128	308
rect	127	310	128	311
rect	127	313	128	314
rect	127	316	128	317
rect	127	319	128	320
rect	127	322	128	323
rect	127	325	128	326
rect	127	328	128	329
rect	127	331	128	332
rect	127	334	128	335
rect	127	337	128	338
rect	127	340	128	341
rect	127	343	128	344
rect	127	346	128	347
rect	127	349	128	350
rect	127	352	128	353
rect	127	355	128	356
rect	127	358	128	359
rect	127	361	128	362
rect	127	364	128	365
rect	127	367	128	368
rect	127	373	128	374
rect	127	376	128	377
rect	127	379	128	380
rect	127	385	128	386
rect	128	1	129	2
rect	128	4	129	5
rect	128	7	129	8
rect	128	10	129	11
rect	128	13	129	14
rect	128	16	129	17
rect	128	19	129	20
rect	128	22	129	23
rect	128	25	129	26
rect	128	28	129	29
rect	128	31	129	32
rect	128	34	129	35
rect	128	37	129	38
rect	128	40	129	41
rect	128	43	129	44
rect	128	46	129	47
rect	128	49	129	50
rect	128	52	129	53
rect	128	55	129	56
rect	128	58	129	59
rect	128	61	129	62
rect	128	64	129	65
rect	128	67	129	68
rect	128	70	129	71
rect	128	73	129	74
rect	128	76	129	77
rect	128	79	129	80
rect	128	82	129	83
rect	128	85	129	86
rect	128	88	129	89
rect	128	91	129	92
rect	128	94	129	95
rect	128	97	129	98
rect	128	100	129	101
rect	128	103	129	104
rect	128	106	129	107
rect	128	109	129	110
rect	128	112	129	113
rect	128	115	129	116
rect	128	118	129	119
rect	128	121	129	122
rect	128	124	129	125
rect	128	127	129	128
rect	128	130	129	131
rect	128	133	129	134
rect	128	136	129	137
rect	128	139	129	140
rect	128	142	129	143
rect	128	145	129	146
rect	128	148	129	149
rect	128	151	129	152
rect	128	154	129	155
rect	128	157	129	158
rect	128	160	129	161
rect	128	163	129	164
rect	128	166	129	167
rect	128	169	129	170
rect	128	172	129	173
rect	128	175	129	176
rect	128	178	129	179
rect	128	181	129	182
rect	128	184	129	185
rect	128	187	129	188
rect	128	190	129	191
rect	128	193	129	194
rect	128	196	129	197
rect	128	199	129	200
rect	128	202	129	203
rect	128	205	129	206
rect	128	208	129	209
rect	128	211	129	212
rect	128	214	129	215
rect	128	217	129	218
rect	128	220	129	221
rect	128	223	129	224
rect	128	226	129	227
rect	128	229	129	230
rect	128	232	129	233
rect	128	235	129	236
rect	128	238	129	239
rect	128	241	129	242
rect	128	244	129	245
rect	128	247	129	248
rect	128	250	129	251
rect	128	253	129	254
rect	128	256	129	257
rect	128	259	129	260
rect	128	262	129	263
rect	128	265	129	266
rect	128	268	129	269
rect	128	271	129	272
rect	128	274	129	275
rect	128	277	129	278
rect	128	280	129	281
rect	128	283	129	284
rect	128	286	129	287
rect	128	289	129	290
rect	128	292	129	293
rect	128	295	129	296
rect	128	298	129	299
rect	128	301	129	302
rect	128	304	129	305
rect	128	307	129	308
rect	128	310	129	311
rect	128	313	129	314
rect	128	316	129	317
rect	128	319	129	320
rect	128	322	129	323
rect	128	325	129	326
rect	128	328	129	329
rect	128	331	129	332
rect	128	334	129	335
rect	128	337	129	338
rect	128	340	129	341
rect	128	343	129	344
rect	128	346	129	347
rect	128	349	129	350
rect	128	352	129	353
rect	128	355	129	356
rect	128	358	129	359
rect	128	361	129	362
rect	128	364	129	365
rect	128	367	129	368
rect	128	373	129	374
rect	128	376	129	377
rect	128	379	129	380
rect	128	385	129	386
rect	129	1	130	2
rect	129	4	130	5
rect	129	7	130	8
rect	129	10	130	11
rect	129	13	130	14
rect	129	16	130	17
rect	129	19	130	20
rect	129	22	130	23
rect	129	25	130	26
rect	129	28	130	29
rect	129	31	130	32
rect	129	34	130	35
rect	129	37	130	38
rect	129	40	130	41
rect	129	43	130	44
rect	129	46	130	47
rect	129	49	130	50
rect	129	52	130	53
rect	129	55	130	56
rect	129	58	130	59
rect	129	61	130	62
rect	129	64	130	65
rect	129	67	130	68
rect	129	70	130	71
rect	129	73	130	74
rect	129	76	130	77
rect	129	79	130	80
rect	129	82	130	83
rect	129	85	130	86
rect	129	88	130	89
rect	129	91	130	92
rect	129	94	130	95
rect	129	97	130	98
rect	129	100	130	101
rect	129	103	130	104
rect	129	106	130	107
rect	129	109	130	110
rect	129	112	130	113
rect	129	115	130	116
rect	129	118	130	119
rect	129	121	130	122
rect	129	124	130	125
rect	129	127	130	128
rect	129	130	130	131
rect	129	133	130	134
rect	129	136	130	137
rect	129	139	130	140
rect	129	142	130	143
rect	129	145	130	146
rect	129	148	130	149
rect	129	151	130	152
rect	129	154	130	155
rect	129	157	130	158
rect	129	160	130	161
rect	129	163	130	164
rect	129	166	130	167
rect	129	169	130	170
rect	129	172	130	173
rect	129	175	130	176
rect	129	178	130	179
rect	129	181	130	182
rect	129	184	130	185
rect	129	187	130	188
rect	129	190	130	191
rect	129	193	130	194
rect	129	196	130	197
rect	129	199	130	200
rect	129	202	130	203
rect	129	205	130	206
rect	129	208	130	209
rect	129	211	130	212
rect	129	214	130	215
rect	129	217	130	218
rect	129	220	130	221
rect	129	223	130	224
rect	129	226	130	227
rect	129	229	130	230
rect	129	232	130	233
rect	129	235	130	236
rect	129	238	130	239
rect	129	241	130	242
rect	129	244	130	245
rect	129	247	130	248
rect	129	250	130	251
rect	129	253	130	254
rect	129	256	130	257
rect	129	259	130	260
rect	129	262	130	263
rect	129	265	130	266
rect	129	268	130	269
rect	129	271	130	272
rect	129	274	130	275
rect	129	277	130	278
rect	129	280	130	281
rect	129	283	130	284
rect	129	286	130	287
rect	129	289	130	290
rect	129	292	130	293
rect	129	295	130	296
rect	129	298	130	299
rect	129	301	130	302
rect	129	304	130	305
rect	129	307	130	308
rect	129	310	130	311
rect	129	313	130	314
rect	129	316	130	317
rect	129	319	130	320
rect	129	322	130	323
rect	129	325	130	326
rect	129	328	130	329
rect	129	331	130	332
rect	129	334	130	335
rect	129	337	130	338
rect	129	340	130	341
rect	129	343	130	344
rect	129	346	130	347
rect	129	349	130	350
rect	129	352	130	353
rect	129	355	130	356
rect	129	358	130	359
rect	129	361	130	362
rect	129	364	130	365
rect	129	367	130	368
rect	129	373	130	374
rect	129	376	130	377
rect	129	379	130	380
rect	129	385	130	386
rect	130	1	131	2
rect	130	4	131	5
rect	130	7	131	8
rect	130	10	131	11
rect	130	13	131	14
rect	130	16	131	17
rect	130	19	131	20
rect	130	22	131	23
rect	130	25	131	26
rect	130	28	131	29
rect	130	31	131	32
rect	130	34	131	35
rect	130	37	131	38
rect	130	40	131	41
rect	130	43	131	44
rect	130	46	131	47
rect	130	49	131	50
rect	130	52	131	53
rect	130	55	131	56
rect	130	58	131	59
rect	130	61	131	62
rect	130	64	131	65
rect	130	67	131	68
rect	130	70	131	71
rect	130	73	131	74
rect	130	76	131	77
rect	130	79	131	80
rect	130	82	131	83
rect	130	85	131	86
rect	130	88	131	89
rect	130	91	131	92
rect	130	94	131	95
rect	130	97	131	98
rect	130	100	131	101
rect	130	103	131	104
rect	130	106	131	107
rect	130	109	131	110
rect	130	112	131	113
rect	130	115	131	116
rect	130	118	131	119
rect	130	121	131	122
rect	130	124	131	125
rect	130	127	131	128
rect	130	130	131	131
rect	130	133	131	134
rect	130	136	131	137
rect	130	139	131	140
rect	130	142	131	143
rect	130	145	131	146
rect	130	148	131	149
rect	130	151	131	152
rect	130	154	131	155
rect	130	157	131	158
rect	130	160	131	161
rect	130	163	131	164
rect	130	166	131	167
rect	130	169	131	170
rect	130	172	131	173
rect	130	175	131	176
rect	130	178	131	179
rect	130	181	131	182
rect	130	184	131	185
rect	130	187	131	188
rect	130	190	131	191
rect	130	193	131	194
rect	130	196	131	197
rect	130	199	131	200
rect	130	202	131	203
rect	130	205	131	206
rect	130	208	131	209
rect	130	211	131	212
rect	130	214	131	215
rect	130	217	131	218
rect	130	220	131	221
rect	130	223	131	224
rect	130	226	131	227
rect	130	229	131	230
rect	130	232	131	233
rect	130	235	131	236
rect	130	238	131	239
rect	130	241	131	242
rect	130	244	131	245
rect	130	247	131	248
rect	130	250	131	251
rect	130	253	131	254
rect	130	256	131	257
rect	130	259	131	260
rect	130	262	131	263
rect	130	265	131	266
rect	130	268	131	269
rect	130	271	131	272
rect	130	274	131	275
rect	130	277	131	278
rect	130	280	131	281
rect	130	283	131	284
rect	130	286	131	287
rect	130	289	131	290
rect	130	292	131	293
rect	130	295	131	296
rect	130	298	131	299
rect	130	301	131	302
rect	130	304	131	305
rect	130	307	131	308
rect	130	310	131	311
rect	130	313	131	314
rect	130	316	131	317
rect	130	319	131	320
rect	130	322	131	323
rect	130	325	131	326
rect	130	328	131	329
rect	130	331	131	332
rect	130	334	131	335
rect	130	340	131	341
rect	130	343	131	344
rect	130	346	131	347
rect	130	349	131	350
rect	130	352	131	353
rect	130	355	131	356
rect	130	358	131	359
rect	130	361	131	362
rect	130	364	131	365
rect	130	367	131	368
rect	130	373	131	374
rect	130	376	131	377
rect	130	379	131	380
rect	130	385	131	386
rect	131	1	132	2
rect	131	4	132	5
rect	131	7	132	8
rect	131	10	132	11
rect	131	13	132	14
rect	131	16	132	17
rect	131	19	132	20
rect	131	22	132	23
rect	131	25	132	26
rect	131	28	132	29
rect	131	31	132	32
rect	131	34	132	35
rect	131	37	132	38
rect	131	40	132	41
rect	131	43	132	44
rect	131	46	132	47
rect	131	49	132	50
rect	131	52	132	53
rect	131	55	132	56
rect	131	58	132	59
rect	131	61	132	62
rect	131	64	132	65
rect	131	67	132	68
rect	131	70	132	71
rect	131	73	132	74
rect	131	76	132	77
rect	131	79	132	80
rect	131	82	132	83
rect	131	85	132	86
rect	131	88	132	89
rect	131	91	132	92
rect	131	94	132	95
rect	131	97	132	98
rect	131	100	132	101
rect	131	103	132	104
rect	131	106	132	107
rect	131	109	132	110
rect	131	112	132	113
rect	131	115	132	116
rect	131	118	132	119
rect	131	121	132	122
rect	131	124	132	125
rect	131	127	132	128
rect	131	130	132	131
rect	131	133	132	134
rect	131	136	132	137
rect	131	139	132	140
rect	131	142	132	143
rect	131	145	132	146
rect	131	148	132	149
rect	131	151	132	152
rect	131	154	132	155
rect	131	157	132	158
rect	131	160	132	161
rect	131	163	132	164
rect	131	166	132	167
rect	131	169	132	170
rect	131	172	132	173
rect	131	175	132	176
rect	131	178	132	179
rect	131	181	132	182
rect	131	184	132	185
rect	131	187	132	188
rect	131	190	132	191
rect	131	193	132	194
rect	131	196	132	197
rect	131	199	132	200
rect	131	202	132	203
rect	131	205	132	206
rect	131	208	132	209
rect	131	211	132	212
rect	131	214	132	215
rect	131	217	132	218
rect	131	220	132	221
rect	131	223	132	224
rect	131	226	132	227
rect	131	229	132	230
rect	131	232	132	233
rect	131	235	132	236
rect	131	238	132	239
rect	131	241	132	242
rect	131	244	132	245
rect	131	247	132	248
rect	131	250	132	251
rect	131	253	132	254
rect	131	256	132	257
rect	131	259	132	260
rect	131	262	132	263
rect	131	265	132	266
rect	131	268	132	269
rect	131	271	132	272
rect	131	274	132	275
rect	131	277	132	278
rect	131	280	132	281
rect	131	283	132	284
rect	131	286	132	287
rect	131	289	132	290
rect	131	292	132	293
rect	131	295	132	296
rect	131	298	132	299
rect	131	301	132	302
rect	131	304	132	305
rect	131	307	132	308
rect	131	310	132	311
rect	131	313	132	314
rect	131	316	132	317
rect	131	319	132	320
rect	131	322	132	323
rect	131	325	132	326
rect	131	328	132	329
rect	131	331	132	332
rect	131	334	132	335
rect	131	340	132	341
rect	131	343	132	344
rect	131	346	132	347
rect	131	349	132	350
rect	131	352	132	353
rect	131	355	132	356
rect	131	358	132	359
rect	131	361	132	362
rect	131	364	132	365
rect	131	367	132	368
rect	131	373	132	374
rect	131	376	132	377
rect	131	379	132	380
rect	131	385	132	386
rect	132	1	133	2
rect	132	4	133	5
rect	132	7	133	8
rect	132	10	133	11
rect	132	13	133	14
rect	132	16	133	17
rect	132	19	133	20
rect	132	22	133	23
rect	132	25	133	26
rect	132	28	133	29
rect	132	31	133	32
rect	132	34	133	35
rect	132	37	133	38
rect	132	40	133	41
rect	132	43	133	44
rect	132	46	133	47
rect	132	49	133	50
rect	132	52	133	53
rect	132	55	133	56
rect	132	58	133	59
rect	132	61	133	62
rect	132	64	133	65
rect	132	67	133	68
rect	132	70	133	71
rect	132	73	133	74
rect	132	76	133	77
rect	132	79	133	80
rect	132	82	133	83
rect	132	85	133	86
rect	132	88	133	89
rect	132	91	133	92
rect	132	94	133	95
rect	132	97	133	98
rect	132	100	133	101
rect	132	103	133	104
rect	132	106	133	107
rect	132	109	133	110
rect	132	112	133	113
rect	132	115	133	116
rect	132	118	133	119
rect	132	121	133	122
rect	132	124	133	125
rect	132	127	133	128
rect	132	130	133	131
rect	132	133	133	134
rect	132	136	133	137
rect	132	139	133	140
rect	132	142	133	143
rect	132	145	133	146
rect	132	148	133	149
rect	132	151	133	152
rect	132	154	133	155
rect	132	157	133	158
rect	132	160	133	161
rect	132	163	133	164
rect	132	166	133	167
rect	132	169	133	170
rect	132	172	133	173
rect	132	175	133	176
rect	132	178	133	179
rect	132	181	133	182
rect	132	184	133	185
rect	132	187	133	188
rect	132	190	133	191
rect	132	193	133	194
rect	132	196	133	197
rect	132	199	133	200
rect	132	202	133	203
rect	132	205	133	206
rect	132	208	133	209
rect	132	211	133	212
rect	132	214	133	215
rect	132	217	133	218
rect	132	220	133	221
rect	132	223	133	224
rect	132	226	133	227
rect	132	229	133	230
rect	132	232	133	233
rect	132	235	133	236
rect	132	238	133	239
rect	132	241	133	242
rect	132	244	133	245
rect	132	247	133	248
rect	132	250	133	251
rect	132	253	133	254
rect	132	256	133	257
rect	132	259	133	260
rect	132	262	133	263
rect	132	265	133	266
rect	132	268	133	269
rect	132	271	133	272
rect	132	274	133	275
rect	132	277	133	278
rect	132	280	133	281
rect	132	283	133	284
rect	132	286	133	287
rect	132	289	133	290
rect	132	292	133	293
rect	132	295	133	296
rect	132	298	133	299
rect	132	301	133	302
rect	132	304	133	305
rect	132	307	133	308
rect	132	310	133	311
rect	132	313	133	314
rect	132	316	133	317
rect	132	319	133	320
rect	132	322	133	323
rect	132	325	133	326
rect	132	328	133	329
rect	132	331	133	332
rect	132	334	133	335
rect	132	340	133	341
rect	132	343	133	344
rect	132	346	133	347
rect	132	349	133	350
rect	132	352	133	353
rect	132	355	133	356
rect	132	358	133	359
rect	132	361	133	362
rect	132	364	133	365
rect	132	367	133	368
rect	132	373	133	374
rect	132	376	133	377
rect	132	379	133	380
rect	132	385	133	386
rect	133	1	134	2
rect	133	4	134	5
rect	133	7	134	8
rect	133	10	134	11
rect	133	13	134	14
rect	133	16	134	17
rect	133	19	134	20
rect	133	22	134	23
rect	133	25	134	26
rect	133	28	134	29
rect	133	31	134	32
rect	133	34	134	35
rect	133	37	134	38
rect	133	40	134	41
rect	133	43	134	44
rect	133	46	134	47
rect	133	49	134	50
rect	133	52	134	53
rect	133	55	134	56
rect	133	58	134	59
rect	133	61	134	62
rect	133	64	134	65
rect	133	67	134	68
rect	133	70	134	71
rect	133	73	134	74
rect	133	76	134	77
rect	133	79	134	80
rect	133	82	134	83
rect	133	85	134	86
rect	133	88	134	89
rect	133	91	134	92
rect	133	94	134	95
rect	133	97	134	98
rect	133	100	134	101
rect	133	103	134	104
rect	133	106	134	107
rect	133	109	134	110
rect	133	112	134	113
rect	133	115	134	116
rect	133	118	134	119
rect	133	121	134	122
rect	133	124	134	125
rect	133	127	134	128
rect	133	130	134	131
rect	133	133	134	134
rect	133	136	134	137
rect	133	139	134	140
rect	133	142	134	143
rect	133	145	134	146
rect	133	148	134	149
rect	133	151	134	152
rect	133	154	134	155
rect	133	157	134	158
rect	133	160	134	161
rect	133	163	134	164
rect	133	166	134	167
rect	133	169	134	170
rect	133	172	134	173
rect	133	175	134	176
rect	133	178	134	179
rect	133	181	134	182
rect	133	184	134	185
rect	133	187	134	188
rect	133	190	134	191
rect	133	193	134	194
rect	133	196	134	197
rect	133	199	134	200
rect	133	202	134	203
rect	133	205	134	206
rect	133	208	134	209
rect	133	211	134	212
rect	133	214	134	215
rect	133	217	134	218
rect	133	220	134	221
rect	133	223	134	224
rect	133	226	134	227
rect	133	229	134	230
rect	133	232	134	233
rect	133	235	134	236
rect	133	238	134	239
rect	133	241	134	242
rect	133	244	134	245
rect	133	247	134	248
rect	133	250	134	251
rect	133	253	134	254
rect	133	256	134	257
rect	133	259	134	260
rect	133	262	134	263
rect	133	265	134	266
rect	133	268	134	269
rect	133	271	134	272
rect	133	274	134	275
rect	133	277	134	278
rect	133	280	134	281
rect	133	283	134	284
rect	133	286	134	287
rect	133	289	134	290
rect	133	292	134	293
rect	133	295	134	296
rect	133	298	134	299
rect	133	301	134	302
rect	133	304	134	305
rect	133	307	134	308
rect	133	310	134	311
rect	133	313	134	314
rect	133	316	134	317
rect	133	319	134	320
rect	133	322	134	323
rect	133	325	134	326
rect	133	328	134	329
rect	133	331	134	332
rect	133	334	134	335
rect	133	340	134	341
rect	133	343	134	344
rect	133	346	134	347
rect	133	349	134	350
rect	133	352	134	353
rect	133	355	134	356
rect	133	358	134	359
rect	133	361	134	362
rect	133	364	134	365
rect	133	367	134	368
rect	133	373	134	374
rect	133	376	134	377
rect	133	379	134	380
rect	133	385	134	386
rect	134	1	135	2
rect	134	4	135	5
rect	134	7	135	8
rect	134	10	135	11
rect	134	13	135	14
rect	134	16	135	17
rect	134	19	135	20
rect	134	22	135	23
rect	134	25	135	26
rect	134	28	135	29
rect	134	31	135	32
rect	134	34	135	35
rect	134	37	135	38
rect	134	40	135	41
rect	134	43	135	44
rect	134	46	135	47
rect	134	49	135	50
rect	134	52	135	53
rect	134	55	135	56
rect	134	58	135	59
rect	134	61	135	62
rect	134	64	135	65
rect	134	67	135	68
rect	134	70	135	71
rect	134	73	135	74
rect	134	76	135	77
rect	134	79	135	80
rect	134	82	135	83
rect	134	85	135	86
rect	134	88	135	89
rect	134	91	135	92
rect	134	94	135	95
rect	134	97	135	98
rect	134	100	135	101
rect	134	103	135	104
rect	134	106	135	107
rect	134	109	135	110
rect	134	112	135	113
rect	134	115	135	116
rect	134	118	135	119
rect	134	121	135	122
rect	134	124	135	125
rect	134	127	135	128
rect	134	130	135	131
rect	134	133	135	134
rect	134	136	135	137
rect	134	139	135	140
rect	134	142	135	143
rect	134	145	135	146
rect	134	148	135	149
rect	134	151	135	152
rect	134	154	135	155
rect	134	157	135	158
rect	134	160	135	161
rect	134	163	135	164
rect	134	166	135	167
rect	134	169	135	170
rect	134	172	135	173
rect	134	175	135	176
rect	134	178	135	179
rect	134	181	135	182
rect	134	184	135	185
rect	134	187	135	188
rect	134	190	135	191
rect	134	193	135	194
rect	134	196	135	197
rect	134	199	135	200
rect	134	202	135	203
rect	134	205	135	206
rect	134	208	135	209
rect	134	211	135	212
rect	134	214	135	215
rect	134	217	135	218
rect	134	220	135	221
rect	134	223	135	224
rect	134	226	135	227
rect	134	229	135	230
rect	134	232	135	233
rect	134	235	135	236
rect	134	238	135	239
rect	134	241	135	242
rect	134	244	135	245
rect	134	247	135	248
rect	134	250	135	251
rect	134	253	135	254
rect	134	256	135	257
rect	134	259	135	260
rect	134	262	135	263
rect	134	265	135	266
rect	134	268	135	269
rect	134	271	135	272
rect	134	274	135	275
rect	134	277	135	278
rect	134	280	135	281
rect	134	283	135	284
rect	134	286	135	287
rect	134	289	135	290
rect	134	292	135	293
rect	134	295	135	296
rect	134	298	135	299
rect	134	301	135	302
rect	134	304	135	305
rect	134	307	135	308
rect	134	310	135	311
rect	134	313	135	314
rect	134	316	135	317
rect	134	319	135	320
rect	134	322	135	323
rect	134	325	135	326
rect	134	328	135	329
rect	134	331	135	332
rect	134	334	135	335
rect	134	340	135	341
rect	134	343	135	344
rect	134	346	135	347
rect	134	349	135	350
rect	134	352	135	353
rect	134	355	135	356
rect	134	358	135	359
rect	134	361	135	362
rect	134	364	135	365
rect	134	367	135	368
rect	134	373	135	374
rect	134	376	135	377
rect	134	379	135	380
rect	134	385	135	386
rect	135	1	136	2
rect	135	4	136	5
rect	135	7	136	8
rect	135	10	136	11
rect	135	13	136	14
rect	135	16	136	17
rect	135	19	136	20
rect	135	22	136	23
rect	135	25	136	26
rect	135	28	136	29
rect	135	31	136	32
rect	135	34	136	35
rect	135	37	136	38
rect	135	40	136	41
rect	135	43	136	44
rect	135	46	136	47
rect	135	49	136	50
rect	135	52	136	53
rect	135	55	136	56
rect	135	58	136	59
rect	135	61	136	62
rect	135	64	136	65
rect	135	67	136	68
rect	135	70	136	71
rect	135	73	136	74
rect	135	76	136	77
rect	135	79	136	80
rect	135	82	136	83
rect	135	85	136	86
rect	135	88	136	89
rect	135	91	136	92
rect	135	94	136	95
rect	135	97	136	98
rect	135	100	136	101
rect	135	103	136	104
rect	135	106	136	107
rect	135	109	136	110
rect	135	112	136	113
rect	135	115	136	116
rect	135	118	136	119
rect	135	121	136	122
rect	135	124	136	125
rect	135	127	136	128
rect	135	130	136	131
rect	135	133	136	134
rect	135	136	136	137
rect	135	139	136	140
rect	135	142	136	143
rect	135	145	136	146
rect	135	148	136	149
rect	135	151	136	152
rect	135	154	136	155
rect	135	157	136	158
rect	135	160	136	161
rect	135	163	136	164
rect	135	166	136	167
rect	135	169	136	170
rect	135	172	136	173
rect	135	175	136	176
rect	135	178	136	179
rect	135	181	136	182
rect	135	184	136	185
rect	135	187	136	188
rect	135	190	136	191
rect	135	193	136	194
rect	135	196	136	197
rect	135	199	136	200
rect	135	202	136	203
rect	135	205	136	206
rect	135	208	136	209
rect	135	211	136	212
rect	135	214	136	215
rect	135	217	136	218
rect	135	220	136	221
rect	135	223	136	224
rect	135	226	136	227
rect	135	229	136	230
rect	135	232	136	233
rect	135	235	136	236
rect	135	238	136	239
rect	135	241	136	242
rect	135	244	136	245
rect	135	247	136	248
rect	135	250	136	251
rect	135	253	136	254
rect	135	256	136	257
rect	135	259	136	260
rect	135	262	136	263
rect	135	265	136	266
rect	135	268	136	269
rect	135	271	136	272
rect	135	274	136	275
rect	135	277	136	278
rect	135	280	136	281
rect	135	283	136	284
rect	135	286	136	287
rect	135	289	136	290
rect	135	292	136	293
rect	135	295	136	296
rect	135	298	136	299
rect	135	301	136	302
rect	135	304	136	305
rect	135	307	136	308
rect	135	310	136	311
rect	135	313	136	314
rect	135	316	136	317
rect	135	319	136	320
rect	135	322	136	323
rect	135	325	136	326
rect	135	328	136	329
rect	135	331	136	332
rect	135	334	136	335
rect	135	340	136	341
rect	135	343	136	344
rect	135	346	136	347
rect	135	349	136	350
rect	135	352	136	353
rect	135	355	136	356
rect	135	358	136	359
rect	135	361	136	362
rect	135	364	136	365
rect	135	367	136	368
rect	135	373	136	374
rect	135	376	136	377
rect	135	379	136	380
rect	135	385	136	386
rect	136	1	137	2
rect	136	4	137	5
rect	136	7	137	8
rect	136	10	137	11
rect	136	13	137	14
rect	136	16	137	17
rect	136	19	137	20
rect	136	22	137	23
rect	136	25	137	26
rect	136	28	137	29
rect	136	31	137	32
rect	136	34	137	35
rect	136	37	137	38
rect	136	40	137	41
rect	136	43	137	44
rect	136	46	137	47
rect	136	49	137	50
rect	136	52	137	53
rect	136	55	137	56
rect	136	58	137	59
rect	136	61	137	62
rect	136	64	137	65
rect	136	67	137	68
rect	136	70	137	71
rect	136	73	137	74
rect	136	76	137	77
rect	136	79	137	80
rect	136	82	137	83
rect	136	85	137	86
rect	136	88	137	89
rect	136	91	137	92
rect	136	94	137	95
rect	136	97	137	98
rect	136	100	137	101
rect	136	103	137	104
rect	136	106	137	107
rect	136	109	137	110
rect	136	112	137	113
rect	136	115	137	116
rect	136	118	137	119
rect	136	121	137	122
rect	136	124	137	125
rect	136	127	137	128
rect	136	130	137	131
rect	136	133	137	134
rect	136	136	137	137
rect	136	139	137	140
rect	136	142	137	143
rect	136	145	137	146
rect	136	148	137	149
rect	136	151	137	152
rect	136	154	137	155
rect	136	157	137	158
rect	136	160	137	161
rect	136	163	137	164
rect	136	166	137	167
rect	136	169	137	170
rect	136	172	137	173
rect	136	175	137	176
rect	136	178	137	179
rect	136	181	137	182
rect	136	184	137	185
rect	136	187	137	188
rect	136	190	137	191
rect	136	193	137	194
rect	136	196	137	197
rect	136	199	137	200
rect	136	202	137	203
rect	136	205	137	206
rect	136	208	137	209
rect	136	211	137	212
rect	136	214	137	215
rect	136	217	137	218
rect	136	220	137	221
rect	136	223	137	224
rect	136	226	137	227
rect	136	229	137	230
rect	136	232	137	233
rect	136	235	137	236
rect	136	238	137	239
rect	136	241	137	242
rect	136	244	137	245
rect	136	247	137	248
rect	136	250	137	251
rect	136	253	137	254
rect	136	256	137	257
rect	136	259	137	260
rect	136	262	137	263
rect	136	265	137	266
rect	136	268	137	269
rect	136	271	137	272
rect	136	274	137	275
rect	136	277	137	278
rect	136	280	137	281
rect	136	283	137	284
rect	136	286	137	287
rect	136	289	137	290
rect	136	292	137	293
rect	136	295	137	296
rect	136	298	137	299
rect	136	301	137	302
rect	136	304	137	305
rect	136	307	137	308
rect	136	310	137	311
rect	136	313	137	314
rect	136	316	137	317
rect	136	319	137	320
rect	136	322	137	323
rect	136	325	137	326
rect	136	328	137	329
rect	136	331	137	332
rect	136	334	137	335
rect	136	340	137	341
rect	136	343	137	344
rect	136	346	137	347
rect	136	349	137	350
rect	136	352	137	353
rect	136	355	137	356
rect	136	358	137	359
rect	136	361	137	362
rect	136	364	137	365
rect	136	367	137	368
rect	136	373	137	374
rect	136	376	137	377
rect	136	379	137	380
rect	136	385	137	386
rect	137	1	138	2
rect	137	4	138	5
rect	137	7	138	8
rect	137	10	138	11
rect	137	13	138	14
rect	137	16	138	17
rect	137	19	138	20
rect	137	22	138	23
rect	137	25	138	26
rect	137	28	138	29
rect	137	31	138	32
rect	137	34	138	35
rect	137	37	138	38
rect	137	40	138	41
rect	137	43	138	44
rect	137	46	138	47
rect	137	49	138	50
rect	137	52	138	53
rect	137	55	138	56
rect	137	58	138	59
rect	137	61	138	62
rect	137	64	138	65
rect	137	67	138	68
rect	137	70	138	71
rect	137	73	138	74
rect	137	76	138	77
rect	137	79	138	80
rect	137	82	138	83
rect	137	85	138	86
rect	137	88	138	89
rect	137	91	138	92
rect	137	94	138	95
rect	137	97	138	98
rect	137	100	138	101
rect	137	103	138	104
rect	137	106	138	107
rect	137	109	138	110
rect	137	112	138	113
rect	137	115	138	116
rect	137	118	138	119
rect	137	121	138	122
rect	137	124	138	125
rect	137	127	138	128
rect	137	130	138	131
rect	137	133	138	134
rect	137	136	138	137
rect	137	139	138	140
rect	137	142	138	143
rect	137	145	138	146
rect	137	148	138	149
rect	137	151	138	152
rect	137	154	138	155
rect	137	157	138	158
rect	137	160	138	161
rect	137	163	138	164
rect	137	166	138	167
rect	137	169	138	170
rect	137	172	138	173
rect	137	175	138	176
rect	137	178	138	179
rect	137	181	138	182
rect	137	184	138	185
rect	137	187	138	188
rect	137	190	138	191
rect	137	193	138	194
rect	137	196	138	197
rect	137	199	138	200
rect	137	202	138	203
rect	137	205	138	206
rect	137	208	138	209
rect	137	211	138	212
rect	137	214	138	215
rect	137	217	138	218
rect	137	220	138	221
rect	137	223	138	224
rect	137	226	138	227
rect	137	229	138	230
rect	137	232	138	233
rect	137	235	138	236
rect	137	238	138	239
rect	137	241	138	242
rect	137	244	138	245
rect	137	247	138	248
rect	137	250	138	251
rect	137	253	138	254
rect	137	256	138	257
rect	137	259	138	260
rect	137	262	138	263
rect	137	265	138	266
rect	137	268	138	269
rect	137	271	138	272
rect	137	274	138	275
rect	137	277	138	278
rect	137	280	138	281
rect	137	283	138	284
rect	137	286	138	287
rect	137	289	138	290
rect	137	292	138	293
rect	137	295	138	296
rect	137	298	138	299
rect	137	301	138	302
rect	137	304	138	305
rect	137	307	138	308
rect	137	310	138	311
rect	137	313	138	314
rect	137	316	138	317
rect	137	319	138	320
rect	137	322	138	323
rect	137	325	138	326
rect	137	328	138	329
rect	137	331	138	332
rect	137	334	138	335
rect	137	340	138	341
rect	137	343	138	344
rect	137	346	138	347
rect	137	349	138	350
rect	137	352	138	353
rect	137	355	138	356
rect	137	358	138	359
rect	137	361	138	362
rect	137	364	138	365
rect	137	367	138	368
rect	137	373	138	374
rect	137	376	138	377
rect	137	379	138	380
rect	137	385	138	386
rect	138	1	139	2
rect	138	4	139	5
rect	138	7	139	8
rect	138	10	139	11
rect	138	13	139	14
rect	138	16	139	17
rect	138	19	139	20
rect	138	22	139	23
rect	138	25	139	26
rect	138	28	139	29
rect	138	31	139	32
rect	138	34	139	35
rect	138	37	139	38
rect	138	40	139	41
rect	138	43	139	44
rect	138	46	139	47
rect	138	49	139	50
rect	138	52	139	53
rect	138	55	139	56
rect	138	58	139	59
rect	138	61	139	62
rect	138	64	139	65
rect	138	67	139	68
rect	138	70	139	71
rect	138	73	139	74
rect	138	76	139	77
rect	138	79	139	80
rect	138	82	139	83
rect	138	85	139	86
rect	138	88	139	89
rect	138	91	139	92
rect	138	94	139	95
rect	138	97	139	98
rect	138	100	139	101
rect	138	103	139	104
rect	138	106	139	107
rect	138	109	139	110
rect	138	112	139	113
rect	138	115	139	116
rect	138	118	139	119
rect	138	121	139	122
rect	138	124	139	125
rect	138	127	139	128
rect	138	130	139	131
rect	138	133	139	134
rect	138	136	139	137
rect	138	139	139	140
rect	138	142	139	143
rect	138	145	139	146
rect	138	148	139	149
rect	138	151	139	152
rect	138	154	139	155
rect	138	157	139	158
rect	138	160	139	161
rect	138	163	139	164
rect	138	166	139	167
rect	138	169	139	170
rect	138	172	139	173
rect	138	175	139	176
rect	138	178	139	179
rect	138	181	139	182
rect	138	184	139	185
rect	138	187	139	188
rect	138	190	139	191
rect	138	193	139	194
rect	138	196	139	197
rect	138	199	139	200
rect	138	202	139	203
rect	138	205	139	206
rect	138	208	139	209
rect	138	211	139	212
rect	138	214	139	215
rect	138	217	139	218
rect	138	220	139	221
rect	138	223	139	224
rect	138	226	139	227
rect	138	229	139	230
rect	138	232	139	233
rect	138	235	139	236
rect	138	238	139	239
rect	138	241	139	242
rect	138	244	139	245
rect	138	247	139	248
rect	138	250	139	251
rect	138	253	139	254
rect	138	256	139	257
rect	138	259	139	260
rect	138	262	139	263
rect	138	265	139	266
rect	138	268	139	269
rect	138	271	139	272
rect	138	274	139	275
rect	138	277	139	278
rect	138	280	139	281
rect	138	283	139	284
rect	138	286	139	287
rect	138	289	139	290
rect	138	292	139	293
rect	138	295	139	296
rect	138	298	139	299
rect	138	301	139	302
rect	138	304	139	305
rect	138	307	139	308
rect	138	310	139	311
rect	138	313	139	314
rect	138	316	139	317
rect	138	319	139	320
rect	138	322	139	323
rect	138	325	139	326
rect	138	328	139	329
rect	138	331	139	332
rect	138	334	139	335
rect	138	340	139	341
rect	138	343	139	344
rect	138	346	139	347
rect	138	349	139	350
rect	138	352	139	353
rect	138	355	139	356
rect	138	358	139	359
rect	138	361	139	362
rect	138	364	139	365
rect	138	367	139	368
rect	138	373	139	374
rect	138	376	139	377
rect	138	379	139	380
rect	138	385	139	386
rect	139	1	140	2
rect	139	4	140	5
rect	139	7	140	8
rect	139	10	140	11
rect	139	13	140	14
rect	139	16	140	17
rect	139	19	140	20
rect	139	22	140	23
rect	139	25	140	26
rect	139	28	140	29
rect	139	31	140	32
rect	139	34	140	35
rect	139	37	140	38
rect	139	40	140	41
rect	139	43	140	44
rect	139	46	140	47
rect	139	49	140	50
rect	139	52	140	53
rect	139	55	140	56
rect	139	58	140	59
rect	139	61	140	62
rect	139	64	140	65
rect	139	67	140	68
rect	139	70	140	71
rect	139	73	140	74
rect	139	76	140	77
rect	139	79	140	80
rect	139	82	140	83
rect	139	85	140	86
rect	139	88	140	89
rect	139	91	140	92
rect	139	94	140	95
rect	139	97	140	98
rect	139	100	140	101
rect	139	103	140	104
rect	139	106	140	107
rect	139	109	140	110
rect	139	112	140	113
rect	139	115	140	116
rect	139	118	140	119
rect	139	121	140	122
rect	139	124	140	125
rect	139	127	140	128
rect	139	130	140	131
rect	139	133	140	134
rect	139	136	140	137
rect	139	139	140	140
rect	139	142	140	143
rect	139	145	140	146
rect	139	148	140	149
rect	139	151	140	152
rect	139	154	140	155
rect	139	157	140	158
rect	139	160	140	161
rect	139	163	140	164
rect	139	166	140	167
rect	139	169	140	170
rect	139	172	140	173
rect	139	175	140	176
rect	139	178	140	179
rect	139	181	140	182
rect	139	184	140	185
rect	139	187	140	188
rect	139	190	140	191
rect	139	193	140	194
rect	139	196	140	197
rect	139	199	140	200
rect	139	202	140	203
rect	139	205	140	206
rect	139	208	140	209
rect	139	211	140	212
rect	139	214	140	215
rect	139	217	140	218
rect	139	220	140	221
rect	139	223	140	224
rect	139	226	140	227
rect	139	229	140	230
rect	139	232	140	233
rect	139	235	140	236
rect	139	238	140	239
rect	139	241	140	242
rect	139	244	140	245
rect	139	247	140	248
rect	139	250	140	251
rect	139	253	140	254
rect	139	256	140	257
rect	139	259	140	260
rect	139	262	140	263
rect	139	265	140	266
rect	139	268	140	269
rect	139	271	140	272
rect	139	274	140	275
rect	139	277	140	278
rect	139	280	140	281
rect	139	283	140	284
rect	139	289	140	290
rect	139	292	140	293
rect	139	295	140	296
rect	139	298	140	299
rect	139	301	140	302
rect	139	304	140	305
rect	139	307	140	308
rect	139	310	140	311
rect	139	313	140	314
rect	139	316	140	317
rect	139	319	140	320
rect	139	322	140	323
rect	139	325	140	326
rect	139	328	140	329
rect	139	331	140	332
rect	139	334	140	335
rect	139	340	140	341
rect	139	343	140	344
rect	139	346	140	347
rect	139	349	140	350
rect	139	352	140	353
rect	139	355	140	356
rect	139	358	140	359
rect	139	361	140	362
rect	139	364	140	365
rect	139	367	140	368
rect	139	373	140	374
rect	139	376	140	377
rect	139	379	140	380
rect	139	385	140	386
rect	140	1	141	2
rect	140	4	141	5
rect	140	7	141	8
rect	140	10	141	11
rect	140	13	141	14
rect	140	16	141	17
rect	140	19	141	20
rect	140	22	141	23
rect	140	25	141	26
rect	140	28	141	29
rect	140	31	141	32
rect	140	34	141	35
rect	140	37	141	38
rect	140	40	141	41
rect	140	43	141	44
rect	140	46	141	47
rect	140	49	141	50
rect	140	52	141	53
rect	140	55	141	56
rect	140	58	141	59
rect	140	61	141	62
rect	140	64	141	65
rect	140	67	141	68
rect	140	70	141	71
rect	140	73	141	74
rect	140	76	141	77
rect	140	79	141	80
rect	140	82	141	83
rect	140	85	141	86
rect	140	88	141	89
rect	140	91	141	92
rect	140	94	141	95
rect	140	97	141	98
rect	140	100	141	101
rect	140	103	141	104
rect	140	106	141	107
rect	140	109	141	110
rect	140	112	141	113
rect	140	115	141	116
rect	140	118	141	119
rect	140	121	141	122
rect	140	124	141	125
rect	140	127	141	128
rect	140	130	141	131
rect	140	133	141	134
rect	140	136	141	137
rect	140	139	141	140
rect	140	142	141	143
rect	140	145	141	146
rect	140	148	141	149
rect	140	151	141	152
rect	140	154	141	155
rect	140	157	141	158
rect	140	160	141	161
rect	140	163	141	164
rect	140	166	141	167
rect	140	169	141	170
rect	140	172	141	173
rect	140	175	141	176
rect	140	178	141	179
rect	140	181	141	182
rect	140	184	141	185
rect	140	187	141	188
rect	140	190	141	191
rect	140	193	141	194
rect	140	196	141	197
rect	140	199	141	200
rect	140	202	141	203
rect	140	205	141	206
rect	140	208	141	209
rect	140	211	141	212
rect	140	214	141	215
rect	140	217	141	218
rect	140	220	141	221
rect	140	223	141	224
rect	140	226	141	227
rect	140	229	141	230
rect	140	232	141	233
rect	140	235	141	236
rect	140	238	141	239
rect	140	241	141	242
rect	140	244	141	245
rect	140	247	141	248
rect	140	250	141	251
rect	140	253	141	254
rect	140	256	141	257
rect	140	259	141	260
rect	140	262	141	263
rect	140	265	141	266
rect	140	268	141	269
rect	140	271	141	272
rect	140	274	141	275
rect	140	277	141	278
rect	140	280	141	281
rect	140	283	141	284
rect	140	286	141	287
rect	140	289	141	290
rect	140	292	141	293
rect	140	295	141	296
rect	140	298	141	299
rect	140	301	141	302
rect	140	304	141	305
rect	140	307	141	308
rect	140	310	141	311
rect	140	313	141	314
rect	140	316	141	317
rect	140	319	141	320
rect	140	322	141	323
rect	140	325	141	326
rect	140	328	141	329
rect	140	331	141	332
rect	140	334	141	335
rect	140	340	141	341
rect	140	343	141	344
rect	140	346	141	347
rect	140	349	141	350
rect	140	352	141	353
rect	140	355	141	356
rect	140	358	141	359
rect	140	361	141	362
rect	140	364	141	365
rect	140	367	141	368
rect	140	373	141	374
rect	140	376	141	377
rect	140	379	141	380
rect	140	385	141	386
rect	141	1	142	2
rect	141	4	142	5
rect	141	7	142	8
rect	141	10	142	11
rect	141	13	142	14
rect	141	16	142	17
rect	141	19	142	20
rect	141	22	142	23
rect	141	25	142	26
rect	141	28	142	29
rect	141	31	142	32
rect	141	34	142	35
rect	141	37	142	38
rect	141	40	142	41
rect	141	43	142	44
rect	141	46	142	47
rect	141	52	142	53
rect	141	55	142	56
rect	141	58	142	59
rect	141	61	142	62
rect	141	64	142	65
rect	141	67	142	68
rect	141	70	142	71
rect	141	73	142	74
rect	141	76	142	77
rect	141	79	142	80
rect	141	82	142	83
rect	141	85	142	86
rect	141	88	142	89
rect	141	91	142	92
rect	141	94	142	95
rect	141	97	142	98
rect	141	100	142	101
rect	141	103	142	104
rect	141	106	142	107
rect	141	109	142	110
rect	141	112	142	113
rect	141	115	142	116
rect	141	118	142	119
rect	141	121	142	122
rect	141	124	142	125
rect	141	127	142	128
rect	141	130	142	131
rect	141	133	142	134
rect	141	136	142	137
rect	141	139	142	140
rect	141	142	142	143
rect	141	145	142	146
rect	141	148	142	149
rect	141	151	142	152
rect	141	154	142	155
rect	141	157	142	158
rect	141	160	142	161
rect	141	163	142	164
rect	141	166	142	167
rect	141	169	142	170
rect	141	172	142	173
rect	141	175	142	176
rect	141	178	142	179
rect	141	181	142	182
rect	141	184	142	185
rect	141	187	142	188
rect	141	190	142	191
rect	141	193	142	194
rect	141	196	142	197
rect	141	199	142	200
rect	141	202	142	203
rect	141	205	142	206
rect	141	208	142	209
rect	141	211	142	212
rect	141	214	142	215
rect	141	217	142	218
rect	141	220	142	221
rect	141	223	142	224
rect	141	226	142	227
rect	141	229	142	230
rect	141	232	142	233
rect	141	235	142	236
rect	141	238	142	239
rect	141	241	142	242
rect	141	244	142	245
rect	141	247	142	248
rect	141	250	142	251
rect	141	253	142	254
rect	141	256	142	257
rect	141	259	142	260
rect	141	262	142	263
rect	141	265	142	266
rect	141	268	142	269
rect	141	271	142	272
rect	141	274	142	275
rect	141	277	142	278
rect	141	280	142	281
rect	141	283	142	284
rect	141	286	142	287
rect	141	289	142	290
rect	141	292	142	293
rect	141	298	142	299
rect	141	301	142	302
rect	141	304	142	305
rect	141	307	142	308
rect	141	310	142	311
rect	141	313	142	314
rect	141	316	142	317
rect	141	319	142	320
rect	141	322	142	323
rect	141	325	142	326
rect	141	328	142	329
rect	141	331	142	332
rect	141	334	142	335
rect	141	340	142	341
rect	141	343	142	344
rect	141	346	142	347
rect	141	349	142	350
rect	141	352	142	353
rect	141	355	142	356
rect	141	358	142	359
rect	141	361	142	362
rect	141	364	142	365
rect	141	367	142	368
rect	141	373	142	374
rect	141	376	142	377
rect	141	379	142	380
rect	141	385	142	386
rect	142	1	143	2
rect	142	4	143	5
rect	142	7	143	8
rect	142	10	143	11
rect	142	13	143	14
rect	142	16	143	17
rect	142	19	143	20
rect	142	22	143	23
rect	142	25	143	26
rect	142	28	143	29
rect	142	31	143	32
rect	142	34	143	35
rect	142	37	143	38
rect	142	40	143	41
rect	142	43	143	44
rect	142	46	143	47
rect	142	49	143	50
rect	142	52	143	53
rect	142	55	143	56
rect	142	58	143	59
rect	142	61	143	62
rect	142	64	143	65
rect	142	67	143	68
rect	142	70	143	71
rect	142	73	143	74
rect	142	76	143	77
rect	142	79	143	80
rect	142	82	143	83
rect	142	85	143	86
rect	142	88	143	89
rect	142	91	143	92
rect	142	94	143	95
rect	142	97	143	98
rect	142	100	143	101
rect	142	103	143	104
rect	142	106	143	107
rect	142	109	143	110
rect	142	112	143	113
rect	142	115	143	116
rect	142	118	143	119
rect	142	121	143	122
rect	142	124	143	125
rect	142	127	143	128
rect	142	130	143	131
rect	142	133	143	134
rect	142	136	143	137
rect	142	139	143	140
rect	142	142	143	143
rect	142	145	143	146
rect	142	148	143	149
rect	142	151	143	152
rect	142	154	143	155
rect	142	157	143	158
rect	142	160	143	161
rect	142	163	143	164
rect	142	166	143	167
rect	142	169	143	170
rect	142	172	143	173
rect	142	175	143	176
rect	142	178	143	179
rect	142	181	143	182
rect	142	184	143	185
rect	142	187	143	188
rect	142	190	143	191
rect	142	193	143	194
rect	142	196	143	197
rect	142	199	143	200
rect	142	202	143	203
rect	142	205	143	206
rect	142	208	143	209
rect	142	211	143	212
rect	142	214	143	215
rect	142	217	143	218
rect	142	220	143	221
rect	142	223	143	224
rect	142	226	143	227
rect	142	229	143	230
rect	142	232	143	233
rect	142	235	143	236
rect	142	238	143	239
rect	142	241	143	242
rect	142	244	143	245
rect	142	247	143	248
rect	142	250	143	251
rect	142	253	143	254
rect	142	256	143	257
rect	142	259	143	260
rect	142	262	143	263
rect	142	265	143	266
rect	142	268	143	269
rect	142	271	143	272
rect	142	274	143	275
rect	142	277	143	278
rect	142	280	143	281
rect	142	283	143	284
rect	142	286	143	287
rect	142	289	143	290
rect	142	292	143	293
rect	142	295	143	296
rect	142	298	143	299
rect	142	301	143	302
rect	142	304	143	305
rect	142	307	143	308
rect	142	310	143	311
rect	142	313	143	314
rect	142	316	143	317
rect	142	319	143	320
rect	142	322	143	323
rect	142	325	143	326
rect	142	328	143	329
rect	142	331	143	332
rect	142	334	143	335
rect	142	340	143	341
rect	142	343	143	344
rect	142	346	143	347
rect	142	349	143	350
rect	142	352	143	353
rect	142	355	143	356
rect	142	358	143	359
rect	142	361	143	362
rect	142	364	143	365
rect	142	367	143	368
rect	142	373	143	374
rect	142	376	143	377
rect	142	379	143	380
rect	142	385	143	386
rect	143	1	144	2
rect	143	4	144	5
rect	143	7	144	8
rect	143	10	144	11
rect	143	13	144	14
rect	143	16	144	17
rect	143	19	144	20
rect	143	22	144	23
rect	143	25	144	26
rect	143	28	144	29
rect	143	31	144	32
rect	143	34	144	35
rect	143	37	144	38
rect	143	40	144	41
rect	143	43	144	44
rect	143	46	144	47
rect	143	49	144	50
rect	143	52	144	53
rect	143	55	144	56
rect	143	58	144	59
rect	143	61	144	62
rect	143	64	144	65
rect	143	67	144	68
rect	143	70	144	71
rect	143	73	144	74
rect	143	76	144	77
rect	143	79	144	80
rect	143	82	144	83
rect	143	85	144	86
rect	143	88	144	89
rect	143	91	144	92
rect	143	94	144	95
rect	143	97	144	98
rect	143	100	144	101
rect	143	103	144	104
rect	143	106	144	107
rect	143	109	144	110
rect	143	112	144	113
rect	143	115	144	116
rect	143	118	144	119
rect	143	121	144	122
rect	143	124	144	125
rect	143	127	144	128
rect	143	130	144	131
rect	143	133	144	134
rect	143	136	144	137
rect	143	139	144	140
rect	143	142	144	143
rect	143	145	144	146
rect	143	148	144	149
rect	143	151	144	152
rect	143	154	144	155
rect	143	157	144	158
rect	143	160	144	161
rect	143	163	144	164
rect	143	166	144	167
rect	143	169	144	170
rect	143	172	144	173
rect	143	175	144	176
rect	143	178	144	179
rect	143	181	144	182
rect	143	184	144	185
rect	143	187	144	188
rect	143	190	144	191
rect	143	193	144	194
rect	143	196	144	197
rect	143	199	144	200
rect	143	202	144	203
rect	143	205	144	206
rect	143	208	144	209
rect	143	211	144	212
rect	143	214	144	215
rect	143	217	144	218
rect	143	220	144	221
rect	143	223	144	224
rect	143	226	144	227
rect	143	229	144	230
rect	143	232	144	233
rect	143	235	144	236
rect	143	238	144	239
rect	143	241	144	242
rect	143	244	144	245
rect	143	247	144	248
rect	143	250	144	251
rect	143	253	144	254
rect	143	256	144	257
rect	143	259	144	260
rect	143	262	144	263
rect	143	265	144	266
rect	143	268	144	269
rect	143	271	144	272
rect	143	274	144	275
rect	143	277	144	278
rect	143	280	144	281
rect	143	283	144	284
rect	143	286	144	287
rect	143	289	144	290
rect	143	292	144	293
rect	143	295	144	296
rect	143	298	144	299
rect	143	301	144	302
rect	143	307	144	308
rect	143	310	144	311
rect	143	313	144	314
rect	143	316	144	317
rect	143	319	144	320
rect	143	322	144	323
rect	143	325	144	326
rect	143	328	144	329
rect	143	331	144	332
rect	143	334	144	335
rect	143	340	144	341
rect	143	343	144	344
rect	143	346	144	347
rect	143	349	144	350
rect	143	352	144	353
rect	143	355	144	356
rect	143	358	144	359
rect	143	361	144	362
rect	143	364	144	365
rect	143	367	144	368
rect	143	373	144	374
rect	143	376	144	377
rect	143	379	144	380
rect	143	385	144	386
rect	144	1	145	2
rect	144	4	145	5
rect	144	7	145	8
rect	144	10	145	11
rect	144	13	145	14
rect	144	16	145	17
rect	144	19	145	20
rect	144	22	145	23
rect	144	25	145	26
rect	144	28	145	29
rect	144	31	145	32
rect	144	34	145	35
rect	144	37	145	38
rect	144	40	145	41
rect	144	43	145	44
rect	144	46	145	47
rect	144	49	145	50
rect	144	52	145	53
rect	144	55	145	56
rect	144	58	145	59
rect	144	61	145	62
rect	144	64	145	65
rect	144	67	145	68
rect	144	70	145	71
rect	144	73	145	74
rect	144	76	145	77
rect	144	79	145	80
rect	144	82	145	83
rect	144	85	145	86
rect	144	88	145	89
rect	144	91	145	92
rect	144	94	145	95
rect	144	97	145	98
rect	144	100	145	101
rect	144	103	145	104
rect	144	106	145	107
rect	144	109	145	110
rect	144	112	145	113
rect	144	115	145	116
rect	144	118	145	119
rect	144	121	145	122
rect	144	124	145	125
rect	144	127	145	128
rect	144	130	145	131
rect	144	133	145	134
rect	144	136	145	137
rect	144	139	145	140
rect	144	142	145	143
rect	144	145	145	146
rect	144	148	145	149
rect	144	151	145	152
rect	144	154	145	155
rect	144	157	145	158
rect	144	160	145	161
rect	144	163	145	164
rect	144	166	145	167
rect	144	169	145	170
rect	144	172	145	173
rect	144	175	145	176
rect	144	178	145	179
rect	144	181	145	182
rect	144	184	145	185
rect	144	187	145	188
rect	144	190	145	191
rect	144	193	145	194
rect	144	196	145	197
rect	144	199	145	200
rect	144	202	145	203
rect	144	205	145	206
rect	144	208	145	209
rect	144	211	145	212
rect	144	214	145	215
rect	144	217	145	218
rect	144	220	145	221
rect	144	223	145	224
rect	144	226	145	227
rect	144	229	145	230
rect	144	232	145	233
rect	144	235	145	236
rect	144	238	145	239
rect	144	241	145	242
rect	144	244	145	245
rect	144	247	145	248
rect	144	250	145	251
rect	144	253	145	254
rect	144	256	145	257
rect	144	259	145	260
rect	144	262	145	263
rect	144	265	145	266
rect	144	268	145	269
rect	144	271	145	272
rect	144	274	145	275
rect	144	277	145	278
rect	144	280	145	281
rect	144	283	145	284
rect	144	286	145	287
rect	144	289	145	290
rect	144	292	145	293
rect	144	295	145	296
rect	144	298	145	299
rect	144	301	145	302
rect	144	307	145	308
rect	144	310	145	311
rect	144	313	145	314
rect	144	316	145	317
rect	144	319	145	320
rect	144	322	145	323
rect	144	325	145	326
rect	144	328	145	329
rect	144	331	145	332
rect	144	334	145	335
rect	144	340	145	341
rect	144	343	145	344
rect	144	346	145	347
rect	144	349	145	350
rect	144	352	145	353
rect	144	355	145	356
rect	144	358	145	359
rect	144	361	145	362
rect	144	364	145	365
rect	144	367	145	368
rect	144	373	145	374
rect	144	376	145	377
rect	144	379	145	380
rect	144	385	145	386
rect	145	1	146	2
rect	145	4	146	5
rect	145	7	146	8
rect	145	10	146	11
rect	145	13	146	14
rect	145	16	146	17
rect	145	19	146	20
rect	145	22	146	23
rect	145	25	146	26
rect	145	28	146	29
rect	145	31	146	32
rect	145	34	146	35
rect	145	37	146	38
rect	145	40	146	41
rect	145	43	146	44
rect	145	46	146	47
rect	145	49	146	50
rect	145	52	146	53
rect	145	55	146	56
rect	145	58	146	59
rect	145	61	146	62
rect	145	64	146	65
rect	145	67	146	68
rect	145	70	146	71
rect	145	73	146	74
rect	145	76	146	77
rect	145	79	146	80
rect	145	82	146	83
rect	145	85	146	86
rect	145	88	146	89
rect	145	91	146	92
rect	145	94	146	95
rect	145	97	146	98
rect	145	100	146	101
rect	145	103	146	104
rect	145	106	146	107
rect	145	109	146	110
rect	145	112	146	113
rect	145	115	146	116
rect	145	118	146	119
rect	145	121	146	122
rect	145	124	146	125
rect	145	127	146	128
rect	145	130	146	131
rect	145	133	146	134
rect	145	136	146	137
rect	145	139	146	140
rect	145	142	146	143
rect	145	145	146	146
rect	145	148	146	149
rect	145	151	146	152
rect	145	154	146	155
rect	145	157	146	158
rect	145	160	146	161
rect	145	163	146	164
rect	145	166	146	167
rect	145	169	146	170
rect	145	172	146	173
rect	145	175	146	176
rect	145	178	146	179
rect	145	181	146	182
rect	145	184	146	185
rect	145	187	146	188
rect	145	190	146	191
rect	145	193	146	194
rect	145	196	146	197
rect	145	199	146	200
rect	145	202	146	203
rect	145	205	146	206
rect	145	208	146	209
rect	145	211	146	212
rect	145	214	146	215
rect	145	217	146	218
rect	145	220	146	221
rect	145	223	146	224
rect	145	226	146	227
rect	145	229	146	230
rect	145	232	146	233
rect	145	235	146	236
rect	145	238	146	239
rect	145	241	146	242
rect	145	244	146	245
rect	145	247	146	248
rect	145	250	146	251
rect	145	253	146	254
rect	145	256	146	257
rect	145	259	146	260
rect	145	262	146	263
rect	145	265	146	266
rect	145	268	146	269
rect	145	271	146	272
rect	145	274	146	275
rect	145	277	146	278
rect	145	280	146	281
rect	145	283	146	284
rect	145	286	146	287
rect	145	289	146	290
rect	145	292	146	293
rect	145	295	146	296
rect	145	298	146	299
rect	145	301	146	302
rect	145	307	146	308
rect	145	310	146	311
rect	145	313	146	314
rect	145	316	146	317
rect	145	319	146	320
rect	145	322	146	323
rect	145	325	146	326
rect	145	328	146	329
rect	145	331	146	332
rect	145	334	146	335
rect	145	340	146	341
rect	145	343	146	344
rect	145	346	146	347
rect	145	349	146	350
rect	145	352	146	353
rect	145	355	146	356
rect	145	358	146	359
rect	145	361	146	362
rect	145	364	146	365
rect	145	367	146	368
rect	145	373	146	374
rect	145	376	146	377
rect	145	379	146	380
rect	145	385	146	386
rect	146	1	147	2
rect	146	4	147	5
rect	146	7	147	8
rect	146	10	147	11
rect	146	13	147	14
rect	146	16	147	17
rect	146	19	147	20
rect	146	22	147	23
rect	146	25	147	26
rect	146	28	147	29
rect	146	31	147	32
rect	146	34	147	35
rect	146	37	147	38
rect	146	40	147	41
rect	146	43	147	44
rect	146	46	147	47
rect	146	49	147	50
rect	146	52	147	53
rect	146	55	147	56
rect	146	58	147	59
rect	146	61	147	62
rect	146	64	147	65
rect	146	67	147	68
rect	146	70	147	71
rect	146	73	147	74
rect	146	76	147	77
rect	146	79	147	80
rect	146	82	147	83
rect	146	85	147	86
rect	146	88	147	89
rect	146	91	147	92
rect	146	94	147	95
rect	146	97	147	98
rect	146	100	147	101
rect	146	103	147	104
rect	146	106	147	107
rect	146	109	147	110
rect	146	112	147	113
rect	146	115	147	116
rect	146	118	147	119
rect	146	121	147	122
rect	146	124	147	125
rect	146	127	147	128
rect	146	130	147	131
rect	146	133	147	134
rect	146	136	147	137
rect	146	139	147	140
rect	146	142	147	143
rect	146	145	147	146
rect	146	148	147	149
rect	146	151	147	152
rect	146	154	147	155
rect	146	157	147	158
rect	146	160	147	161
rect	146	163	147	164
rect	146	166	147	167
rect	146	169	147	170
rect	146	172	147	173
rect	146	175	147	176
rect	146	178	147	179
rect	146	181	147	182
rect	146	184	147	185
rect	146	187	147	188
rect	146	190	147	191
rect	146	193	147	194
rect	146	196	147	197
rect	146	199	147	200
rect	146	202	147	203
rect	146	205	147	206
rect	146	208	147	209
rect	146	211	147	212
rect	146	214	147	215
rect	146	217	147	218
rect	146	220	147	221
rect	146	223	147	224
rect	146	226	147	227
rect	146	229	147	230
rect	146	232	147	233
rect	146	235	147	236
rect	146	238	147	239
rect	146	241	147	242
rect	146	244	147	245
rect	146	247	147	248
rect	146	250	147	251
rect	146	253	147	254
rect	146	256	147	257
rect	146	259	147	260
rect	146	262	147	263
rect	146	265	147	266
rect	146	268	147	269
rect	146	271	147	272
rect	146	274	147	275
rect	146	277	147	278
rect	146	280	147	281
rect	146	283	147	284
rect	146	286	147	287
rect	146	289	147	290
rect	146	292	147	293
rect	146	295	147	296
rect	146	298	147	299
rect	146	301	147	302
rect	146	307	147	308
rect	146	310	147	311
rect	146	313	147	314
rect	146	316	147	317
rect	146	319	147	320
rect	146	322	147	323
rect	146	325	147	326
rect	146	328	147	329
rect	146	331	147	332
rect	146	334	147	335
rect	146	340	147	341
rect	146	343	147	344
rect	146	346	147	347
rect	146	349	147	350
rect	146	352	147	353
rect	146	355	147	356
rect	146	358	147	359
rect	146	361	147	362
rect	146	364	147	365
rect	146	367	147	368
rect	146	373	147	374
rect	146	376	147	377
rect	146	379	147	380
rect	146	385	147	386
rect	147	1	148	2
rect	147	4	148	5
rect	147	7	148	8
rect	147	10	148	11
rect	147	13	148	14
rect	147	16	148	17
rect	147	19	148	20
rect	147	22	148	23
rect	147	25	148	26
rect	147	28	148	29
rect	147	31	148	32
rect	147	34	148	35
rect	147	37	148	38
rect	147	40	148	41
rect	147	43	148	44
rect	147	46	148	47
rect	147	49	148	50
rect	147	52	148	53
rect	147	55	148	56
rect	147	58	148	59
rect	147	61	148	62
rect	147	64	148	65
rect	147	67	148	68
rect	147	70	148	71
rect	147	73	148	74
rect	147	76	148	77
rect	147	79	148	80
rect	147	82	148	83
rect	147	85	148	86
rect	147	88	148	89
rect	147	91	148	92
rect	147	94	148	95
rect	147	97	148	98
rect	147	100	148	101
rect	147	103	148	104
rect	147	106	148	107
rect	147	109	148	110
rect	147	112	148	113
rect	147	115	148	116
rect	147	118	148	119
rect	147	121	148	122
rect	147	124	148	125
rect	147	127	148	128
rect	147	130	148	131
rect	147	133	148	134
rect	147	136	148	137
rect	147	139	148	140
rect	147	142	148	143
rect	147	145	148	146
rect	147	148	148	149
rect	147	151	148	152
rect	147	154	148	155
rect	147	157	148	158
rect	147	160	148	161
rect	147	163	148	164
rect	147	166	148	167
rect	147	169	148	170
rect	147	172	148	173
rect	147	175	148	176
rect	147	178	148	179
rect	147	181	148	182
rect	147	184	148	185
rect	147	187	148	188
rect	147	190	148	191
rect	147	193	148	194
rect	147	196	148	197
rect	147	199	148	200
rect	147	202	148	203
rect	147	205	148	206
rect	147	208	148	209
rect	147	211	148	212
rect	147	214	148	215
rect	147	217	148	218
rect	147	220	148	221
rect	147	223	148	224
rect	147	226	148	227
rect	147	229	148	230
rect	147	232	148	233
rect	147	235	148	236
rect	147	238	148	239
rect	147	241	148	242
rect	147	244	148	245
rect	147	247	148	248
rect	147	250	148	251
rect	147	253	148	254
rect	147	256	148	257
rect	147	259	148	260
rect	147	262	148	263
rect	147	265	148	266
rect	147	268	148	269
rect	147	271	148	272
rect	147	274	148	275
rect	147	277	148	278
rect	147	280	148	281
rect	147	283	148	284
rect	147	286	148	287
rect	147	289	148	290
rect	147	292	148	293
rect	147	295	148	296
rect	147	298	148	299
rect	147	301	148	302
rect	147	307	148	308
rect	147	310	148	311
rect	147	313	148	314
rect	147	316	148	317
rect	147	319	148	320
rect	147	322	148	323
rect	147	325	148	326
rect	147	328	148	329
rect	147	331	148	332
rect	147	334	148	335
rect	147	340	148	341
rect	147	343	148	344
rect	147	346	148	347
rect	147	349	148	350
rect	147	352	148	353
rect	147	355	148	356
rect	147	358	148	359
rect	147	361	148	362
rect	147	364	148	365
rect	147	367	148	368
rect	147	373	148	374
rect	147	376	148	377
rect	147	379	148	380
rect	147	385	148	386
rect	148	1	149	2
rect	148	4	149	5
rect	148	7	149	8
rect	148	10	149	11
rect	148	13	149	14
rect	148	16	149	17
rect	148	19	149	20
rect	148	22	149	23
rect	148	25	149	26
rect	148	28	149	29
rect	148	31	149	32
rect	148	34	149	35
rect	148	37	149	38
rect	148	40	149	41
rect	148	43	149	44
rect	148	46	149	47
rect	148	49	149	50
rect	148	52	149	53
rect	148	55	149	56
rect	148	58	149	59
rect	148	61	149	62
rect	148	64	149	65
rect	148	67	149	68
rect	148	70	149	71
rect	148	73	149	74
rect	148	76	149	77
rect	148	79	149	80
rect	148	82	149	83
rect	148	85	149	86
rect	148	88	149	89
rect	148	91	149	92
rect	148	94	149	95
rect	148	97	149	98
rect	148	100	149	101
rect	148	103	149	104
rect	148	106	149	107
rect	148	109	149	110
rect	148	112	149	113
rect	148	115	149	116
rect	148	118	149	119
rect	148	121	149	122
rect	148	124	149	125
rect	148	127	149	128
rect	148	130	149	131
rect	148	133	149	134
rect	148	136	149	137
rect	148	139	149	140
rect	148	142	149	143
rect	148	145	149	146
rect	148	148	149	149
rect	148	151	149	152
rect	148	154	149	155
rect	148	157	149	158
rect	148	160	149	161
rect	148	163	149	164
rect	148	166	149	167
rect	148	169	149	170
rect	148	172	149	173
rect	148	175	149	176
rect	148	178	149	179
rect	148	181	149	182
rect	148	184	149	185
rect	148	187	149	188
rect	148	190	149	191
rect	148	193	149	194
rect	148	196	149	197
rect	148	199	149	200
rect	148	202	149	203
rect	148	205	149	206
rect	148	208	149	209
rect	148	211	149	212
rect	148	214	149	215
rect	148	217	149	218
rect	148	220	149	221
rect	148	223	149	224
rect	148	226	149	227
rect	148	229	149	230
rect	148	232	149	233
rect	148	235	149	236
rect	148	238	149	239
rect	148	241	149	242
rect	148	244	149	245
rect	148	247	149	248
rect	148	250	149	251
rect	148	253	149	254
rect	148	256	149	257
rect	148	259	149	260
rect	148	262	149	263
rect	148	265	149	266
rect	148	268	149	269
rect	148	271	149	272
rect	148	274	149	275
rect	148	277	149	278
rect	148	280	149	281
rect	148	283	149	284
rect	148	286	149	287
rect	148	289	149	290
rect	148	292	149	293
rect	148	295	149	296
rect	148	298	149	299
rect	148	301	149	302
rect	148	307	149	308
rect	148	310	149	311
rect	148	313	149	314
rect	148	316	149	317
rect	148	319	149	320
rect	148	322	149	323
rect	148	325	149	326
rect	148	328	149	329
rect	148	331	149	332
rect	148	334	149	335
rect	148	340	149	341
rect	148	343	149	344
rect	148	346	149	347
rect	148	349	149	350
rect	148	352	149	353
rect	148	355	149	356
rect	148	358	149	359
rect	148	361	149	362
rect	148	364	149	365
rect	148	367	149	368
rect	148	373	149	374
rect	148	376	149	377
rect	148	379	149	380
rect	148	385	149	386
rect	149	1	150	2
rect	149	4	150	5
rect	149	7	150	8
rect	149	10	150	11
rect	149	13	150	14
rect	149	16	150	17
rect	149	19	150	20
rect	149	22	150	23
rect	149	25	150	26
rect	149	28	150	29
rect	149	31	150	32
rect	149	34	150	35
rect	149	37	150	38
rect	149	40	150	41
rect	149	43	150	44
rect	149	46	150	47
rect	149	49	150	50
rect	149	52	150	53
rect	149	55	150	56
rect	149	58	150	59
rect	149	61	150	62
rect	149	64	150	65
rect	149	67	150	68
rect	149	70	150	71
rect	149	73	150	74
rect	149	76	150	77
rect	149	79	150	80
rect	149	82	150	83
rect	149	85	150	86
rect	149	88	150	89
rect	149	91	150	92
rect	149	94	150	95
rect	149	97	150	98
rect	149	100	150	101
rect	149	103	150	104
rect	149	106	150	107
rect	149	109	150	110
rect	149	112	150	113
rect	149	115	150	116
rect	149	118	150	119
rect	149	121	150	122
rect	149	124	150	125
rect	149	127	150	128
rect	149	130	150	131
rect	149	133	150	134
rect	149	136	150	137
rect	149	139	150	140
rect	149	142	150	143
rect	149	145	150	146
rect	149	148	150	149
rect	149	151	150	152
rect	149	154	150	155
rect	149	157	150	158
rect	149	160	150	161
rect	149	163	150	164
rect	149	166	150	167
rect	149	169	150	170
rect	149	172	150	173
rect	149	175	150	176
rect	149	178	150	179
rect	149	181	150	182
rect	149	184	150	185
rect	149	187	150	188
rect	149	190	150	191
rect	149	193	150	194
rect	149	196	150	197
rect	149	199	150	200
rect	149	202	150	203
rect	149	205	150	206
rect	149	208	150	209
rect	149	211	150	212
rect	149	214	150	215
rect	149	217	150	218
rect	149	220	150	221
rect	149	223	150	224
rect	149	226	150	227
rect	149	229	150	230
rect	149	232	150	233
rect	149	235	150	236
rect	149	238	150	239
rect	149	241	150	242
rect	149	244	150	245
rect	149	247	150	248
rect	149	250	150	251
rect	149	253	150	254
rect	149	256	150	257
rect	149	259	150	260
rect	149	262	150	263
rect	149	265	150	266
rect	149	268	150	269
rect	149	271	150	272
rect	149	274	150	275
rect	149	277	150	278
rect	149	280	150	281
rect	149	283	150	284
rect	149	286	150	287
rect	149	289	150	290
rect	149	292	150	293
rect	149	295	150	296
rect	149	298	150	299
rect	149	301	150	302
rect	149	307	150	308
rect	149	310	150	311
rect	149	313	150	314
rect	149	316	150	317
rect	149	319	150	320
rect	149	322	150	323
rect	149	325	150	326
rect	149	328	150	329
rect	149	331	150	332
rect	149	334	150	335
rect	149	340	150	341
rect	149	343	150	344
rect	149	346	150	347
rect	149	349	150	350
rect	149	352	150	353
rect	149	355	150	356
rect	149	358	150	359
rect	149	361	150	362
rect	149	364	150	365
rect	149	367	150	368
rect	149	373	150	374
rect	149	376	150	377
rect	149	379	150	380
rect	149	385	150	386
rect	150	1	151	2
rect	150	4	151	5
rect	150	7	151	8
rect	150	10	151	11
rect	150	13	151	14
rect	150	16	151	17
rect	150	19	151	20
rect	150	22	151	23
rect	150	25	151	26
rect	150	28	151	29
rect	150	31	151	32
rect	150	34	151	35
rect	150	37	151	38
rect	150	40	151	41
rect	150	43	151	44
rect	150	46	151	47
rect	150	49	151	50
rect	150	52	151	53
rect	150	55	151	56
rect	150	58	151	59
rect	150	61	151	62
rect	150	64	151	65
rect	150	67	151	68
rect	150	70	151	71
rect	150	73	151	74
rect	150	76	151	77
rect	150	79	151	80
rect	150	82	151	83
rect	150	85	151	86
rect	150	88	151	89
rect	150	91	151	92
rect	150	94	151	95
rect	150	97	151	98
rect	150	100	151	101
rect	150	103	151	104
rect	150	106	151	107
rect	150	109	151	110
rect	150	112	151	113
rect	150	115	151	116
rect	150	118	151	119
rect	150	121	151	122
rect	150	124	151	125
rect	150	127	151	128
rect	150	130	151	131
rect	150	133	151	134
rect	150	136	151	137
rect	150	139	151	140
rect	150	142	151	143
rect	150	145	151	146
rect	150	148	151	149
rect	150	151	151	152
rect	150	154	151	155
rect	150	157	151	158
rect	150	160	151	161
rect	150	163	151	164
rect	150	166	151	167
rect	150	169	151	170
rect	150	172	151	173
rect	150	175	151	176
rect	150	178	151	179
rect	150	181	151	182
rect	150	184	151	185
rect	150	187	151	188
rect	150	190	151	191
rect	150	193	151	194
rect	150	196	151	197
rect	150	199	151	200
rect	150	202	151	203
rect	150	205	151	206
rect	150	208	151	209
rect	150	211	151	212
rect	150	214	151	215
rect	150	217	151	218
rect	150	220	151	221
rect	150	223	151	224
rect	150	226	151	227
rect	150	229	151	230
rect	150	232	151	233
rect	150	235	151	236
rect	150	238	151	239
rect	150	241	151	242
rect	150	244	151	245
rect	150	247	151	248
rect	150	250	151	251
rect	150	253	151	254
rect	150	256	151	257
rect	150	259	151	260
rect	150	262	151	263
rect	150	265	151	266
rect	150	268	151	269
rect	150	271	151	272
rect	150	274	151	275
rect	150	277	151	278
rect	150	280	151	281
rect	150	283	151	284
rect	150	286	151	287
rect	150	289	151	290
rect	150	292	151	293
rect	150	295	151	296
rect	150	298	151	299
rect	150	301	151	302
rect	150	307	151	308
rect	150	310	151	311
rect	150	313	151	314
rect	150	316	151	317
rect	150	319	151	320
rect	150	322	151	323
rect	150	325	151	326
rect	150	328	151	329
rect	150	331	151	332
rect	150	334	151	335
rect	150	340	151	341
rect	150	343	151	344
rect	150	346	151	347
rect	150	349	151	350
rect	150	352	151	353
rect	150	355	151	356
rect	150	358	151	359
rect	150	361	151	362
rect	150	364	151	365
rect	150	367	151	368
rect	150	373	151	374
rect	150	376	151	377
rect	150	379	151	380
rect	150	385	151	386
rect	151	1	152	2
rect	151	4	152	5
rect	151	7	152	8
rect	151	10	152	11
rect	151	13	152	14
rect	151	16	152	17
rect	151	19	152	20
rect	151	22	152	23
rect	151	25	152	26
rect	151	28	152	29
rect	151	31	152	32
rect	151	34	152	35
rect	151	37	152	38
rect	151	40	152	41
rect	151	43	152	44
rect	151	46	152	47
rect	151	49	152	50
rect	151	52	152	53
rect	151	55	152	56
rect	151	58	152	59
rect	151	61	152	62
rect	151	64	152	65
rect	151	67	152	68
rect	151	70	152	71
rect	151	73	152	74
rect	151	76	152	77
rect	151	79	152	80
rect	151	82	152	83
rect	151	85	152	86
rect	151	88	152	89
rect	151	91	152	92
rect	151	94	152	95
rect	151	97	152	98
rect	151	100	152	101
rect	151	103	152	104
rect	151	106	152	107
rect	151	109	152	110
rect	151	112	152	113
rect	151	115	152	116
rect	151	118	152	119
rect	151	121	152	122
rect	151	124	152	125
rect	151	127	152	128
rect	151	130	152	131
rect	151	133	152	134
rect	151	136	152	137
rect	151	139	152	140
rect	151	142	152	143
rect	151	145	152	146
rect	151	148	152	149
rect	151	151	152	152
rect	151	154	152	155
rect	151	157	152	158
rect	151	160	152	161
rect	151	163	152	164
rect	151	166	152	167
rect	151	169	152	170
rect	151	172	152	173
rect	151	175	152	176
rect	151	178	152	179
rect	151	181	152	182
rect	151	184	152	185
rect	151	187	152	188
rect	151	190	152	191
rect	151	193	152	194
rect	151	196	152	197
rect	151	199	152	200
rect	151	202	152	203
rect	151	205	152	206
rect	151	208	152	209
rect	151	211	152	212
rect	151	214	152	215
rect	151	217	152	218
rect	151	220	152	221
rect	151	223	152	224
rect	151	226	152	227
rect	151	229	152	230
rect	151	232	152	233
rect	151	235	152	236
rect	151	238	152	239
rect	151	241	152	242
rect	151	244	152	245
rect	151	247	152	248
rect	151	250	152	251
rect	151	253	152	254
rect	151	256	152	257
rect	151	259	152	260
rect	151	262	152	263
rect	151	265	152	266
rect	151	268	152	269
rect	151	271	152	272
rect	151	274	152	275
rect	151	277	152	278
rect	151	280	152	281
rect	151	283	152	284
rect	151	286	152	287
rect	151	289	152	290
rect	151	292	152	293
rect	151	295	152	296
rect	151	298	152	299
rect	151	301	152	302
rect	151	307	152	308
rect	151	310	152	311
rect	151	313	152	314
rect	151	316	152	317
rect	151	319	152	320
rect	151	322	152	323
rect	151	325	152	326
rect	151	328	152	329
rect	151	331	152	332
rect	151	334	152	335
rect	151	340	152	341
rect	151	343	152	344
rect	151	346	152	347
rect	151	349	152	350
rect	151	352	152	353
rect	151	355	152	356
rect	151	358	152	359
rect	151	361	152	362
rect	151	364	152	365
rect	151	367	152	368
rect	151	373	152	374
rect	151	376	152	377
rect	151	379	152	380
rect	151	385	152	386
rect	152	1	153	2
rect	152	4	153	5
rect	152	7	153	8
rect	152	10	153	11
rect	152	13	153	14
rect	152	16	153	17
rect	152	19	153	20
rect	152	22	153	23
rect	152	25	153	26
rect	152	28	153	29
rect	152	31	153	32
rect	152	34	153	35
rect	152	37	153	38
rect	152	40	153	41
rect	152	43	153	44
rect	152	46	153	47
rect	152	49	153	50
rect	152	52	153	53
rect	152	55	153	56
rect	152	58	153	59
rect	152	61	153	62
rect	152	64	153	65
rect	152	67	153	68
rect	152	70	153	71
rect	152	73	153	74
rect	152	76	153	77
rect	152	79	153	80
rect	152	82	153	83
rect	152	85	153	86
rect	152	88	153	89
rect	152	91	153	92
rect	152	94	153	95
rect	152	97	153	98
rect	152	100	153	101
rect	152	103	153	104
rect	152	106	153	107
rect	152	109	153	110
rect	152	112	153	113
rect	152	115	153	116
rect	152	118	153	119
rect	152	121	153	122
rect	152	124	153	125
rect	152	127	153	128
rect	152	130	153	131
rect	152	133	153	134
rect	152	136	153	137
rect	152	142	153	143
rect	152	145	153	146
rect	152	148	153	149
rect	152	151	153	152
rect	152	154	153	155
rect	152	157	153	158
rect	152	160	153	161
rect	152	163	153	164
rect	152	166	153	167
rect	152	169	153	170
rect	152	172	153	173
rect	152	175	153	176
rect	152	178	153	179
rect	152	181	153	182
rect	152	184	153	185
rect	152	187	153	188
rect	152	190	153	191
rect	152	193	153	194
rect	152	196	153	197
rect	152	199	153	200
rect	152	202	153	203
rect	152	205	153	206
rect	152	208	153	209
rect	152	211	153	212
rect	152	214	153	215
rect	152	217	153	218
rect	152	220	153	221
rect	152	223	153	224
rect	152	226	153	227
rect	152	229	153	230
rect	152	232	153	233
rect	152	235	153	236
rect	152	238	153	239
rect	152	241	153	242
rect	152	244	153	245
rect	152	247	153	248
rect	152	250	153	251
rect	152	253	153	254
rect	152	256	153	257
rect	152	259	153	260
rect	152	262	153	263
rect	152	265	153	266
rect	152	268	153	269
rect	152	271	153	272
rect	152	274	153	275
rect	152	277	153	278
rect	152	280	153	281
rect	152	283	153	284
rect	152	286	153	287
rect	152	289	153	290
rect	152	292	153	293
rect	152	295	153	296
rect	152	298	153	299
rect	152	301	153	302
rect	152	307	153	308
rect	152	310	153	311
rect	152	313	153	314
rect	152	316	153	317
rect	152	319	153	320
rect	152	322	153	323
rect	152	325	153	326
rect	152	328	153	329
rect	152	331	153	332
rect	152	334	153	335
rect	152	340	153	341
rect	152	343	153	344
rect	152	346	153	347
rect	152	349	153	350
rect	152	352	153	353
rect	152	355	153	356
rect	152	358	153	359
rect	152	361	153	362
rect	152	364	153	365
rect	152	367	153	368
rect	152	373	153	374
rect	152	376	153	377
rect	152	379	153	380
rect	152	385	153	386
rect	153	1	154	2
rect	153	4	154	5
rect	153	7	154	8
rect	153	10	154	11
rect	153	13	154	14
rect	153	16	154	17
rect	153	19	154	20
rect	153	22	154	23
rect	153	25	154	26
rect	153	28	154	29
rect	153	31	154	32
rect	153	34	154	35
rect	153	37	154	38
rect	153	40	154	41
rect	153	43	154	44
rect	153	46	154	47
rect	153	49	154	50
rect	153	52	154	53
rect	153	55	154	56
rect	153	58	154	59
rect	153	61	154	62
rect	153	64	154	65
rect	153	67	154	68
rect	153	70	154	71
rect	153	73	154	74
rect	153	76	154	77
rect	153	79	154	80
rect	153	82	154	83
rect	153	85	154	86
rect	153	88	154	89
rect	153	91	154	92
rect	153	94	154	95
rect	153	97	154	98
rect	153	100	154	101
rect	153	103	154	104
rect	153	106	154	107
rect	153	109	154	110
rect	153	112	154	113
rect	153	115	154	116
rect	153	118	154	119
rect	153	121	154	122
rect	153	124	154	125
rect	153	127	154	128
rect	153	130	154	131
rect	153	133	154	134
rect	153	136	154	137
rect	153	139	154	140
rect	153	142	154	143
rect	153	145	154	146
rect	153	148	154	149
rect	153	151	154	152
rect	153	154	154	155
rect	153	157	154	158
rect	153	160	154	161
rect	153	163	154	164
rect	153	166	154	167
rect	153	169	154	170
rect	153	172	154	173
rect	153	175	154	176
rect	153	178	154	179
rect	153	181	154	182
rect	153	184	154	185
rect	153	187	154	188
rect	153	190	154	191
rect	153	193	154	194
rect	153	196	154	197
rect	153	199	154	200
rect	153	202	154	203
rect	153	205	154	206
rect	153	208	154	209
rect	153	211	154	212
rect	153	214	154	215
rect	153	217	154	218
rect	153	220	154	221
rect	153	223	154	224
rect	153	226	154	227
rect	153	229	154	230
rect	153	232	154	233
rect	153	235	154	236
rect	153	238	154	239
rect	153	241	154	242
rect	153	244	154	245
rect	153	247	154	248
rect	153	250	154	251
rect	153	253	154	254
rect	153	256	154	257
rect	153	259	154	260
rect	153	262	154	263
rect	153	265	154	266
rect	153	268	154	269
rect	153	271	154	272
rect	153	274	154	275
rect	153	277	154	278
rect	153	280	154	281
rect	153	283	154	284
rect	153	286	154	287
rect	153	289	154	290
rect	153	292	154	293
rect	153	295	154	296
rect	153	298	154	299
rect	153	301	154	302
rect	153	307	154	308
rect	153	310	154	311
rect	153	313	154	314
rect	153	316	154	317
rect	153	319	154	320
rect	153	322	154	323
rect	153	325	154	326
rect	153	328	154	329
rect	153	331	154	332
rect	153	334	154	335
rect	153	340	154	341
rect	153	343	154	344
rect	153	346	154	347
rect	153	349	154	350
rect	153	352	154	353
rect	153	355	154	356
rect	153	358	154	359
rect	153	361	154	362
rect	153	364	154	365
rect	153	367	154	368
rect	153	373	154	374
rect	153	376	154	377
rect	153	379	154	380
rect	153	385	154	386
rect	154	1	155	2
rect	154	4	155	5
rect	154	7	155	8
rect	154	10	155	11
rect	154	13	155	14
rect	154	16	155	17
rect	154	19	155	20
rect	154	22	155	23
rect	154	25	155	26
rect	154	28	155	29
rect	154	31	155	32
rect	154	34	155	35
rect	154	37	155	38
rect	154	40	155	41
rect	154	43	155	44
rect	154	46	155	47
rect	154	49	155	50
rect	154	52	155	53
rect	154	55	155	56
rect	154	58	155	59
rect	154	61	155	62
rect	154	64	155	65
rect	154	67	155	68
rect	154	70	155	71
rect	154	73	155	74
rect	154	76	155	77
rect	154	79	155	80
rect	154	82	155	83
rect	154	85	155	86
rect	154	88	155	89
rect	154	91	155	92
rect	154	94	155	95
rect	154	97	155	98
rect	154	100	155	101
rect	154	103	155	104
rect	154	106	155	107
rect	154	109	155	110
rect	154	112	155	113
rect	154	115	155	116
rect	154	118	155	119
rect	154	121	155	122
rect	154	124	155	125
rect	154	127	155	128
rect	154	130	155	131
rect	154	133	155	134
rect	154	136	155	137
rect	154	139	155	140
rect	154	142	155	143
rect	154	145	155	146
rect	154	148	155	149
rect	154	151	155	152
rect	154	154	155	155
rect	154	157	155	158
rect	154	160	155	161
rect	154	163	155	164
rect	154	166	155	167
rect	154	169	155	170
rect	154	172	155	173
rect	154	175	155	176
rect	154	178	155	179
rect	154	181	155	182
rect	154	184	155	185
rect	154	187	155	188
rect	154	190	155	191
rect	154	193	155	194
rect	154	196	155	197
rect	154	199	155	200
rect	154	202	155	203
rect	154	205	155	206
rect	154	208	155	209
rect	154	211	155	212
rect	154	214	155	215
rect	154	217	155	218
rect	154	220	155	221
rect	154	223	155	224
rect	154	226	155	227
rect	154	229	155	230
rect	154	232	155	233
rect	154	235	155	236
rect	154	238	155	239
rect	154	241	155	242
rect	154	244	155	245
rect	154	247	155	248
rect	154	250	155	251
rect	154	253	155	254
rect	154	256	155	257
rect	154	259	155	260
rect	154	262	155	263
rect	154	265	155	266
rect	154	268	155	269
rect	154	271	155	272
rect	154	274	155	275
rect	154	277	155	278
rect	154	280	155	281
rect	154	283	155	284
rect	154	286	155	287
rect	154	289	155	290
rect	154	292	155	293
rect	154	295	155	296
rect	154	298	155	299
rect	154	301	155	302
rect	154	307	155	308
rect	154	310	155	311
rect	154	313	155	314
rect	154	316	155	317
rect	154	319	155	320
rect	154	322	155	323
rect	154	325	155	326
rect	154	328	155	329
rect	154	331	155	332
rect	154	334	155	335
rect	154	340	155	341
rect	154	343	155	344
rect	154	349	155	350
rect	154	352	155	353
rect	154	355	155	356
rect	154	358	155	359
rect	154	361	155	362
rect	154	364	155	365
rect	154	367	155	368
rect	154	373	155	374
rect	154	376	155	377
rect	154	379	155	380
rect	154	385	155	386
rect	155	1	156	2
rect	155	4	156	5
rect	155	7	156	8
rect	155	10	156	11
rect	155	13	156	14
rect	155	16	156	17
rect	155	19	156	20
rect	155	22	156	23
rect	155	25	156	26
rect	155	28	156	29
rect	155	31	156	32
rect	155	34	156	35
rect	155	37	156	38
rect	155	40	156	41
rect	155	43	156	44
rect	155	46	156	47
rect	155	49	156	50
rect	155	52	156	53
rect	155	55	156	56
rect	155	58	156	59
rect	155	61	156	62
rect	155	64	156	65
rect	155	67	156	68
rect	155	70	156	71
rect	155	73	156	74
rect	155	76	156	77
rect	155	79	156	80
rect	155	82	156	83
rect	155	85	156	86
rect	155	88	156	89
rect	155	91	156	92
rect	155	94	156	95
rect	155	97	156	98
rect	155	100	156	101
rect	155	103	156	104
rect	155	106	156	107
rect	155	109	156	110
rect	155	112	156	113
rect	155	115	156	116
rect	155	118	156	119
rect	155	121	156	122
rect	155	124	156	125
rect	155	127	156	128
rect	155	130	156	131
rect	155	133	156	134
rect	155	136	156	137
rect	155	139	156	140
rect	155	142	156	143
rect	155	145	156	146
rect	155	148	156	149
rect	155	151	156	152
rect	155	154	156	155
rect	155	157	156	158
rect	155	160	156	161
rect	155	163	156	164
rect	155	166	156	167
rect	155	169	156	170
rect	155	172	156	173
rect	155	175	156	176
rect	155	178	156	179
rect	155	181	156	182
rect	155	184	156	185
rect	155	187	156	188
rect	155	190	156	191
rect	155	193	156	194
rect	155	196	156	197
rect	155	199	156	200
rect	155	202	156	203
rect	155	205	156	206
rect	155	208	156	209
rect	155	211	156	212
rect	155	214	156	215
rect	155	217	156	218
rect	155	220	156	221
rect	155	223	156	224
rect	155	226	156	227
rect	155	229	156	230
rect	155	232	156	233
rect	155	235	156	236
rect	155	238	156	239
rect	155	241	156	242
rect	155	244	156	245
rect	155	247	156	248
rect	155	250	156	251
rect	155	253	156	254
rect	155	256	156	257
rect	155	259	156	260
rect	155	262	156	263
rect	155	265	156	266
rect	155	268	156	269
rect	155	271	156	272
rect	155	274	156	275
rect	155	277	156	278
rect	155	280	156	281
rect	155	283	156	284
rect	155	286	156	287
rect	155	289	156	290
rect	155	292	156	293
rect	155	295	156	296
rect	155	298	156	299
rect	155	301	156	302
rect	155	307	156	308
rect	155	310	156	311
rect	155	313	156	314
rect	155	316	156	317
rect	155	319	156	320
rect	155	322	156	323
rect	155	325	156	326
rect	155	328	156	329
rect	155	331	156	332
rect	155	334	156	335
rect	155	343	156	344
rect	155	346	156	347
rect	155	349	156	350
rect	155	352	156	353
rect	155	355	156	356
rect	155	358	156	359
rect	155	361	156	362
rect	155	364	156	365
rect	155	367	156	368
rect	155	373	156	374
rect	155	376	156	377
rect	155	379	156	380
rect	155	385	156	386
rect	156	1	157	2
rect	156	4	157	5
rect	156	7	157	8
rect	156	10	157	11
rect	156	13	157	14
rect	156	16	157	17
rect	156	19	157	20
rect	156	22	157	23
rect	156	25	157	26
rect	156	28	157	29
rect	156	31	157	32
rect	156	34	157	35
rect	156	37	157	38
rect	156	40	157	41
rect	156	43	157	44
rect	156	46	157	47
rect	156	49	157	50
rect	156	52	157	53
rect	156	55	157	56
rect	156	58	157	59
rect	156	61	157	62
rect	156	64	157	65
rect	156	67	157	68
rect	156	70	157	71
rect	156	73	157	74
rect	156	76	157	77
rect	156	79	157	80
rect	156	82	157	83
rect	156	85	157	86
rect	156	88	157	89
rect	156	91	157	92
rect	156	94	157	95
rect	156	97	157	98
rect	156	100	157	101
rect	156	103	157	104
rect	156	106	157	107
rect	156	109	157	110
rect	156	112	157	113
rect	156	115	157	116
rect	156	118	157	119
rect	156	121	157	122
rect	156	124	157	125
rect	156	127	157	128
rect	156	130	157	131
rect	156	133	157	134
rect	156	136	157	137
rect	156	139	157	140
rect	156	142	157	143
rect	156	145	157	146
rect	156	148	157	149
rect	156	151	157	152
rect	156	154	157	155
rect	156	157	157	158
rect	156	160	157	161
rect	156	163	157	164
rect	156	166	157	167
rect	156	169	157	170
rect	156	172	157	173
rect	156	175	157	176
rect	156	178	157	179
rect	156	181	157	182
rect	156	184	157	185
rect	156	187	157	188
rect	156	190	157	191
rect	156	193	157	194
rect	156	196	157	197
rect	156	199	157	200
rect	156	202	157	203
rect	156	205	157	206
rect	156	208	157	209
rect	156	211	157	212
rect	156	214	157	215
rect	156	217	157	218
rect	156	220	157	221
rect	156	223	157	224
rect	156	226	157	227
rect	156	229	157	230
rect	156	232	157	233
rect	156	235	157	236
rect	156	238	157	239
rect	156	241	157	242
rect	156	244	157	245
rect	156	247	157	248
rect	156	250	157	251
rect	156	253	157	254
rect	156	256	157	257
rect	156	259	157	260
rect	156	262	157	263
rect	156	265	157	266
rect	156	268	157	269
rect	156	271	157	272
rect	156	274	157	275
rect	156	277	157	278
rect	156	280	157	281
rect	156	283	157	284
rect	156	286	157	287
rect	156	289	157	290
rect	156	292	157	293
rect	156	298	157	299
rect	156	301	157	302
rect	156	307	157	308
rect	156	310	157	311
rect	156	313	157	314
rect	156	316	157	317
rect	156	319	157	320
rect	156	322	157	323
rect	156	325	157	326
rect	156	328	157	329
rect	156	331	157	332
rect	156	334	157	335
rect	156	343	157	344
rect	156	346	157	347
rect	156	349	157	350
rect	156	352	157	353
rect	156	355	157	356
rect	156	358	157	359
rect	156	361	157	362
rect	156	364	157	365
rect	156	367	157	368
rect	156	373	157	374
rect	156	376	157	377
rect	156	379	157	380
rect	156	385	157	386
rect	157	1	158	2
rect	157	4	158	5
rect	157	7	158	8
rect	157	10	158	11
rect	157	13	158	14
rect	157	16	158	17
rect	157	19	158	20
rect	157	22	158	23
rect	157	25	158	26
rect	157	28	158	29
rect	157	31	158	32
rect	157	34	158	35
rect	157	37	158	38
rect	157	40	158	41
rect	157	43	158	44
rect	157	46	158	47
rect	157	49	158	50
rect	157	52	158	53
rect	157	55	158	56
rect	157	58	158	59
rect	157	61	158	62
rect	157	64	158	65
rect	157	67	158	68
rect	157	70	158	71
rect	157	73	158	74
rect	157	76	158	77
rect	157	79	158	80
rect	157	82	158	83
rect	157	85	158	86
rect	157	88	158	89
rect	157	91	158	92
rect	157	94	158	95
rect	157	97	158	98
rect	157	100	158	101
rect	157	103	158	104
rect	157	106	158	107
rect	157	109	158	110
rect	157	112	158	113
rect	157	115	158	116
rect	157	118	158	119
rect	157	121	158	122
rect	157	124	158	125
rect	157	127	158	128
rect	157	130	158	131
rect	157	133	158	134
rect	157	136	158	137
rect	157	139	158	140
rect	157	142	158	143
rect	157	145	158	146
rect	157	148	158	149
rect	157	151	158	152
rect	157	154	158	155
rect	157	157	158	158
rect	157	160	158	161
rect	157	163	158	164
rect	157	166	158	167
rect	157	169	158	170
rect	157	172	158	173
rect	157	175	158	176
rect	157	178	158	179
rect	157	181	158	182
rect	157	184	158	185
rect	157	187	158	188
rect	157	190	158	191
rect	157	193	158	194
rect	157	196	158	197
rect	157	199	158	200
rect	157	202	158	203
rect	157	205	158	206
rect	157	208	158	209
rect	157	211	158	212
rect	157	214	158	215
rect	157	217	158	218
rect	157	220	158	221
rect	157	223	158	224
rect	157	226	158	227
rect	157	229	158	230
rect	157	232	158	233
rect	157	235	158	236
rect	157	238	158	239
rect	157	241	158	242
rect	157	244	158	245
rect	157	247	158	248
rect	157	250	158	251
rect	157	253	158	254
rect	157	256	158	257
rect	157	259	158	260
rect	157	262	158	263
rect	157	265	158	266
rect	157	268	158	269
rect	157	271	158	272
rect	157	274	158	275
rect	157	277	158	278
rect	157	280	158	281
rect	157	283	158	284
rect	157	286	158	287
rect	157	289	158	290
rect	157	292	158	293
rect	157	295	158	296
rect	157	298	158	299
rect	157	301	158	302
rect	157	307	158	308
rect	157	310	158	311
rect	157	313	158	314
rect	157	316	158	317
rect	157	319	158	320
rect	157	322	158	323
rect	157	325	158	326
rect	157	328	158	329
rect	157	331	158	332
rect	157	334	158	335
rect	157	337	158	338
rect	157	340	158	341
rect	157	343	158	344
rect	157	346	158	347
rect	157	349	158	350
rect	157	352	158	353
rect	157	355	158	356
rect	157	358	158	359
rect	157	361	158	362
rect	157	364	158	365
rect	157	367	158	368
rect	157	370	158	371
rect	157	373	158	374
rect	157	376	158	377
rect	157	379	158	380
rect	157	385	158	386
rect	158	1	159	2
rect	158	4	159	5
rect	158	7	159	8
rect	158	10	159	11
rect	158	13	159	14
rect	158	16	159	17
rect	158	19	159	20
rect	158	22	159	23
rect	158	25	159	26
rect	158	28	159	29
rect	158	31	159	32
rect	158	34	159	35
rect	158	37	159	38
rect	158	40	159	41
rect	158	43	159	44
rect	158	46	159	47
rect	158	49	159	50
rect	158	52	159	53
rect	158	55	159	56
rect	158	58	159	59
rect	158	61	159	62
rect	158	64	159	65
rect	158	67	159	68
rect	158	70	159	71
rect	158	73	159	74
rect	158	76	159	77
rect	158	79	159	80
rect	158	85	159	86
rect	158	88	159	89
rect	158	91	159	92
rect	158	94	159	95
rect	158	97	159	98
rect	158	100	159	101
rect	158	103	159	104
rect	158	106	159	107
rect	158	109	159	110
rect	158	112	159	113
rect	158	115	159	116
rect	158	118	159	119
rect	158	121	159	122
rect	158	124	159	125
rect	158	127	159	128
rect	158	130	159	131
rect	158	133	159	134
rect	158	136	159	137
rect	158	139	159	140
rect	158	142	159	143
rect	158	145	159	146
rect	158	148	159	149
rect	158	151	159	152
rect	158	154	159	155
rect	158	157	159	158
rect	158	160	159	161
rect	158	163	159	164
rect	158	166	159	167
rect	158	169	159	170
rect	158	172	159	173
rect	158	175	159	176
rect	158	178	159	179
rect	158	181	159	182
rect	158	184	159	185
rect	158	187	159	188
rect	158	190	159	191
rect	158	193	159	194
rect	158	196	159	197
rect	158	199	159	200
rect	158	202	159	203
rect	158	205	159	206
rect	158	208	159	209
rect	158	211	159	212
rect	158	214	159	215
rect	158	217	159	218
rect	158	220	159	221
rect	158	223	159	224
rect	158	226	159	227
rect	158	229	159	230
rect	158	232	159	233
rect	158	235	159	236
rect	158	238	159	239
rect	158	241	159	242
rect	158	244	159	245
rect	158	247	159	248
rect	158	250	159	251
rect	158	253	159	254
rect	158	256	159	257
rect	158	259	159	260
rect	158	262	159	263
rect	158	265	159	266
rect	158	268	159	269
rect	158	271	159	272
rect	158	274	159	275
rect	158	277	159	278
rect	158	283	159	284
rect	158	286	159	287
rect	158	289	159	290
rect	158	292	159	293
rect	158	295	159	296
rect	158	298	159	299
rect	158	301	159	302
rect	158	307	159	308
rect	158	310	159	311
rect	158	313	159	314
rect	158	316	159	317
rect	158	322	159	323
rect	158	325	159	326
rect	158	328	159	329
rect	158	331	159	332
rect	158	334	159	335
rect	158	337	159	338
rect	158	340	159	341
rect	158	343	159	344
rect	158	346	159	347
rect	158	349	159	350
rect	158	352	159	353
rect	158	355	159	356
rect	158	358	159	359
rect	158	361	159	362
rect	158	364	159	365
rect	158	367	159	368
rect	158	370	159	371
rect	158	373	159	374
rect	158	376	159	377
rect	158	379	159	380
rect	158	385	159	386
rect	159	1	160	2
rect	159	4	160	5
rect	159	7	160	8
rect	159	10	160	11
rect	159	13	160	14
rect	159	16	160	17
rect	159	19	160	20
rect	159	22	160	23
rect	159	25	160	26
rect	159	28	160	29
rect	159	31	160	32
rect	159	34	160	35
rect	159	37	160	38
rect	159	40	160	41
rect	159	43	160	44
rect	159	46	160	47
rect	159	49	160	50
rect	159	52	160	53
rect	159	55	160	56
rect	159	58	160	59
rect	159	61	160	62
rect	159	64	160	65
rect	159	67	160	68
rect	159	70	160	71
rect	159	73	160	74
rect	159	76	160	77
rect	159	79	160	80
rect	159	82	160	83
rect	159	85	160	86
rect	159	88	160	89
rect	159	91	160	92
rect	159	94	160	95
rect	159	97	160	98
rect	159	100	160	101
rect	159	103	160	104
rect	159	106	160	107
rect	159	109	160	110
rect	159	112	160	113
rect	159	115	160	116
rect	159	118	160	119
rect	159	121	160	122
rect	159	124	160	125
rect	159	127	160	128
rect	159	130	160	131
rect	159	133	160	134
rect	159	136	160	137
rect	159	139	160	140
rect	159	142	160	143
rect	159	145	160	146
rect	159	148	160	149
rect	159	151	160	152
rect	159	154	160	155
rect	159	157	160	158
rect	159	160	160	161
rect	159	163	160	164
rect	159	166	160	167
rect	159	169	160	170
rect	159	172	160	173
rect	159	175	160	176
rect	159	178	160	179
rect	159	181	160	182
rect	159	184	160	185
rect	159	187	160	188
rect	159	190	160	191
rect	159	193	160	194
rect	159	196	160	197
rect	159	199	160	200
rect	159	202	160	203
rect	159	205	160	206
rect	159	208	160	209
rect	159	211	160	212
rect	159	214	160	215
rect	159	217	160	218
rect	159	220	160	221
rect	159	223	160	224
rect	159	226	160	227
rect	159	229	160	230
rect	159	232	160	233
rect	159	235	160	236
rect	159	238	160	239
rect	159	241	160	242
rect	159	244	160	245
rect	159	247	160	248
rect	159	250	160	251
rect	159	253	160	254
rect	159	256	160	257
rect	159	259	160	260
rect	159	262	160	263
rect	159	265	160	266
rect	159	268	160	269
rect	159	271	160	272
rect	159	274	160	275
rect	159	277	160	278
rect	159	280	160	281
rect	159	283	160	284
rect	159	286	160	287
rect	159	289	160	290
rect	159	292	160	293
rect	159	295	160	296
rect	159	298	160	299
rect	159	301	160	302
rect	159	307	160	308
rect	159	310	160	311
rect	159	313	160	314
rect	159	316	160	317
rect	159	319	160	320
rect	159	322	160	323
rect	159	325	160	326
rect	159	328	160	329
rect	159	331	160	332
rect	159	334	160	335
rect	159	337	160	338
rect	159	340	160	341
rect	159	343	160	344
rect	159	346	160	347
rect	159	349	160	350
rect	159	352	160	353
rect	159	355	160	356
rect	159	358	160	359
rect	159	361	160	362
rect	159	364	160	365
rect	159	367	160	368
rect	159	370	160	371
rect	159	373	160	374
rect	159	376	160	377
rect	159	379	160	380
rect	159	385	160	386
rect	160	1	161	2
rect	160	4	161	5
rect	160	7	161	8
rect	160	10	161	11
rect	160	13	161	14
rect	160	16	161	17
rect	160	19	161	20
rect	160	22	161	23
rect	160	25	161	26
rect	160	28	161	29
rect	160	31	161	32
rect	160	34	161	35
rect	160	37	161	38
rect	160	40	161	41
rect	160	43	161	44
rect	160	46	161	47
rect	160	49	161	50
rect	160	52	161	53
rect	160	55	161	56
rect	160	58	161	59
rect	160	61	161	62
rect	160	64	161	65
rect	160	67	161	68
rect	160	70	161	71
rect	160	73	161	74
rect	160	76	161	77
rect	160	79	161	80
rect	160	82	161	83
rect	160	85	161	86
rect	160	88	161	89
rect	160	91	161	92
rect	160	94	161	95
rect	160	97	161	98
rect	160	100	161	101
rect	160	103	161	104
rect	160	106	161	107
rect	160	109	161	110
rect	160	112	161	113
rect	160	115	161	116
rect	160	118	161	119
rect	160	121	161	122
rect	160	124	161	125
rect	160	127	161	128
rect	160	130	161	131
rect	160	133	161	134
rect	160	136	161	137
rect	160	139	161	140
rect	160	142	161	143
rect	160	145	161	146
rect	160	148	161	149
rect	160	151	161	152
rect	160	154	161	155
rect	160	157	161	158
rect	160	160	161	161
rect	160	163	161	164
rect	160	166	161	167
rect	160	169	161	170
rect	160	172	161	173
rect	160	175	161	176
rect	160	178	161	179
rect	160	181	161	182
rect	160	184	161	185
rect	160	187	161	188
rect	160	190	161	191
rect	160	193	161	194
rect	160	196	161	197
rect	160	199	161	200
rect	160	202	161	203
rect	160	205	161	206
rect	160	208	161	209
rect	160	211	161	212
rect	160	214	161	215
rect	160	217	161	218
rect	160	220	161	221
rect	160	223	161	224
rect	160	226	161	227
rect	160	229	161	230
rect	160	232	161	233
rect	160	235	161	236
rect	160	238	161	239
rect	160	241	161	242
rect	160	244	161	245
rect	160	247	161	248
rect	160	250	161	251
rect	160	253	161	254
rect	160	256	161	257
rect	160	259	161	260
rect	160	262	161	263
rect	160	265	161	266
rect	160	268	161	269
rect	160	271	161	272
rect	160	274	161	275
rect	160	277	161	278
rect	160	280	161	281
rect	160	283	161	284
rect	160	286	161	287
rect	160	289	161	290
rect	160	292	161	293
rect	160	295	161	296
rect	160	298	161	299
rect	160	301	161	302
rect	160	307	161	308
rect	160	310	161	311
rect	160	313	161	314
rect	160	316	161	317
rect	160	319	161	320
rect	160	322	161	323
rect	160	325	161	326
rect	160	331	161	332
rect	160	334	161	335
rect	160	346	161	347
rect	160	349	161	350
rect	160	352	161	353
rect	160	355	161	356
rect	160	358	161	359
rect	160	361	161	362
rect	160	364	161	365
rect	160	367	161	368
rect	161	1	162	2
rect	161	4	162	5
rect	161	7	162	8
rect	161	10	162	11
rect	161	13	162	14
rect	161	16	162	17
rect	161	19	162	20
rect	161	22	162	23
rect	161	25	162	26
rect	161	28	162	29
rect	161	31	162	32
rect	161	34	162	35
rect	161	37	162	38
rect	161	40	162	41
rect	161	43	162	44
rect	161	46	162	47
rect	161	49	162	50
rect	161	52	162	53
rect	161	55	162	56
rect	161	58	162	59
rect	161	61	162	62
rect	161	64	162	65
rect	161	67	162	68
rect	161	70	162	71
rect	161	73	162	74
rect	161	76	162	77
rect	161	79	162	80
rect	161	82	162	83
rect	161	85	162	86
rect	161	88	162	89
rect	161	91	162	92
rect	161	94	162	95
rect	161	97	162	98
rect	161	100	162	101
rect	161	103	162	104
rect	161	106	162	107
rect	161	109	162	110
rect	161	112	162	113
rect	161	115	162	116
rect	161	118	162	119
rect	161	121	162	122
rect	161	124	162	125
rect	161	127	162	128
rect	161	130	162	131
rect	161	133	162	134
rect	161	136	162	137
rect	161	139	162	140
rect	161	142	162	143
rect	161	145	162	146
rect	161	148	162	149
rect	161	151	162	152
rect	161	154	162	155
rect	161	157	162	158
rect	161	160	162	161
rect	161	163	162	164
rect	161	166	162	167
rect	161	169	162	170
rect	161	172	162	173
rect	161	175	162	176
rect	161	178	162	179
rect	161	181	162	182
rect	161	184	162	185
rect	161	187	162	188
rect	161	190	162	191
rect	161	193	162	194
rect	161	196	162	197
rect	161	199	162	200
rect	161	202	162	203
rect	161	205	162	206
rect	161	208	162	209
rect	161	211	162	212
rect	161	214	162	215
rect	161	217	162	218
rect	161	220	162	221
rect	161	223	162	224
rect	161	226	162	227
rect	161	229	162	230
rect	161	232	162	233
rect	161	235	162	236
rect	161	238	162	239
rect	161	241	162	242
rect	161	244	162	245
rect	161	247	162	248
rect	161	250	162	251
rect	161	253	162	254
rect	161	256	162	257
rect	161	259	162	260
rect	161	262	162	263
rect	161	265	162	266
rect	161	268	162	269
rect	161	271	162	272
rect	161	274	162	275
rect	161	277	162	278
rect	161	280	162	281
rect	161	283	162	284
rect	161	286	162	287
rect	161	289	162	290
rect	161	292	162	293
rect	161	295	162	296
rect	161	298	162	299
rect	161	301	162	302
rect	161	307	162	308
rect	161	310	162	311
rect	161	313	162	314
rect	161	316	162	317
rect	161	319	162	320
rect	161	322	162	323
rect	161	325	162	326
rect	161	331	162	332
rect	161	334	162	335
rect	161	346	162	347
rect	161	349	162	350
rect	161	352	162	353
rect	161	355	162	356
rect	161	358	162	359
rect	161	361	162	362
rect	161	364	162	365
rect	161	367	162	368
rect	162	1	163	2
rect	162	4	163	5
rect	162	7	163	8
rect	162	10	163	11
rect	162	13	163	14
rect	162	16	163	17
rect	162	19	163	20
rect	162	22	163	23
rect	162	25	163	26
rect	162	28	163	29
rect	162	31	163	32
rect	162	34	163	35
rect	162	37	163	38
rect	162	40	163	41
rect	162	43	163	44
rect	162	46	163	47
rect	162	49	163	50
rect	162	52	163	53
rect	162	55	163	56
rect	162	58	163	59
rect	162	61	163	62
rect	162	64	163	65
rect	162	67	163	68
rect	162	70	163	71
rect	162	73	163	74
rect	162	76	163	77
rect	162	79	163	80
rect	162	82	163	83
rect	162	85	163	86
rect	162	88	163	89
rect	162	91	163	92
rect	162	94	163	95
rect	162	97	163	98
rect	162	100	163	101
rect	162	103	163	104
rect	162	106	163	107
rect	162	109	163	110
rect	162	112	163	113
rect	162	115	163	116
rect	162	118	163	119
rect	162	121	163	122
rect	162	124	163	125
rect	162	127	163	128
rect	162	130	163	131
rect	162	133	163	134
rect	162	136	163	137
rect	162	139	163	140
rect	162	142	163	143
rect	162	145	163	146
rect	162	148	163	149
rect	162	151	163	152
rect	162	154	163	155
rect	162	157	163	158
rect	162	160	163	161
rect	162	163	163	164
rect	162	166	163	167
rect	162	169	163	170
rect	162	172	163	173
rect	162	175	163	176
rect	162	178	163	179
rect	162	181	163	182
rect	162	184	163	185
rect	162	187	163	188
rect	162	190	163	191
rect	162	193	163	194
rect	162	196	163	197
rect	162	199	163	200
rect	162	202	163	203
rect	162	205	163	206
rect	162	208	163	209
rect	162	211	163	212
rect	162	214	163	215
rect	162	217	163	218
rect	162	220	163	221
rect	162	223	163	224
rect	162	226	163	227
rect	162	229	163	230
rect	162	232	163	233
rect	162	235	163	236
rect	162	238	163	239
rect	162	241	163	242
rect	162	244	163	245
rect	162	247	163	248
rect	162	250	163	251
rect	162	253	163	254
rect	162	256	163	257
rect	162	259	163	260
rect	162	262	163	263
rect	162	265	163	266
rect	162	268	163	269
rect	162	271	163	272
rect	162	274	163	275
rect	162	277	163	278
rect	162	280	163	281
rect	162	283	163	284
rect	162	286	163	287
rect	162	289	163	290
rect	162	292	163	293
rect	162	295	163	296
rect	162	298	163	299
rect	162	301	163	302
rect	162	307	163	308
rect	162	310	163	311
rect	162	313	163	314
rect	162	316	163	317
rect	162	319	163	320
rect	162	322	163	323
rect	162	325	163	326
rect	162	331	163	332
rect	162	334	163	335
rect	162	346	163	347
rect	162	349	163	350
rect	162	352	163	353
rect	162	355	163	356
rect	162	358	163	359
rect	162	361	163	362
rect	162	364	163	365
rect	162	367	163	368
rect	163	1	164	2
rect	163	4	164	5
rect	163	7	164	8
rect	163	10	164	11
rect	163	13	164	14
rect	163	16	164	17
rect	163	19	164	20
rect	163	22	164	23
rect	163	25	164	26
rect	163	28	164	29
rect	163	31	164	32
rect	163	34	164	35
rect	163	37	164	38
rect	163	40	164	41
rect	163	43	164	44
rect	163	46	164	47
rect	163	49	164	50
rect	163	52	164	53
rect	163	55	164	56
rect	163	58	164	59
rect	163	61	164	62
rect	163	64	164	65
rect	163	67	164	68
rect	163	70	164	71
rect	163	73	164	74
rect	163	76	164	77
rect	163	79	164	80
rect	163	82	164	83
rect	163	85	164	86
rect	163	88	164	89
rect	163	91	164	92
rect	163	94	164	95
rect	163	97	164	98
rect	163	100	164	101
rect	163	103	164	104
rect	163	106	164	107
rect	163	109	164	110
rect	163	112	164	113
rect	163	115	164	116
rect	163	118	164	119
rect	163	121	164	122
rect	163	124	164	125
rect	163	127	164	128
rect	163	130	164	131
rect	163	133	164	134
rect	163	136	164	137
rect	163	139	164	140
rect	163	142	164	143
rect	163	145	164	146
rect	163	148	164	149
rect	163	151	164	152
rect	163	154	164	155
rect	163	157	164	158
rect	163	160	164	161
rect	163	163	164	164
rect	163	166	164	167
rect	163	169	164	170
rect	163	172	164	173
rect	163	175	164	176
rect	163	178	164	179
rect	163	181	164	182
rect	163	184	164	185
rect	163	187	164	188
rect	163	190	164	191
rect	163	193	164	194
rect	163	196	164	197
rect	163	199	164	200
rect	163	202	164	203
rect	163	205	164	206
rect	163	208	164	209
rect	163	211	164	212
rect	163	214	164	215
rect	163	217	164	218
rect	163	220	164	221
rect	163	223	164	224
rect	163	226	164	227
rect	163	229	164	230
rect	163	232	164	233
rect	163	235	164	236
rect	163	238	164	239
rect	163	241	164	242
rect	163	244	164	245
rect	163	247	164	248
rect	163	250	164	251
rect	163	253	164	254
rect	163	256	164	257
rect	163	259	164	260
rect	163	262	164	263
rect	163	265	164	266
rect	163	268	164	269
rect	163	271	164	272
rect	163	274	164	275
rect	163	277	164	278
rect	163	280	164	281
rect	163	283	164	284
rect	163	286	164	287
rect	163	289	164	290
rect	163	292	164	293
rect	163	295	164	296
rect	163	298	164	299
rect	163	301	164	302
rect	163	307	164	308
rect	163	310	164	311
rect	163	313	164	314
rect	163	316	164	317
rect	163	319	164	320
rect	163	322	164	323
rect	163	325	164	326
rect	163	331	164	332
rect	163	334	164	335
rect	163	346	164	347
rect	163	349	164	350
rect	163	352	164	353
rect	163	355	164	356
rect	163	358	164	359
rect	163	361	164	362
rect	163	364	164	365
rect	163	367	164	368
rect	164	1	165	2
rect	164	4	165	5
rect	164	7	165	8
rect	164	10	165	11
rect	164	13	165	14
rect	164	16	165	17
rect	164	19	165	20
rect	164	22	165	23
rect	164	25	165	26
rect	164	28	165	29
rect	164	31	165	32
rect	164	34	165	35
rect	164	37	165	38
rect	164	40	165	41
rect	164	43	165	44
rect	164	46	165	47
rect	164	49	165	50
rect	164	52	165	53
rect	164	55	165	56
rect	164	58	165	59
rect	164	61	165	62
rect	164	64	165	65
rect	164	67	165	68
rect	164	70	165	71
rect	164	73	165	74
rect	164	76	165	77
rect	164	79	165	80
rect	164	82	165	83
rect	164	85	165	86
rect	164	88	165	89
rect	164	91	165	92
rect	164	94	165	95
rect	164	97	165	98
rect	164	100	165	101
rect	164	103	165	104
rect	164	106	165	107
rect	164	109	165	110
rect	164	112	165	113
rect	164	115	165	116
rect	164	118	165	119
rect	164	121	165	122
rect	164	124	165	125
rect	164	127	165	128
rect	164	130	165	131
rect	164	133	165	134
rect	164	136	165	137
rect	164	139	165	140
rect	164	142	165	143
rect	164	145	165	146
rect	164	148	165	149
rect	164	151	165	152
rect	164	154	165	155
rect	164	157	165	158
rect	164	160	165	161
rect	164	163	165	164
rect	164	166	165	167
rect	164	169	165	170
rect	164	172	165	173
rect	164	175	165	176
rect	164	178	165	179
rect	164	181	165	182
rect	164	184	165	185
rect	164	187	165	188
rect	164	190	165	191
rect	164	193	165	194
rect	164	196	165	197
rect	164	199	165	200
rect	164	202	165	203
rect	164	205	165	206
rect	164	208	165	209
rect	164	211	165	212
rect	164	214	165	215
rect	164	217	165	218
rect	164	220	165	221
rect	164	223	165	224
rect	164	226	165	227
rect	164	229	165	230
rect	164	232	165	233
rect	164	235	165	236
rect	164	238	165	239
rect	164	241	165	242
rect	164	244	165	245
rect	164	247	165	248
rect	164	250	165	251
rect	164	253	165	254
rect	164	256	165	257
rect	164	259	165	260
rect	164	262	165	263
rect	164	265	165	266
rect	164	268	165	269
rect	164	271	165	272
rect	164	274	165	275
rect	164	277	165	278
rect	164	280	165	281
rect	164	283	165	284
rect	164	286	165	287
rect	164	289	165	290
rect	164	292	165	293
rect	164	295	165	296
rect	164	298	165	299
rect	164	301	165	302
rect	164	307	165	308
rect	164	310	165	311
rect	164	313	165	314
rect	164	316	165	317
rect	164	319	165	320
rect	164	322	165	323
rect	164	325	165	326
rect	164	331	165	332
rect	164	334	165	335
rect	164	346	165	347
rect	164	349	165	350
rect	164	352	165	353
rect	164	355	165	356
rect	164	358	165	359
rect	164	361	165	362
rect	164	364	165	365
rect	164	367	165	368
rect	165	1	166	2
rect	165	4	166	5
rect	165	7	166	8
rect	165	10	166	11
rect	165	13	166	14
rect	165	16	166	17
rect	165	19	166	20
rect	165	22	166	23
rect	165	25	166	26
rect	165	28	166	29
rect	165	31	166	32
rect	165	34	166	35
rect	165	37	166	38
rect	165	40	166	41
rect	165	43	166	44
rect	165	46	166	47
rect	165	49	166	50
rect	165	52	166	53
rect	165	55	166	56
rect	165	58	166	59
rect	165	61	166	62
rect	165	64	166	65
rect	165	67	166	68
rect	165	70	166	71
rect	165	73	166	74
rect	165	76	166	77
rect	165	79	166	80
rect	165	82	166	83
rect	165	85	166	86
rect	165	88	166	89
rect	165	91	166	92
rect	165	94	166	95
rect	165	97	166	98
rect	165	100	166	101
rect	165	103	166	104
rect	165	106	166	107
rect	165	109	166	110
rect	165	112	166	113
rect	165	115	166	116
rect	165	118	166	119
rect	165	121	166	122
rect	165	124	166	125
rect	165	127	166	128
rect	165	130	166	131
rect	165	133	166	134
rect	165	136	166	137
rect	165	139	166	140
rect	165	142	166	143
rect	165	145	166	146
rect	165	148	166	149
rect	165	151	166	152
rect	165	154	166	155
rect	165	157	166	158
rect	165	160	166	161
rect	165	163	166	164
rect	165	166	166	167
rect	165	169	166	170
rect	165	172	166	173
rect	165	175	166	176
rect	165	178	166	179
rect	165	181	166	182
rect	165	184	166	185
rect	165	187	166	188
rect	165	190	166	191
rect	165	193	166	194
rect	165	196	166	197
rect	165	199	166	200
rect	165	202	166	203
rect	165	205	166	206
rect	165	208	166	209
rect	165	211	166	212
rect	165	214	166	215
rect	165	217	166	218
rect	165	220	166	221
rect	165	223	166	224
rect	165	226	166	227
rect	165	229	166	230
rect	165	232	166	233
rect	165	235	166	236
rect	165	238	166	239
rect	165	241	166	242
rect	165	244	166	245
rect	165	247	166	248
rect	165	250	166	251
rect	165	253	166	254
rect	165	256	166	257
rect	165	259	166	260
rect	165	262	166	263
rect	165	265	166	266
rect	165	268	166	269
rect	165	271	166	272
rect	165	274	166	275
rect	165	277	166	278
rect	165	280	166	281
rect	165	283	166	284
rect	165	286	166	287
rect	165	289	166	290
rect	165	292	166	293
rect	165	295	166	296
rect	165	298	166	299
rect	165	301	166	302
rect	165	307	166	308
rect	165	310	166	311
rect	165	313	166	314
rect	165	316	166	317
rect	165	319	166	320
rect	165	322	166	323
rect	165	325	166	326
rect	165	331	166	332
rect	165	334	166	335
rect	165	346	166	347
rect	165	349	166	350
rect	165	352	166	353
rect	165	355	166	356
rect	165	358	166	359
rect	165	361	166	362
rect	165	364	166	365
rect	165	367	166	368
rect	166	1	167	2
rect	166	4	167	5
rect	166	7	167	8
rect	166	10	167	11
rect	166	13	167	14
rect	166	16	167	17
rect	166	19	167	20
rect	166	22	167	23
rect	166	25	167	26
rect	166	28	167	29
rect	166	31	167	32
rect	166	34	167	35
rect	166	37	167	38
rect	166	40	167	41
rect	166	43	167	44
rect	166	46	167	47
rect	166	49	167	50
rect	166	52	167	53
rect	166	55	167	56
rect	166	58	167	59
rect	166	61	167	62
rect	166	64	167	65
rect	166	67	167	68
rect	166	70	167	71
rect	166	73	167	74
rect	166	76	167	77
rect	166	79	167	80
rect	166	82	167	83
rect	166	85	167	86
rect	166	88	167	89
rect	166	91	167	92
rect	166	94	167	95
rect	166	97	167	98
rect	166	100	167	101
rect	166	103	167	104
rect	166	106	167	107
rect	166	109	167	110
rect	166	112	167	113
rect	166	115	167	116
rect	166	118	167	119
rect	166	121	167	122
rect	166	124	167	125
rect	166	127	167	128
rect	166	130	167	131
rect	166	133	167	134
rect	166	136	167	137
rect	166	139	167	140
rect	166	142	167	143
rect	166	145	167	146
rect	166	148	167	149
rect	166	151	167	152
rect	166	154	167	155
rect	166	157	167	158
rect	166	160	167	161
rect	166	163	167	164
rect	166	166	167	167
rect	166	169	167	170
rect	166	172	167	173
rect	166	175	167	176
rect	166	178	167	179
rect	166	181	167	182
rect	166	184	167	185
rect	166	187	167	188
rect	166	190	167	191
rect	166	193	167	194
rect	166	196	167	197
rect	166	199	167	200
rect	166	202	167	203
rect	166	205	167	206
rect	166	208	167	209
rect	166	211	167	212
rect	166	214	167	215
rect	166	217	167	218
rect	166	220	167	221
rect	166	223	167	224
rect	166	226	167	227
rect	166	229	167	230
rect	166	232	167	233
rect	166	235	167	236
rect	166	238	167	239
rect	166	241	167	242
rect	166	244	167	245
rect	166	247	167	248
rect	166	250	167	251
rect	166	253	167	254
rect	166	256	167	257
rect	166	259	167	260
rect	166	262	167	263
rect	166	265	167	266
rect	166	268	167	269
rect	166	271	167	272
rect	166	274	167	275
rect	166	277	167	278
rect	166	280	167	281
rect	166	283	167	284
rect	166	286	167	287
rect	166	289	167	290
rect	166	292	167	293
rect	166	295	167	296
rect	166	298	167	299
rect	166	301	167	302
rect	166	307	167	308
rect	166	310	167	311
rect	166	313	167	314
rect	166	316	167	317
rect	166	319	167	320
rect	166	322	167	323
rect	166	325	167	326
rect	166	331	167	332
rect	166	334	167	335
rect	166	346	167	347
rect	166	349	167	350
rect	166	352	167	353
rect	166	355	167	356
rect	166	358	167	359
rect	166	361	167	362
rect	166	364	167	365
rect	166	367	167	368
rect	167	1	168	2
rect	167	4	168	5
rect	167	7	168	8
rect	167	10	168	11
rect	167	13	168	14
rect	167	16	168	17
rect	167	19	168	20
rect	167	22	168	23
rect	167	25	168	26
rect	167	28	168	29
rect	167	31	168	32
rect	167	34	168	35
rect	167	37	168	38
rect	167	40	168	41
rect	167	43	168	44
rect	167	49	168	50
rect	167	52	168	53
rect	167	55	168	56
rect	167	58	168	59
rect	167	61	168	62
rect	167	64	168	65
rect	167	67	168	68
rect	167	70	168	71
rect	167	73	168	74
rect	167	76	168	77
rect	167	79	168	80
rect	167	82	168	83
rect	167	85	168	86
rect	167	88	168	89
rect	167	91	168	92
rect	167	94	168	95
rect	167	97	168	98
rect	167	100	168	101
rect	167	103	168	104
rect	167	106	168	107
rect	167	109	168	110
rect	167	112	168	113
rect	167	115	168	116
rect	167	118	168	119
rect	167	121	168	122
rect	167	124	168	125
rect	167	127	168	128
rect	167	130	168	131
rect	167	133	168	134
rect	167	136	168	137
rect	167	139	168	140
rect	167	142	168	143
rect	167	145	168	146
rect	167	148	168	149
rect	167	151	168	152
rect	167	154	168	155
rect	167	157	168	158
rect	167	160	168	161
rect	167	163	168	164
rect	167	166	168	167
rect	167	169	168	170
rect	167	172	168	173
rect	167	175	168	176
rect	167	178	168	179
rect	167	181	168	182
rect	167	184	168	185
rect	167	187	168	188
rect	167	190	168	191
rect	167	193	168	194
rect	167	196	168	197
rect	167	199	168	200
rect	167	202	168	203
rect	167	205	168	206
rect	167	208	168	209
rect	167	211	168	212
rect	167	214	168	215
rect	167	217	168	218
rect	167	220	168	221
rect	167	223	168	224
rect	167	226	168	227
rect	167	229	168	230
rect	167	232	168	233
rect	167	235	168	236
rect	167	238	168	239
rect	167	241	168	242
rect	167	244	168	245
rect	167	247	168	248
rect	167	250	168	251
rect	167	253	168	254
rect	167	256	168	257
rect	167	259	168	260
rect	167	262	168	263
rect	167	265	168	266
rect	167	268	168	269
rect	167	271	168	272
rect	167	274	168	275
rect	167	277	168	278
rect	167	280	168	281
rect	167	283	168	284
rect	167	286	168	287
rect	167	289	168	290
rect	167	292	168	293
rect	167	295	168	296
rect	167	298	168	299
rect	167	301	168	302
rect	167	307	168	308
rect	167	310	168	311
rect	167	313	168	314
rect	167	316	168	317
rect	167	319	168	320
rect	167	322	168	323
rect	167	325	168	326
rect	167	331	168	332
rect	167	334	168	335
rect	167	346	168	347
rect	167	349	168	350
rect	167	352	168	353
rect	167	355	168	356
rect	167	361	168	362
rect	167	364	168	365
rect	167	367	168	368
rect	168	1	169	2
rect	168	4	169	5
rect	168	7	169	8
rect	168	10	169	11
rect	168	13	169	14
rect	168	16	169	17
rect	168	19	169	20
rect	168	22	169	23
rect	168	25	169	26
rect	168	28	169	29
rect	168	31	169	32
rect	168	34	169	35
rect	168	37	169	38
rect	168	40	169	41
rect	168	43	169	44
rect	168	46	169	47
rect	168	49	169	50
rect	168	52	169	53
rect	168	55	169	56
rect	168	58	169	59
rect	168	61	169	62
rect	168	64	169	65
rect	168	67	169	68
rect	168	70	169	71
rect	168	73	169	74
rect	168	76	169	77
rect	168	79	169	80
rect	168	82	169	83
rect	168	85	169	86
rect	168	88	169	89
rect	168	91	169	92
rect	168	94	169	95
rect	168	97	169	98
rect	168	100	169	101
rect	168	103	169	104
rect	168	106	169	107
rect	168	109	169	110
rect	168	112	169	113
rect	168	115	169	116
rect	168	118	169	119
rect	168	121	169	122
rect	168	124	169	125
rect	168	127	169	128
rect	168	130	169	131
rect	168	133	169	134
rect	168	136	169	137
rect	168	139	169	140
rect	168	142	169	143
rect	168	145	169	146
rect	168	148	169	149
rect	168	151	169	152
rect	168	154	169	155
rect	168	157	169	158
rect	168	160	169	161
rect	168	163	169	164
rect	168	166	169	167
rect	168	169	169	170
rect	168	172	169	173
rect	168	175	169	176
rect	168	178	169	179
rect	168	181	169	182
rect	168	184	169	185
rect	168	187	169	188
rect	168	190	169	191
rect	168	193	169	194
rect	168	196	169	197
rect	168	199	169	200
rect	168	202	169	203
rect	168	205	169	206
rect	168	208	169	209
rect	168	211	169	212
rect	168	214	169	215
rect	168	217	169	218
rect	168	220	169	221
rect	168	223	169	224
rect	168	226	169	227
rect	168	229	169	230
rect	168	232	169	233
rect	168	235	169	236
rect	168	238	169	239
rect	168	241	169	242
rect	168	244	169	245
rect	168	247	169	248
rect	168	250	169	251
rect	168	253	169	254
rect	168	256	169	257
rect	168	259	169	260
rect	168	262	169	263
rect	168	265	169	266
rect	168	268	169	269
rect	168	271	169	272
rect	168	274	169	275
rect	168	277	169	278
rect	168	280	169	281
rect	168	283	169	284
rect	168	286	169	287
rect	168	289	169	290
rect	168	292	169	293
rect	168	295	169	296
rect	168	298	169	299
rect	168	301	169	302
rect	168	307	169	308
rect	168	310	169	311
rect	168	313	169	314
rect	168	316	169	317
rect	168	319	169	320
rect	168	322	169	323
rect	168	325	169	326
rect	168	331	169	332
rect	168	334	169	335
rect	168	346	169	347
rect	168	349	169	350
rect	168	352	169	353
rect	168	355	169	356
rect	168	358	169	359
rect	168	361	169	362
rect	168	364	169	365
rect	168	367	169	368
rect	169	1	170	2
rect	169	4	170	5
rect	169	7	170	8
rect	169	10	170	11
rect	169	13	170	14
rect	169	16	170	17
rect	169	19	170	20
rect	169	22	170	23
rect	169	25	170	26
rect	169	28	170	29
rect	169	31	170	32
rect	169	34	170	35
rect	169	37	170	38
rect	169	40	170	41
rect	169	43	170	44
rect	169	46	170	47
rect	169	49	170	50
rect	169	52	170	53
rect	169	55	170	56
rect	169	58	170	59
rect	169	61	170	62
rect	169	64	170	65
rect	169	67	170	68
rect	169	70	170	71
rect	169	73	170	74
rect	169	76	170	77
rect	169	79	170	80
rect	169	82	170	83
rect	169	85	170	86
rect	169	88	170	89
rect	169	91	170	92
rect	169	94	170	95
rect	169	97	170	98
rect	169	100	170	101
rect	169	103	170	104
rect	169	106	170	107
rect	169	109	170	110
rect	169	112	170	113
rect	169	115	170	116
rect	169	118	170	119
rect	169	121	170	122
rect	169	124	170	125
rect	169	127	170	128
rect	169	130	170	131
rect	169	133	170	134
rect	169	136	170	137
rect	169	139	170	140
rect	169	142	170	143
rect	169	145	170	146
rect	169	148	170	149
rect	169	151	170	152
rect	169	154	170	155
rect	169	157	170	158
rect	169	160	170	161
rect	169	163	170	164
rect	169	166	170	167
rect	169	169	170	170
rect	169	172	170	173
rect	169	175	170	176
rect	169	178	170	179
rect	169	181	170	182
rect	169	184	170	185
rect	169	187	170	188
rect	169	190	170	191
rect	169	193	170	194
rect	169	196	170	197
rect	169	199	170	200
rect	169	202	170	203
rect	169	205	170	206
rect	169	208	170	209
rect	169	211	170	212
rect	169	214	170	215
rect	169	217	170	218
rect	169	220	170	221
rect	169	223	170	224
rect	169	226	170	227
rect	169	229	170	230
rect	169	232	170	233
rect	169	235	170	236
rect	169	238	170	239
rect	169	241	170	242
rect	169	244	170	245
rect	169	247	170	248
rect	169	250	170	251
rect	169	253	170	254
rect	169	256	170	257
rect	169	259	170	260
rect	169	262	170	263
rect	169	265	170	266
rect	169	268	170	269
rect	169	271	170	272
rect	169	274	170	275
rect	169	277	170	278
rect	169	280	170	281
rect	169	283	170	284
rect	169	286	170	287
rect	169	289	170	290
rect	169	292	170	293
rect	169	295	170	296
rect	169	298	170	299
rect	169	301	170	302
rect	169	307	170	308
rect	169	310	170	311
rect	169	313	170	314
rect	169	316	170	317
rect	169	319	170	320
rect	169	322	170	323
rect	169	325	170	326
rect	169	331	170	332
rect	169	334	170	335
rect	169	346	170	347
rect	169	349	170	350
rect	169	352	170	353
rect	169	355	170	356
rect	169	358	170	359
rect	169	361	170	362
rect	169	364	170	365
rect	169	367	170	368
rect	170	1	171	2
rect	170	4	171	5
rect	170	7	171	8
rect	170	10	171	11
rect	170	13	171	14
rect	170	16	171	17
rect	170	19	171	20
rect	170	22	171	23
rect	170	25	171	26
rect	170	28	171	29
rect	170	31	171	32
rect	170	34	171	35
rect	170	37	171	38
rect	170	40	171	41
rect	170	43	171	44
rect	170	46	171	47
rect	170	49	171	50
rect	170	52	171	53
rect	170	55	171	56
rect	170	58	171	59
rect	170	61	171	62
rect	170	64	171	65
rect	170	67	171	68
rect	170	70	171	71
rect	170	73	171	74
rect	170	76	171	77
rect	170	79	171	80
rect	170	82	171	83
rect	170	85	171	86
rect	170	88	171	89
rect	170	91	171	92
rect	170	94	171	95
rect	170	97	171	98
rect	170	100	171	101
rect	170	103	171	104
rect	170	106	171	107
rect	170	109	171	110
rect	170	112	171	113
rect	170	115	171	116
rect	170	118	171	119
rect	170	121	171	122
rect	170	124	171	125
rect	170	127	171	128
rect	170	130	171	131
rect	170	133	171	134
rect	170	136	171	137
rect	170	139	171	140
rect	170	142	171	143
rect	170	145	171	146
rect	170	148	171	149
rect	170	151	171	152
rect	170	154	171	155
rect	170	157	171	158
rect	170	160	171	161
rect	170	163	171	164
rect	170	166	171	167
rect	170	169	171	170
rect	170	172	171	173
rect	170	175	171	176
rect	170	178	171	179
rect	170	181	171	182
rect	170	184	171	185
rect	170	187	171	188
rect	170	190	171	191
rect	170	193	171	194
rect	170	196	171	197
rect	170	199	171	200
rect	170	202	171	203
rect	170	205	171	206
rect	170	208	171	209
rect	170	211	171	212
rect	170	214	171	215
rect	170	217	171	218
rect	170	220	171	221
rect	170	223	171	224
rect	170	226	171	227
rect	170	229	171	230
rect	170	232	171	233
rect	170	235	171	236
rect	170	238	171	239
rect	170	241	171	242
rect	170	244	171	245
rect	170	247	171	248
rect	170	250	171	251
rect	170	253	171	254
rect	170	256	171	257
rect	170	259	171	260
rect	170	262	171	263
rect	170	265	171	266
rect	170	268	171	269
rect	170	271	171	272
rect	170	274	171	275
rect	170	277	171	278
rect	170	280	171	281
rect	170	283	171	284
rect	170	286	171	287
rect	170	289	171	290
rect	170	292	171	293
rect	170	295	171	296
rect	170	298	171	299
rect	170	301	171	302
rect	170	307	171	308
rect	170	310	171	311
rect	170	313	171	314
rect	170	316	171	317
rect	170	319	171	320
rect	170	322	171	323
rect	170	325	171	326
rect	170	331	171	332
rect	170	334	171	335
rect	170	346	171	347
rect	170	349	171	350
rect	170	352	171	353
rect	170	355	171	356
rect	170	358	171	359
rect	170	361	171	362
rect	170	364	171	365
rect	170	367	171	368
rect	171	1	172	2
rect	171	7	172	8
rect	171	10	172	11
rect	171	13	172	14
rect	171	16	172	17
rect	171	19	172	20
rect	171	22	172	23
rect	171	25	172	26
rect	171	28	172	29
rect	171	31	172	32
rect	171	34	172	35
rect	171	37	172	38
rect	171	40	172	41
rect	171	43	172	44
rect	171	46	172	47
rect	171	49	172	50
rect	171	52	172	53
rect	171	55	172	56
rect	171	58	172	59
rect	171	61	172	62
rect	171	64	172	65
rect	171	67	172	68
rect	171	70	172	71
rect	171	73	172	74
rect	171	76	172	77
rect	171	79	172	80
rect	171	82	172	83
rect	171	85	172	86
rect	171	88	172	89
rect	171	91	172	92
rect	171	94	172	95
rect	171	97	172	98
rect	171	100	172	101
rect	171	103	172	104
rect	171	106	172	107
rect	171	109	172	110
rect	171	112	172	113
rect	171	115	172	116
rect	171	118	172	119
rect	171	121	172	122
rect	171	124	172	125
rect	171	127	172	128
rect	171	130	172	131
rect	171	133	172	134
rect	171	136	172	137
rect	171	139	172	140
rect	171	142	172	143
rect	171	145	172	146
rect	171	148	172	149
rect	171	151	172	152
rect	171	154	172	155
rect	171	157	172	158
rect	171	160	172	161
rect	171	163	172	164
rect	171	166	172	167
rect	171	169	172	170
rect	171	172	172	173
rect	171	175	172	176
rect	171	178	172	179
rect	171	181	172	182
rect	171	184	172	185
rect	171	187	172	188
rect	171	190	172	191
rect	171	193	172	194
rect	171	196	172	197
rect	171	199	172	200
rect	171	202	172	203
rect	171	205	172	206
rect	171	208	172	209
rect	171	211	172	212
rect	171	214	172	215
rect	171	217	172	218
rect	171	220	172	221
rect	171	223	172	224
rect	171	226	172	227
rect	171	229	172	230
rect	171	232	172	233
rect	171	235	172	236
rect	171	238	172	239
rect	171	241	172	242
rect	171	244	172	245
rect	171	247	172	248
rect	171	250	172	251
rect	171	253	172	254
rect	171	256	172	257
rect	171	259	172	260
rect	171	262	172	263
rect	171	265	172	266
rect	171	268	172	269
rect	171	271	172	272
rect	171	274	172	275
rect	171	277	172	278
rect	171	280	172	281
rect	171	283	172	284
rect	171	286	172	287
rect	171	289	172	290
rect	171	292	172	293
rect	171	295	172	296
rect	171	298	172	299
rect	171	301	172	302
rect	171	307	172	308
rect	171	310	172	311
rect	171	313	172	314
rect	171	316	172	317
rect	171	322	172	323
rect	171	325	172	326
rect	171	331	172	332
rect	171	334	172	335
rect	171	346	172	347
rect	171	349	172	350
rect	171	352	172	353
rect	171	355	172	356
rect	171	358	172	359
rect	171	361	172	362
rect	171	364	172	365
rect	171	367	172	368
rect	172	1	173	2
rect	172	4	173	5
rect	172	7	173	8
rect	172	10	173	11
rect	172	13	173	14
rect	172	16	173	17
rect	172	19	173	20
rect	172	22	173	23
rect	172	25	173	26
rect	172	28	173	29
rect	172	31	173	32
rect	172	34	173	35
rect	172	37	173	38
rect	172	40	173	41
rect	172	43	173	44
rect	172	46	173	47
rect	172	49	173	50
rect	172	52	173	53
rect	172	55	173	56
rect	172	58	173	59
rect	172	61	173	62
rect	172	64	173	65
rect	172	67	173	68
rect	172	70	173	71
rect	172	73	173	74
rect	172	76	173	77
rect	172	79	173	80
rect	172	82	173	83
rect	172	85	173	86
rect	172	88	173	89
rect	172	91	173	92
rect	172	94	173	95
rect	172	97	173	98
rect	172	100	173	101
rect	172	103	173	104
rect	172	106	173	107
rect	172	109	173	110
rect	172	112	173	113
rect	172	115	173	116
rect	172	118	173	119
rect	172	121	173	122
rect	172	124	173	125
rect	172	127	173	128
rect	172	130	173	131
rect	172	133	173	134
rect	172	136	173	137
rect	172	139	173	140
rect	172	142	173	143
rect	172	145	173	146
rect	172	148	173	149
rect	172	151	173	152
rect	172	154	173	155
rect	172	157	173	158
rect	172	160	173	161
rect	172	163	173	164
rect	172	166	173	167
rect	172	169	173	170
rect	172	172	173	173
rect	172	175	173	176
rect	172	178	173	179
rect	172	181	173	182
rect	172	184	173	185
rect	172	187	173	188
rect	172	190	173	191
rect	172	193	173	194
rect	172	196	173	197
rect	172	199	173	200
rect	172	202	173	203
rect	172	205	173	206
rect	172	208	173	209
rect	172	211	173	212
rect	172	214	173	215
rect	172	217	173	218
rect	172	220	173	221
rect	172	223	173	224
rect	172	226	173	227
rect	172	229	173	230
rect	172	232	173	233
rect	172	235	173	236
rect	172	238	173	239
rect	172	241	173	242
rect	172	244	173	245
rect	172	247	173	248
rect	172	250	173	251
rect	172	253	173	254
rect	172	256	173	257
rect	172	259	173	260
rect	172	262	173	263
rect	172	265	173	266
rect	172	268	173	269
rect	172	271	173	272
rect	172	274	173	275
rect	172	277	173	278
rect	172	280	173	281
rect	172	283	173	284
rect	172	286	173	287
rect	172	289	173	290
rect	172	292	173	293
rect	172	295	173	296
rect	172	298	173	299
rect	172	301	173	302
rect	172	307	173	308
rect	172	310	173	311
rect	172	313	173	314
rect	172	316	173	317
rect	172	319	173	320
rect	172	322	173	323
rect	172	325	173	326
rect	172	331	173	332
rect	172	334	173	335
rect	172	346	173	347
rect	172	349	173	350
rect	172	352	173	353
rect	172	355	173	356
rect	172	358	173	359
rect	172	361	173	362
rect	172	364	173	365
rect	172	367	173	368
rect	173	1	174	2
rect	173	4	174	5
rect	173	7	174	8
rect	173	10	174	11
rect	173	13	174	14
rect	173	16	174	17
rect	173	19	174	20
rect	173	22	174	23
rect	173	25	174	26
rect	173	28	174	29
rect	173	31	174	32
rect	173	34	174	35
rect	173	37	174	38
rect	173	40	174	41
rect	173	43	174	44
rect	173	46	174	47
rect	173	49	174	50
rect	173	52	174	53
rect	173	55	174	56
rect	173	58	174	59
rect	173	61	174	62
rect	173	64	174	65
rect	173	67	174	68
rect	173	70	174	71
rect	173	73	174	74
rect	173	76	174	77
rect	173	79	174	80
rect	173	82	174	83
rect	173	85	174	86
rect	173	88	174	89
rect	173	91	174	92
rect	173	94	174	95
rect	173	97	174	98
rect	173	100	174	101
rect	173	103	174	104
rect	173	106	174	107
rect	173	109	174	110
rect	173	112	174	113
rect	173	115	174	116
rect	173	118	174	119
rect	173	121	174	122
rect	173	124	174	125
rect	173	127	174	128
rect	173	130	174	131
rect	173	133	174	134
rect	173	136	174	137
rect	173	139	174	140
rect	173	142	174	143
rect	173	145	174	146
rect	173	148	174	149
rect	173	151	174	152
rect	173	154	174	155
rect	173	157	174	158
rect	173	160	174	161
rect	173	163	174	164
rect	173	166	174	167
rect	173	169	174	170
rect	173	172	174	173
rect	173	175	174	176
rect	173	178	174	179
rect	173	181	174	182
rect	173	184	174	185
rect	173	187	174	188
rect	173	190	174	191
rect	173	193	174	194
rect	173	196	174	197
rect	173	199	174	200
rect	173	202	174	203
rect	173	205	174	206
rect	173	208	174	209
rect	173	211	174	212
rect	173	214	174	215
rect	173	217	174	218
rect	173	220	174	221
rect	173	223	174	224
rect	173	226	174	227
rect	173	229	174	230
rect	173	232	174	233
rect	173	235	174	236
rect	173	238	174	239
rect	173	241	174	242
rect	173	244	174	245
rect	173	247	174	248
rect	173	250	174	251
rect	173	253	174	254
rect	173	256	174	257
rect	173	259	174	260
rect	173	262	174	263
rect	173	265	174	266
rect	173	268	174	269
rect	173	271	174	272
rect	173	274	174	275
rect	173	277	174	278
rect	173	280	174	281
rect	173	283	174	284
rect	173	286	174	287
rect	173	289	174	290
rect	173	292	174	293
rect	173	295	174	296
rect	173	298	174	299
rect	173	301	174	302
rect	173	307	174	308
rect	173	310	174	311
rect	173	313	174	314
rect	173	316	174	317
rect	173	322	174	323
rect	173	325	174	326
rect	173	331	174	332
rect	173	334	174	335
rect	173	346	174	347
rect	173	349	174	350
rect	173	355	174	356
rect	173	361	174	362
rect	173	364	174	365
rect	173	367	174	368
rect	174	1	175	2
rect	174	4	175	5
rect	174	7	175	8
rect	174	10	175	11
rect	174	13	175	14
rect	174	16	175	17
rect	174	19	175	20
rect	174	22	175	23
rect	174	25	175	26
rect	174	28	175	29
rect	174	31	175	32
rect	174	34	175	35
rect	174	37	175	38
rect	174	40	175	41
rect	174	43	175	44
rect	174	46	175	47
rect	174	49	175	50
rect	174	52	175	53
rect	174	55	175	56
rect	174	58	175	59
rect	174	61	175	62
rect	174	64	175	65
rect	174	67	175	68
rect	174	70	175	71
rect	174	73	175	74
rect	174	76	175	77
rect	174	79	175	80
rect	174	82	175	83
rect	174	85	175	86
rect	174	88	175	89
rect	174	91	175	92
rect	174	94	175	95
rect	174	97	175	98
rect	174	100	175	101
rect	174	103	175	104
rect	174	106	175	107
rect	174	109	175	110
rect	174	112	175	113
rect	174	115	175	116
rect	174	118	175	119
rect	174	121	175	122
rect	174	124	175	125
rect	174	127	175	128
rect	174	130	175	131
rect	174	133	175	134
rect	174	136	175	137
rect	174	139	175	140
rect	174	142	175	143
rect	174	145	175	146
rect	174	148	175	149
rect	174	151	175	152
rect	174	154	175	155
rect	174	157	175	158
rect	174	160	175	161
rect	174	163	175	164
rect	174	166	175	167
rect	174	169	175	170
rect	174	172	175	173
rect	174	175	175	176
rect	174	178	175	179
rect	174	181	175	182
rect	174	184	175	185
rect	174	187	175	188
rect	174	190	175	191
rect	174	193	175	194
rect	174	196	175	197
rect	174	199	175	200
rect	174	202	175	203
rect	174	205	175	206
rect	174	208	175	209
rect	174	211	175	212
rect	174	214	175	215
rect	174	217	175	218
rect	174	220	175	221
rect	174	223	175	224
rect	174	226	175	227
rect	174	229	175	230
rect	174	232	175	233
rect	174	235	175	236
rect	174	238	175	239
rect	174	241	175	242
rect	174	244	175	245
rect	174	247	175	248
rect	174	250	175	251
rect	174	253	175	254
rect	174	256	175	257
rect	174	259	175	260
rect	174	262	175	263
rect	174	265	175	266
rect	174	268	175	269
rect	174	271	175	272
rect	174	274	175	275
rect	174	277	175	278
rect	174	280	175	281
rect	174	283	175	284
rect	174	286	175	287
rect	174	289	175	290
rect	174	292	175	293
rect	174	295	175	296
rect	174	298	175	299
rect	174	301	175	302
rect	174	307	175	308
rect	174	310	175	311
rect	174	313	175	314
rect	174	316	175	317
rect	174	322	175	323
rect	174	325	175	326
rect	174	331	175	332
rect	174	334	175	335
rect	174	346	175	347
rect	174	349	175	350
rect	174	355	175	356
rect	174	361	175	362
rect	174	364	175	365
rect	174	367	175	368
rect	175	1	176	2
rect	175	4	176	5
rect	175	7	176	8
rect	175	10	176	11
rect	175	13	176	14
rect	175	16	176	17
rect	175	19	176	20
rect	175	22	176	23
rect	175	25	176	26
rect	175	28	176	29
rect	175	31	176	32
rect	175	34	176	35
rect	175	37	176	38
rect	175	40	176	41
rect	175	43	176	44
rect	175	46	176	47
rect	175	49	176	50
rect	175	52	176	53
rect	175	55	176	56
rect	175	58	176	59
rect	175	61	176	62
rect	175	64	176	65
rect	175	67	176	68
rect	175	70	176	71
rect	175	73	176	74
rect	175	76	176	77
rect	175	79	176	80
rect	175	82	176	83
rect	175	85	176	86
rect	175	88	176	89
rect	175	91	176	92
rect	175	94	176	95
rect	175	97	176	98
rect	175	100	176	101
rect	175	103	176	104
rect	175	106	176	107
rect	175	109	176	110
rect	175	112	176	113
rect	175	115	176	116
rect	175	118	176	119
rect	175	121	176	122
rect	175	124	176	125
rect	175	127	176	128
rect	175	130	176	131
rect	175	133	176	134
rect	175	136	176	137
rect	175	139	176	140
rect	175	142	176	143
rect	175	145	176	146
rect	175	148	176	149
rect	175	151	176	152
rect	175	154	176	155
rect	175	157	176	158
rect	175	160	176	161
rect	175	163	176	164
rect	175	166	176	167
rect	175	169	176	170
rect	175	172	176	173
rect	175	175	176	176
rect	175	178	176	179
rect	175	181	176	182
rect	175	184	176	185
rect	175	187	176	188
rect	175	190	176	191
rect	175	193	176	194
rect	175	196	176	197
rect	175	199	176	200
rect	175	202	176	203
rect	175	205	176	206
rect	175	208	176	209
rect	175	211	176	212
rect	175	214	176	215
rect	175	217	176	218
rect	175	220	176	221
rect	175	223	176	224
rect	175	226	176	227
rect	175	229	176	230
rect	175	232	176	233
rect	175	235	176	236
rect	175	238	176	239
rect	175	241	176	242
rect	175	244	176	245
rect	175	247	176	248
rect	175	250	176	251
rect	175	253	176	254
rect	175	256	176	257
rect	175	259	176	260
rect	175	262	176	263
rect	175	265	176	266
rect	175	268	176	269
rect	175	271	176	272
rect	175	274	176	275
rect	175	277	176	278
rect	175	280	176	281
rect	175	283	176	284
rect	175	286	176	287
rect	175	289	176	290
rect	175	292	176	293
rect	175	295	176	296
rect	175	298	176	299
rect	175	301	176	302
rect	175	307	176	308
rect	175	310	176	311
rect	175	313	176	314
rect	175	316	176	317
rect	175	322	176	323
rect	175	325	176	326
rect	175	331	176	332
rect	175	334	176	335
rect	175	346	176	347
rect	175	349	176	350
rect	175	355	176	356
rect	175	361	176	362
rect	175	364	176	365
rect	175	367	176	368
rect	176	1	177	2
rect	176	4	177	5
rect	176	7	177	8
rect	176	10	177	11
rect	176	13	177	14
rect	176	16	177	17
rect	176	19	177	20
rect	176	22	177	23
rect	176	25	177	26
rect	176	28	177	29
rect	176	31	177	32
rect	176	34	177	35
rect	176	37	177	38
rect	176	40	177	41
rect	176	43	177	44
rect	176	46	177	47
rect	176	49	177	50
rect	176	52	177	53
rect	176	55	177	56
rect	176	58	177	59
rect	176	61	177	62
rect	176	64	177	65
rect	176	67	177	68
rect	176	70	177	71
rect	176	73	177	74
rect	176	76	177	77
rect	176	79	177	80
rect	176	82	177	83
rect	176	85	177	86
rect	176	88	177	89
rect	176	91	177	92
rect	176	94	177	95
rect	176	97	177	98
rect	176	100	177	101
rect	176	103	177	104
rect	176	106	177	107
rect	176	109	177	110
rect	176	112	177	113
rect	176	115	177	116
rect	176	118	177	119
rect	176	121	177	122
rect	176	124	177	125
rect	176	127	177	128
rect	176	130	177	131
rect	176	133	177	134
rect	176	136	177	137
rect	176	139	177	140
rect	176	142	177	143
rect	176	145	177	146
rect	176	148	177	149
rect	176	151	177	152
rect	176	154	177	155
rect	176	157	177	158
rect	176	160	177	161
rect	176	163	177	164
rect	176	166	177	167
rect	176	169	177	170
rect	176	172	177	173
rect	176	175	177	176
rect	176	178	177	179
rect	176	181	177	182
rect	176	184	177	185
rect	176	187	177	188
rect	176	190	177	191
rect	176	193	177	194
rect	176	196	177	197
rect	176	199	177	200
rect	176	202	177	203
rect	176	205	177	206
rect	176	208	177	209
rect	176	211	177	212
rect	176	214	177	215
rect	176	217	177	218
rect	176	220	177	221
rect	176	223	177	224
rect	176	226	177	227
rect	176	229	177	230
rect	176	232	177	233
rect	176	235	177	236
rect	176	238	177	239
rect	176	241	177	242
rect	176	244	177	245
rect	176	247	177	248
rect	176	250	177	251
rect	176	253	177	254
rect	176	256	177	257
rect	176	259	177	260
rect	176	262	177	263
rect	176	265	177	266
rect	176	268	177	269
rect	176	271	177	272
rect	176	274	177	275
rect	176	277	177	278
rect	176	280	177	281
rect	176	283	177	284
rect	176	286	177	287
rect	176	289	177	290
rect	176	292	177	293
rect	176	295	177	296
rect	176	298	177	299
rect	176	301	177	302
rect	176	307	177	308
rect	176	310	177	311
rect	176	313	177	314
rect	176	316	177	317
rect	176	322	177	323
rect	176	325	177	326
rect	176	331	177	332
rect	176	334	177	335
rect	176	346	177	347
rect	176	349	177	350
rect	176	355	177	356
rect	176	361	177	362
rect	176	364	177	365
rect	176	367	177	368
rect	177	1	178	2
rect	177	4	178	5
rect	177	7	178	8
rect	177	10	178	11
rect	177	13	178	14
rect	177	16	178	17
rect	177	19	178	20
rect	177	22	178	23
rect	177	25	178	26
rect	177	28	178	29
rect	177	31	178	32
rect	177	34	178	35
rect	177	37	178	38
rect	177	40	178	41
rect	177	43	178	44
rect	177	46	178	47
rect	177	49	178	50
rect	177	52	178	53
rect	177	55	178	56
rect	177	58	178	59
rect	177	61	178	62
rect	177	64	178	65
rect	177	67	178	68
rect	177	70	178	71
rect	177	73	178	74
rect	177	76	178	77
rect	177	79	178	80
rect	177	82	178	83
rect	177	85	178	86
rect	177	88	178	89
rect	177	91	178	92
rect	177	94	178	95
rect	177	97	178	98
rect	177	100	178	101
rect	177	103	178	104
rect	177	106	178	107
rect	177	109	178	110
rect	177	112	178	113
rect	177	115	178	116
rect	177	118	178	119
rect	177	121	178	122
rect	177	124	178	125
rect	177	127	178	128
rect	177	130	178	131
rect	177	133	178	134
rect	177	136	178	137
rect	177	139	178	140
rect	177	142	178	143
rect	177	145	178	146
rect	177	148	178	149
rect	177	151	178	152
rect	177	154	178	155
rect	177	157	178	158
rect	177	160	178	161
rect	177	163	178	164
rect	177	166	178	167
rect	177	169	178	170
rect	177	172	178	173
rect	177	175	178	176
rect	177	178	178	179
rect	177	181	178	182
rect	177	184	178	185
rect	177	187	178	188
rect	177	190	178	191
rect	177	193	178	194
rect	177	196	178	197
rect	177	199	178	200
rect	177	202	178	203
rect	177	205	178	206
rect	177	208	178	209
rect	177	211	178	212
rect	177	214	178	215
rect	177	217	178	218
rect	177	220	178	221
rect	177	223	178	224
rect	177	226	178	227
rect	177	229	178	230
rect	177	232	178	233
rect	177	235	178	236
rect	177	238	178	239
rect	177	241	178	242
rect	177	244	178	245
rect	177	247	178	248
rect	177	250	178	251
rect	177	253	178	254
rect	177	256	178	257
rect	177	259	178	260
rect	177	262	178	263
rect	177	265	178	266
rect	177	268	178	269
rect	177	271	178	272
rect	177	274	178	275
rect	177	277	178	278
rect	177	280	178	281
rect	177	283	178	284
rect	177	286	178	287
rect	177	289	178	290
rect	177	292	178	293
rect	177	295	178	296
rect	177	298	178	299
rect	177	301	178	302
rect	177	307	178	308
rect	177	310	178	311
rect	177	313	178	314
rect	177	316	178	317
rect	177	322	178	323
rect	177	325	178	326
rect	177	331	178	332
rect	177	334	178	335
rect	177	346	178	347
rect	177	349	178	350
rect	177	355	178	356
rect	177	361	178	362
rect	177	364	178	365
rect	177	367	178	368
rect	178	1	179	2
rect	178	4	179	5
rect	178	7	179	8
rect	178	10	179	11
rect	178	13	179	14
rect	178	16	179	17
rect	178	19	179	20
rect	178	22	179	23
rect	178	25	179	26
rect	178	28	179	29
rect	178	31	179	32
rect	178	34	179	35
rect	178	37	179	38
rect	178	40	179	41
rect	178	43	179	44
rect	178	46	179	47
rect	178	49	179	50
rect	178	52	179	53
rect	178	55	179	56
rect	178	58	179	59
rect	178	61	179	62
rect	178	64	179	65
rect	178	67	179	68
rect	178	70	179	71
rect	178	73	179	74
rect	178	76	179	77
rect	178	79	179	80
rect	178	82	179	83
rect	178	85	179	86
rect	178	88	179	89
rect	178	91	179	92
rect	178	94	179	95
rect	178	97	179	98
rect	178	100	179	101
rect	178	103	179	104
rect	178	106	179	107
rect	178	109	179	110
rect	178	112	179	113
rect	178	115	179	116
rect	178	118	179	119
rect	178	121	179	122
rect	178	124	179	125
rect	178	127	179	128
rect	178	130	179	131
rect	178	133	179	134
rect	178	136	179	137
rect	178	139	179	140
rect	178	142	179	143
rect	178	145	179	146
rect	178	148	179	149
rect	178	151	179	152
rect	178	154	179	155
rect	178	157	179	158
rect	178	160	179	161
rect	178	163	179	164
rect	178	166	179	167
rect	178	169	179	170
rect	178	172	179	173
rect	178	175	179	176
rect	178	178	179	179
rect	178	181	179	182
rect	178	184	179	185
rect	178	187	179	188
rect	178	190	179	191
rect	178	193	179	194
rect	178	196	179	197
rect	178	199	179	200
rect	178	202	179	203
rect	178	205	179	206
rect	178	208	179	209
rect	178	211	179	212
rect	178	214	179	215
rect	178	217	179	218
rect	178	220	179	221
rect	178	223	179	224
rect	178	226	179	227
rect	178	229	179	230
rect	178	232	179	233
rect	178	235	179	236
rect	178	238	179	239
rect	178	241	179	242
rect	178	244	179	245
rect	178	247	179	248
rect	178	250	179	251
rect	178	253	179	254
rect	178	256	179	257
rect	178	259	179	260
rect	178	262	179	263
rect	178	265	179	266
rect	178	268	179	269
rect	178	271	179	272
rect	178	274	179	275
rect	178	277	179	278
rect	178	280	179	281
rect	178	283	179	284
rect	178	286	179	287
rect	178	289	179	290
rect	178	292	179	293
rect	178	295	179	296
rect	178	298	179	299
rect	178	301	179	302
rect	178	307	179	308
rect	178	310	179	311
rect	178	313	179	314
rect	178	316	179	317
rect	178	322	179	323
rect	178	325	179	326
rect	178	331	179	332
rect	178	334	179	335
rect	178	346	179	347
rect	178	349	179	350
rect	178	355	179	356
rect	178	361	179	362
rect	178	364	179	365
rect	178	367	179	368
rect	179	1	180	2
rect	179	4	180	5
rect	179	7	180	8
rect	179	10	180	11
rect	179	13	180	14
rect	179	16	180	17
rect	179	19	180	20
rect	179	22	180	23
rect	179	25	180	26
rect	179	28	180	29
rect	179	31	180	32
rect	179	34	180	35
rect	179	37	180	38
rect	179	40	180	41
rect	179	43	180	44
rect	179	46	180	47
rect	179	49	180	50
rect	179	52	180	53
rect	179	55	180	56
rect	179	58	180	59
rect	179	61	180	62
rect	179	64	180	65
rect	179	67	180	68
rect	179	70	180	71
rect	179	73	180	74
rect	179	76	180	77
rect	179	79	180	80
rect	179	82	180	83
rect	179	85	180	86
rect	179	88	180	89
rect	179	91	180	92
rect	179	94	180	95
rect	179	97	180	98
rect	179	100	180	101
rect	179	103	180	104
rect	179	106	180	107
rect	179	109	180	110
rect	179	112	180	113
rect	179	115	180	116
rect	179	118	180	119
rect	179	121	180	122
rect	179	124	180	125
rect	179	127	180	128
rect	179	130	180	131
rect	179	133	180	134
rect	179	136	180	137
rect	179	139	180	140
rect	179	142	180	143
rect	179	145	180	146
rect	179	148	180	149
rect	179	151	180	152
rect	179	154	180	155
rect	179	157	180	158
rect	179	160	180	161
rect	179	163	180	164
rect	179	166	180	167
rect	179	169	180	170
rect	179	172	180	173
rect	179	175	180	176
rect	179	178	180	179
rect	179	181	180	182
rect	179	184	180	185
rect	179	187	180	188
rect	179	190	180	191
rect	179	193	180	194
rect	179	196	180	197
rect	179	199	180	200
rect	179	202	180	203
rect	179	205	180	206
rect	179	208	180	209
rect	179	211	180	212
rect	179	214	180	215
rect	179	217	180	218
rect	179	220	180	221
rect	179	223	180	224
rect	179	226	180	227
rect	179	229	180	230
rect	179	232	180	233
rect	179	235	180	236
rect	179	238	180	239
rect	179	241	180	242
rect	179	244	180	245
rect	179	247	180	248
rect	179	250	180	251
rect	179	253	180	254
rect	179	256	180	257
rect	179	259	180	260
rect	179	262	180	263
rect	179	265	180	266
rect	179	268	180	269
rect	179	271	180	272
rect	179	274	180	275
rect	179	277	180	278
rect	179	280	180	281
rect	179	283	180	284
rect	179	286	180	287
rect	179	289	180	290
rect	179	292	180	293
rect	179	295	180	296
rect	179	298	180	299
rect	179	301	180	302
rect	179	307	180	308
rect	179	310	180	311
rect	179	313	180	314
rect	179	316	180	317
rect	179	322	180	323
rect	179	325	180	326
rect	179	331	180	332
rect	179	334	180	335
rect	179	346	180	347
rect	179	349	180	350
rect	179	355	180	356
rect	179	361	180	362
rect	179	364	180	365
rect	179	367	180	368
rect	180	1	181	2
rect	180	4	181	5
rect	180	7	181	8
rect	180	10	181	11
rect	180	13	181	14
rect	180	16	181	17
rect	180	19	181	20
rect	180	22	181	23
rect	180	25	181	26
rect	180	28	181	29
rect	180	31	181	32
rect	180	34	181	35
rect	180	37	181	38
rect	180	40	181	41
rect	180	43	181	44
rect	180	46	181	47
rect	180	49	181	50
rect	180	52	181	53
rect	180	55	181	56
rect	180	58	181	59
rect	180	61	181	62
rect	180	64	181	65
rect	180	67	181	68
rect	180	70	181	71
rect	180	73	181	74
rect	180	76	181	77
rect	180	79	181	80
rect	180	82	181	83
rect	180	85	181	86
rect	180	88	181	89
rect	180	91	181	92
rect	180	94	181	95
rect	180	97	181	98
rect	180	100	181	101
rect	180	103	181	104
rect	180	106	181	107
rect	180	109	181	110
rect	180	112	181	113
rect	180	115	181	116
rect	180	118	181	119
rect	180	121	181	122
rect	180	124	181	125
rect	180	127	181	128
rect	180	130	181	131
rect	180	133	181	134
rect	180	136	181	137
rect	180	139	181	140
rect	180	142	181	143
rect	180	145	181	146
rect	180	148	181	149
rect	180	151	181	152
rect	180	154	181	155
rect	180	157	181	158
rect	180	160	181	161
rect	180	163	181	164
rect	180	166	181	167
rect	180	169	181	170
rect	180	172	181	173
rect	180	175	181	176
rect	180	178	181	179
rect	180	181	181	182
rect	180	184	181	185
rect	180	187	181	188
rect	180	190	181	191
rect	180	193	181	194
rect	180	196	181	197
rect	180	199	181	200
rect	180	202	181	203
rect	180	205	181	206
rect	180	208	181	209
rect	180	211	181	212
rect	180	214	181	215
rect	180	217	181	218
rect	180	220	181	221
rect	180	223	181	224
rect	180	226	181	227
rect	180	229	181	230
rect	180	232	181	233
rect	180	235	181	236
rect	180	238	181	239
rect	180	241	181	242
rect	180	244	181	245
rect	180	247	181	248
rect	180	250	181	251
rect	180	253	181	254
rect	180	256	181	257
rect	180	259	181	260
rect	180	262	181	263
rect	180	265	181	266
rect	180	268	181	269
rect	180	271	181	272
rect	180	274	181	275
rect	180	277	181	278
rect	180	280	181	281
rect	180	283	181	284
rect	180	286	181	287
rect	180	289	181	290
rect	180	292	181	293
rect	180	295	181	296
rect	180	298	181	299
rect	180	301	181	302
rect	180	310	181	311
rect	180	313	181	314
rect	180	316	181	317
rect	180	322	181	323
rect	180	325	181	326
rect	180	331	181	332
rect	180	334	181	335
rect	180	346	181	347
rect	180	349	181	350
rect	180	355	181	356
rect	180	361	181	362
rect	180	364	181	365
rect	180	367	181	368
rect	181	1	182	2
rect	181	4	182	5
rect	181	7	182	8
rect	181	10	182	11
rect	181	13	182	14
rect	181	16	182	17
rect	181	19	182	20
rect	181	22	182	23
rect	181	25	182	26
rect	181	28	182	29
rect	181	31	182	32
rect	181	34	182	35
rect	181	37	182	38
rect	181	40	182	41
rect	181	43	182	44
rect	181	46	182	47
rect	181	49	182	50
rect	181	52	182	53
rect	181	55	182	56
rect	181	58	182	59
rect	181	61	182	62
rect	181	64	182	65
rect	181	67	182	68
rect	181	70	182	71
rect	181	73	182	74
rect	181	76	182	77
rect	181	79	182	80
rect	181	82	182	83
rect	181	85	182	86
rect	181	88	182	89
rect	181	91	182	92
rect	181	94	182	95
rect	181	97	182	98
rect	181	100	182	101
rect	181	103	182	104
rect	181	106	182	107
rect	181	109	182	110
rect	181	112	182	113
rect	181	115	182	116
rect	181	118	182	119
rect	181	121	182	122
rect	181	124	182	125
rect	181	127	182	128
rect	181	130	182	131
rect	181	133	182	134
rect	181	136	182	137
rect	181	139	182	140
rect	181	142	182	143
rect	181	145	182	146
rect	181	148	182	149
rect	181	151	182	152
rect	181	154	182	155
rect	181	157	182	158
rect	181	160	182	161
rect	181	163	182	164
rect	181	166	182	167
rect	181	169	182	170
rect	181	172	182	173
rect	181	175	182	176
rect	181	178	182	179
rect	181	181	182	182
rect	181	184	182	185
rect	181	187	182	188
rect	181	190	182	191
rect	181	193	182	194
rect	181	196	182	197
rect	181	199	182	200
rect	181	202	182	203
rect	181	205	182	206
rect	181	208	182	209
rect	181	211	182	212
rect	181	214	182	215
rect	181	217	182	218
rect	181	220	182	221
rect	181	223	182	224
rect	181	226	182	227
rect	181	229	182	230
rect	181	232	182	233
rect	181	235	182	236
rect	181	238	182	239
rect	181	241	182	242
rect	181	244	182	245
rect	181	247	182	248
rect	181	250	182	251
rect	181	253	182	254
rect	181	256	182	257
rect	181	259	182	260
rect	181	262	182	263
rect	181	265	182	266
rect	181	268	182	269
rect	181	271	182	272
rect	181	274	182	275
rect	181	277	182	278
rect	181	280	182	281
rect	181	283	182	284
rect	181	286	182	287
rect	181	289	182	290
rect	181	292	182	293
rect	181	295	182	296
rect	181	298	182	299
rect	181	301	182	302
rect	181	307	182	308
rect	181	310	182	311
rect	181	313	182	314
rect	181	316	182	317
rect	181	322	182	323
rect	181	325	182	326
rect	181	331	182	332
rect	181	334	182	335
rect	181	346	182	347
rect	181	349	182	350
rect	181	355	182	356
rect	181	361	182	362
rect	181	364	182	365
rect	181	367	182	368
rect	182	1	183	2
rect	182	4	183	5
rect	182	7	183	8
rect	182	10	183	11
rect	182	13	183	14
rect	182	16	183	17
rect	182	19	183	20
rect	182	22	183	23
rect	182	25	183	26
rect	182	28	183	29
rect	182	31	183	32
rect	182	34	183	35
rect	182	37	183	38
rect	182	40	183	41
rect	182	43	183	44
rect	182	46	183	47
rect	182	49	183	50
rect	182	52	183	53
rect	182	55	183	56
rect	182	58	183	59
rect	182	61	183	62
rect	182	64	183	65
rect	182	67	183	68
rect	182	70	183	71
rect	182	73	183	74
rect	182	76	183	77
rect	182	79	183	80
rect	182	82	183	83
rect	182	85	183	86
rect	182	88	183	89
rect	182	91	183	92
rect	182	94	183	95
rect	182	97	183	98
rect	182	100	183	101
rect	182	103	183	104
rect	182	106	183	107
rect	182	109	183	110
rect	182	112	183	113
rect	182	115	183	116
rect	182	118	183	119
rect	182	121	183	122
rect	182	124	183	125
rect	182	127	183	128
rect	182	130	183	131
rect	182	133	183	134
rect	182	136	183	137
rect	182	139	183	140
rect	182	142	183	143
rect	182	145	183	146
rect	182	148	183	149
rect	182	151	183	152
rect	182	154	183	155
rect	182	157	183	158
rect	182	160	183	161
rect	182	163	183	164
rect	182	166	183	167
rect	182	169	183	170
rect	182	172	183	173
rect	182	175	183	176
rect	182	178	183	179
rect	182	181	183	182
rect	182	184	183	185
rect	182	187	183	188
rect	182	190	183	191
rect	182	193	183	194
rect	182	196	183	197
rect	182	199	183	200
rect	182	202	183	203
rect	182	205	183	206
rect	182	208	183	209
rect	182	211	183	212
rect	182	214	183	215
rect	182	217	183	218
rect	182	220	183	221
rect	182	223	183	224
rect	182	226	183	227
rect	182	229	183	230
rect	182	232	183	233
rect	182	235	183	236
rect	182	238	183	239
rect	182	241	183	242
rect	182	244	183	245
rect	182	247	183	248
rect	182	250	183	251
rect	182	253	183	254
rect	182	256	183	257
rect	182	259	183	260
rect	182	262	183	263
rect	182	268	183	269
rect	182	271	183	272
rect	182	274	183	275
rect	182	277	183	278
rect	182	280	183	281
rect	182	283	183	284
rect	182	286	183	287
rect	182	289	183	290
rect	182	292	183	293
rect	182	295	183	296
rect	182	298	183	299
rect	182	301	183	302
rect	182	307	183	308
rect	182	310	183	311
rect	182	313	183	314
rect	182	316	183	317
rect	182	322	183	323
rect	182	325	183	326
rect	182	331	183	332
rect	182	334	183	335
rect	182	346	183	347
rect	182	349	183	350
rect	182	355	183	356
rect	182	361	183	362
rect	182	364	183	365
rect	182	367	183	368
rect	183	1	184	2
rect	183	4	184	5
rect	183	7	184	8
rect	183	10	184	11
rect	183	13	184	14
rect	183	16	184	17
rect	183	19	184	20
rect	183	22	184	23
rect	183	25	184	26
rect	183	28	184	29
rect	183	31	184	32
rect	183	34	184	35
rect	183	37	184	38
rect	183	40	184	41
rect	183	43	184	44
rect	183	46	184	47
rect	183	49	184	50
rect	183	52	184	53
rect	183	55	184	56
rect	183	58	184	59
rect	183	61	184	62
rect	183	64	184	65
rect	183	67	184	68
rect	183	70	184	71
rect	183	73	184	74
rect	183	76	184	77
rect	183	79	184	80
rect	183	82	184	83
rect	183	85	184	86
rect	183	88	184	89
rect	183	91	184	92
rect	183	94	184	95
rect	183	97	184	98
rect	183	100	184	101
rect	183	103	184	104
rect	183	106	184	107
rect	183	109	184	110
rect	183	112	184	113
rect	183	115	184	116
rect	183	118	184	119
rect	183	121	184	122
rect	183	124	184	125
rect	183	127	184	128
rect	183	130	184	131
rect	183	133	184	134
rect	183	136	184	137
rect	183	139	184	140
rect	183	142	184	143
rect	183	145	184	146
rect	183	148	184	149
rect	183	151	184	152
rect	183	154	184	155
rect	183	157	184	158
rect	183	160	184	161
rect	183	163	184	164
rect	183	166	184	167
rect	183	169	184	170
rect	183	172	184	173
rect	183	175	184	176
rect	183	178	184	179
rect	183	181	184	182
rect	183	184	184	185
rect	183	187	184	188
rect	183	190	184	191
rect	183	193	184	194
rect	183	196	184	197
rect	183	199	184	200
rect	183	202	184	203
rect	183	205	184	206
rect	183	208	184	209
rect	183	211	184	212
rect	183	214	184	215
rect	183	217	184	218
rect	183	220	184	221
rect	183	223	184	224
rect	183	226	184	227
rect	183	229	184	230
rect	183	232	184	233
rect	183	235	184	236
rect	183	238	184	239
rect	183	241	184	242
rect	183	244	184	245
rect	183	247	184	248
rect	183	250	184	251
rect	183	253	184	254
rect	183	256	184	257
rect	183	259	184	260
rect	183	262	184	263
rect	183	265	184	266
rect	183	268	184	269
rect	183	271	184	272
rect	183	274	184	275
rect	183	277	184	278
rect	183	280	184	281
rect	183	283	184	284
rect	183	286	184	287
rect	183	289	184	290
rect	183	292	184	293
rect	183	295	184	296
rect	183	298	184	299
rect	183	301	184	302
rect	183	307	184	308
rect	183	310	184	311
rect	183	313	184	314
rect	183	316	184	317
rect	183	322	184	323
rect	183	325	184	326
rect	183	331	184	332
rect	183	334	184	335
rect	183	346	184	347
rect	183	349	184	350
rect	183	355	184	356
rect	183	361	184	362
rect	183	364	184	365
rect	183	367	184	368
rect	184	1	185	2
rect	184	4	185	5
rect	184	7	185	8
rect	184	10	185	11
rect	184	13	185	14
rect	184	16	185	17
rect	184	19	185	20
rect	184	22	185	23
rect	184	25	185	26
rect	184	28	185	29
rect	184	31	185	32
rect	184	34	185	35
rect	184	37	185	38
rect	184	40	185	41
rect	184	43	185	44
rect	184	46	185	47
rect	184	49	185	50
rect	184	52	185	53
rect	184	55	185	56
rect	184	58	185	59
rect	184	61	185	62
rect	184	64	185	65
rect	184	67	185	68
rect	184	70	185	71
rect	184	73	185	74
rect	184	76	185	77
rect	184	79	185	80
rect	184	82	185	83
rect	184	85	185	86
rect	184	88	185	89
rect	184	91	185	92
rect	184	94	185	95
rect	184	97	185	98
rect	184	100	185	101
rect	184	103	185	104
rect	184	106	185	107
rect	184	109	185	110
rect	184	112	185	113
rect	184	115	185	116
rect	184	118	185	119
rect	184	121	185	122
rect	184	124	185	125
rect	184	127	185	128
rect	184	130	185	131
rect	184	133	185	134
rect	184	136	185	137
rect	184	139	185	140
rect	184	142	185	143
rect	184	145	185	146
rect	184	148	185	149
rect	184	151	185	152
rect	184	154	185	155
rect	184	157	185	158
rect	184	160	185	161
rect	184	163	185	164
rect	184	166	185	167
rect	184	169	185	170
rect	184	172	185	173
rect	184	175	185	176
rect	184	178	185	179
rect	184	181	185	182
rect	184	184	185	185
rect	184	187	185	188
rect	184	190	185	191
rect	184	193	185	194
rect	184	196	185	197
rect	184	199	185	200
rect	184	202	185	203
rect	184	205	185	206
rect	184	208	185	209
rect	184	211	185	212
rect	184	214	185	215
rect	184	217	185	218
rect	184	220	185	221
rect	184	223	185	224
rect	184	226	185	227
rect	184	229	185	230
rect	184	232	185	233
rect	184	235	185	236
rect	184	238	185	239
rect	184	241	185	242
rect	184	244	185	245
rect	184	247	185	248
rect	184	250	185	251
rect	184	253	185	254
rect	184	256	185	257
rect	184	259	185	260
rect	184	262	185	263
rect	184	265	185	266
rect	184	268	185	269
rect	184	271	185	272
rect	184	274	185	275
rect	184	277	185	278
rect	184	280	185	281
rect	184	283	185	284
rect	184	286	185	287
rect	184	289	185	290
rect	184	292	185	293
rect	184	295	185	296
rect	184	298	185	299
rect	184	301	185	302
rect	184	307	185	308
rect	184	310	185	311
rect	184	313	185	314
rect	184	316	185	317
rect	184	322	185	323
rect	184	325	185	326
rect	184	331	185	332
rect	184	334	185	335
rect	184	346	185	347
rect	184	349	185	350
rect	184	355	185	356
rect	184	361	185	362
rect	184	364	185	365
rect	184	367	185	368
rect	185	1	186	2
rect	185	4	186	5
rect	185	7	186	8
rect	185	10	186	11
rect	185	13	186	14
rect	185	16	186	17
rect	185	19	186	20
rect	185	22	186	23
rect	185	25	186	26
rect	185	28	186	29
rect	185	31	186	32
rect	185	34	186	35
rect	185	37	186	38
rect	185	40	186	41
rect	185	43	186	44
rect	185	46	186	47
rect	185	49	186	50
rect	185	52	186	53
rect	185	55	186	56
rect	185	58	186	59
rect	185	61	186	62
rect	185	64	186	65
rect	185	67	186	68
rect	185	70	186	71
rect	185	73	186	74
rect	185	76	186	77
rect	185	79	186	80
rect	185	82	186	83
rect	185	85	186	86
rect	185	88	186	89
rect	185	91	186	92
rect	185	94	186	95
rect	185	97	186	98
rect	185	100	186	101
rect	185	103	186	104
rect	185	106	186	107
rect	185	109	186	110
rect	185	112	186	113
rect	185	115	186	116
rect	185	118	186	119
rect	185	121	186	122
rect	185	124	186	125
rect	185	127	186	128
rect	185	130	186	131
rect	185	133	186	134
rect	185	136	186	137
rect	185	139	186	140
rect	185	142	186	143
rect	185	145	186	146
rect	185	148	186	149
rect	185	151	186	152
rect	185	154	186	155
rect	185	157	186	158
rect	185	160	186	161
rect	185	163	186	164
rect	185	166	186	167
rect	185	169	186	170
rect	185	172	186	173
rect	185	175	186	176
rect	185	178	186	179
rect	185	181	186	182
rect	185	184	186	185
rect	185	187	186	188
rect	185	190	186	191
rect	185	193	186	194
rect	185	196	186	197
rect	185	199	186	200
rect	185	202	186	203
rect	185	205	186	206
rect	185	208	186	209
rect	185	211	186	212
rect	185	214	186	215
rect	185	217	186	218
rect	185	220	186	221
rect	185	223	186	224
rect	185	226	186	227
rect	185	229	186	230
rect	185	232	186	233
rect	185	235	186	236
rect	185	238	186	239
rect	185	241	186	242
rect	185	244	186	245
rect	185	247	186	248
rect	185	250	186	251
rect	185	253	186	254
rect	185	256	186	257
rect	185	259	186	260
rect	185	262	186	263
rect	185	265	186	266
rect	185	268	186	269
rect	185	271	186	272
rect	185	274	186	275
rect	185	277	186	278
rect	185	280	186	281
rect	185	283	186	284
rect	185	286	186	287
rect	185	289	186	290
rect	185	292	186	293
rect	185	295	186	296
rect	185	298	186	299
rect	185	301	186	302
rect	185	307	186	308
rect	185	310	186	311
rect	185	313	186	314
rect	185	316	186	317
rect	185	322	186	323
rect	185	325	186	326
rect	185	331	186	332
rect	185	334	186	335
rect	185	346	186	347
rect	185	349	186	350
rect	185	355	186	356
rect	185	361	186	362
rect	185	364	186	365
rect	185	367	186	368
rect	186	1	187	2
rect	186	4	187	5
rect	186	7	187	8
rect	186	10	187	11
rect	186	13	187	14
rect	186	16	187	17
rect	186	19	187	20
rect	186	22	187	23
rect	186	25	187	26
rect	186	28	187	29
rect	186	31	187	32
rect	186	34	187	35
rect	186	37	187	38
rect	186	40	187	41
rect	186	43	187	44
rect	186	46	187	47
rect	186	49	187	50
rect	186	52	187	53
rect	186	55	187	56
rect	186	58	187	59
rect	186	61	187	62
rect	186	64	187	65
rect	186	67	187	68
rect	186	70	187	71
rect	186	73	187	74
rect	186	76	187	77
rect	186	79	187	80
rect	186	82	187	83
rect	186	85	187	86
rect	186	88	187	89
rect	186	91	187	92
rect	186	94	187	95
rect	186	97	187	98
rect	186	100	187	101
rect	186	103	187	104
rect	186	106	187	107
rect	186	109	187	110
rect	186	112	187	113
rect	186	115	187	116
rect	186	118	187	119
rect	186	121	187	122
rect	186	124	187	125
rect	186	127	187	128
rect	186	130	187	131
rect	186	133	187	134
rect	186	136	187	137
rect	186	139	187	140
rect	186	142	187	143
rect	186	145	187	146
rect	186	148	187	149
rect	186	151	187	152
rect	186	154	187	155
rect	186	157	187	158
rect	186	160	187	161
rect	186	163	187	164
rect	186	166	187	167
rect	186	169	187	170
rect	186	172	187	173
rect	186	175	187	176
rect	186	178	187	179
rect	186	181	187	182
rect	186	184	187	185
rect	186	187	187	188
rect	186	190	187	191
rect	186	193	187	194
rect	186	196	187	197
rect	186	199	187	200
rect	186	202	187	203
rect	186	205	187	206
rect	186	208	187	209
rect	186	211	187	212
rect	186	214	187	215
rect	186	217	187	218
rect	186	220	187	221
rect	186	223	187	224
rect	186	226	187	227
rect	186	229	187	230
rect	186	232	187	233
rect	186	235	187	236
rect	186	238	187	239
rect	186	241	187	242
rect	186	244	187	245
rect	186	247	187	248
rect	186	250	187	251
rect	186	253	187	254
rect	186	256	187	257
rect	186	259	187	260
rect	186	262	187	263
rect	186	265	187	266
rect	186	268	187	269
rect	186	271	187	272
rect	186	274	187	275
rect	186	277	187	278
rect	186	280	187	281
rect	186	283	187	284
rect	186	286	187	287
rect	186	289	187	290
rect	186	292	187	293
rect	186	295	187	296
rect	186	298	187	299
rect	186	301	187	302
rect	186	307	187	308
rect	186	310	187	311
rect	186	313	187	314
rect	186	316	187	317
rect	186	322	187	323
rect	186	325	187	326
rect	186	331	187	332
rect	186	334	187	335
rect	186	346	187	347
rect	186	349	187	350
rect	186	355	187	356
rect	186	361	187	362
rect	186	364	187	365
rect	186	367	187	368
rect	187	4	188	5
rect	187	7	188	8
rect	187	10	188	11
rect	187	13	188	14
rect	187	16	188	17
rect	187	19	188	20
rect	187	22	188	23
rect	187	25	188	26
rect	187	28	188	29
rect	187	31	188	32
rect	187	34	188	35
rect	187	37	188	38
rect	187	40	188	41
rect	187	43	188	44
rect	187	46	188	47
rect	187	49	188	50
rect	187	52	188	53
rect	187	55	188	56
rect	187	58	188	59
rect	187	61	188	62
rect	187	64	188	65
rect	187	67	188	68
rect	187	70	188	71
rect	187	73	188	74
rect	187	76	188	77
rect	187	79	188	80
rect	187	82	188	83
rect	187	85	188	86
rect	187	88	188	89
rect	187	91	188	92
rect	187	94	188	95
rect	187	97	188	98
rect	187	100	188	101
rect	187	103	188	104
rect	187	106	188	107
rect	187	109	188	110
rect	187	112	188	113
rect	187	115	188	116
rect	187	118	188	119
rect	187	121	188	122
rect	187	124	188	125
rect	187	127	188	128
rect	187	130	188	131
rect	187	133	188	134
rect	187	136	188	137
rect	187	139	188	140
rect	187	142	188	143
rect	187	145	188	146
rect	187	148	188	149
rect	187	151	188	152
rect	187	154	188	155
rect	187	157	188	158
rect	187	160	188	161
rect	187	163	188	164
rect	187	166	188	167
rect	187	169	188	170
rect	187	172	188	173
rect	187	175	188	176
rect	187	178	188	179
rect	187	181	188	182
rect	187	184	188	185
rect	187	187	188	188
rect	187	190	188	191
rect	187	193	188	194
rect	187	196	188	197
rect	187	199	188	200
rect	187	202	188	203
rect	187	205	188	206
rect	187	208	188	209
rect	187	211	188	212
rect	187	214	188	215
rect	187	217	188	218
rect	187	220	188	221
rect	187	223	188	224
rect	187	226	188	227
rect	187	229	188	230
rect	187	232	188	233
rect	187	235	188	236
rect	187	238	188	239
rect	187	241	188	242
rect	187	244	188	245
rect	187	247	188	248
rect	187	250	188	251
rect	187	253	188	254
rect	187	256	188	257
rect	187	259	188	260
rect	187	262	188	263
rect	187	265	188	266
rect	187	268	188	269
rect	187	271	188	272
rect	187	274	188	275
rect	187	277	188	278
rect	187	280	188	281
rect	187	283	188	284
rect	187	286	188	287
rect	187	289	188	290
rect	187	292	188	293
rect	187	295	188	296
rect	187	298	188	299
rect	187	301	188	302
rect	187	307	188	308
rect	187	310	188	311
rect	187	313	188	314
rect	187	316	188	317
rect	187	322	188	323
rect	187	325	188	326
rect	187	331	188	332
rect	187	334	188	335
rect	187	346	188	347
rect	187	349	188	350
rect	187	364	188	365
rect	188	4	189	5
rect	188	7	189	8
rect	188	10	189	11
rect	188	13	189	14
rect	188	16	189	17
rect	188	22	189	23
rect	188	25	189	26
rect	188	28	189	29
rect	188	31	189	32
rect	188	34	189	35
rect	188	37	189	38
rect	188	40	189	41
rect	188	43	189	44
rect	188	46	189	47
rect	188	49	189	50
rect	188	52	189	53
rect	188	55	189	56
rect	188	58	189	59
rect	188	61	189	62
rect	188	64	189	65
rect	188	67	189	68
rect	188	70	189	71
rect	188	73	189	74
rect	188	76	189	77
rect	188	79	189	80
rect	188	82	189	83
rect	188	85	189	86
rect	188	88	189	89
rect	188	91	189	92
rect	188	94	189	95
rect	188	97	189	98
rect	188	100	189	101
rect	188	103	189	104
rect	188	106	189	107
rect	188	109	189	110
rect	188	112	189	113
rect	188	115	189	116
rect	188	118	189	119
rect	188	121	189	122
rect	188	124	189	125
rect	188	127	189	128
rect	188	130	189	131
rect	188	133	189	134
rect	188	136	189	137
rect	188	139	189	140
rect	188	142	189	143
rect	188	145	189	146
rect	188	148	189	149
rect	188	151	189	152
rect	188	154	189	155
rect	188	157	189	158
rect	188	160	189	161
rect	188	163	189	164
rect	188	166	189	167
rect	188	169	189	170
rect	188	172	189	173
rect	188	175	189	176
rect	188	178	189	179
rect	188	181	189	182
rect	188	184	189	185
rect	188	187	189	188
rect	188	190	189	191
rect	188	193	189	194
rect	188	196	189	197
rect	188	199	189	200
rect	188	202	189	203
rect	188	205	189	206
rect	188	208	189	209
rect	188	211	189	212
rect	188	214	189	215
rect	188	217	189	218
rect	188	220	189	221
rect	188	223	189	224
rect	188	226	189	227
rect	188	229	189	230
rect	188	235	189	236
rect	188	238	189	239
rect	188	241	189	242
rect	188	244	189	245
rect	188	247	189	248
rect	188	250	189	251
rect	188	253	189	254
rect	188	256	189	257
rect	188	259	189	260
rect	188	262	189	263
rect	188	265	189	266
rect	188	268	189	269
rect	188	271	189	272
rect	188	274	189	275
rect	188	277	189	278
rect	188	280	189	281
rect	188	283	189	284
rect	188	286	189	287
rect	188	289	189	290
rect	188	292	189	293
rect	188	295	189	296
rect	188	298	189	299
rect	188	301	189	302
rect	188	307	189	308
rect	188	310	189	311
rect	188	313	189	314
rect	188	316	189	317
rect	188	322	189	323
rect	188	325	189	326
rect	188	331	189	332
rect	188	334	189	335
rect	188	346	189	347
rect	188	349	189	350
rect	188	364	189	365
rect	189	4	190	5
rect	189	7	190	8
rect	189	10	190	11
rect	189	13	190	14
rect	189	16	190	17
rect	189	19	190	20
rect	189	22	190	23
rect	189	25	190	26
rect	189	28	190	29
rect	189	31	190	32
rect	189	34	190	35
rect	189	37	190	38
rect	189	40	190	41
rect	189	43	190	44
rect	189	46	190	47
rect	189	49	190	50
rect	189	52	190	53
rect	189	55	190	56
rect	189	58	190	59
rect	189	61	190	62
rect	189	64	190	65
rect	189	67	190	68
rect	189	70	190	71
rect	189	73	190	74
rect	189	76	190	77
rect	189	79	190	80
rect	189	82	190	83
rect	189	85	190	86
rect	189	88	190	89
rect	189	91	190	92
rect	189	94	190	95
rect	189	97	190	98
rect	189	100	190	101
rect	189	103	190	104
rect	189	106	190	107
rect	189	109	190	110
rect	189	112	190	113
rect	189	115	190	116
rect	189	118	190	119
rect	189	121	190	122
rect	189	124	190	125
rect	189	127	190	128
rect	189	130	190	131
rect	189	133	190	134
rect	189	136	190	137
rect	189	139	190	140
rect	189	142	190	143
rect	189	145	190	146
rect	189	148	190	149
rect	189	151	190	152
rect	189	154	190	155
rect	189	157	190	158
rect	189	160	190	161
rect	189	163	190	164
rect	189	166	190	167
rect	189	169	190	170
rect	189	172	190	173
rect	189	175	190	176
rect	189	178	190	179
rect	189	181	190	182
rect	189	184	190	185
rect	189	187	190	188
rect	189	190	190	191
rect	189	193	190	194
rect	189	196	190	197
rect	189	199	190	200
rect	189	202	190	203
rect	189	205	190	206
rect	189	208	190	209
rect	189	211	190	212
rect	189	214	190	215
rect	189	217	190	218
rect	189	220	190	221
rect	189	223	190	224
rect	189	226	190	227
rect	189	229	190	230
rect	189	232	190	233
rect	189	235	190	236
rect	189	238	190	239
rect	189	241	190	242
rect	189	244	190	245
rect	189	247	190	248
rect	189	250	190	251
rect	189	253	190	254
rect	189	256	190	257
rect	189	259	190	260
rect	189	262	190	263
rect	189	265	190	266
rect	189	268	190	269
rect	189	271	190	272
rect	189	274	190	275
rect	189	277	190	278
rect	189	280	190	281
rect	189	283	190	284
rect	189	286	190	287
rect	189	289	190	290
rect	189	292	190	293
rect	189	295	190	296
rect	189	298	190	299
rect	189	301	190	302
rect	189	307	190	308
rect	189	310	190	311
rect	189	313	190	314
rect	189	316	190	317
rect	189	322	190	323
rect	189	325	190	326
rect	189	331	190	332
rect	189	334	190	335
rect	189	346	190	347
rect	189	349	190	350
rect	189	355	190	356
rect	189	358	190	359
rect	189	364	190	365
rect	190	7	191	8
rect	190	10	191	11
rect	190	13	191	14
rect	190	16	191	17
rect	190	19	191	20
rect	190	22	191	23
rect	190	25	191	26
rect	190	28	191	29
rect	190	31	191	32
rect	190	34	191	35
rect	190	37	191	38
rect	190	40	191	41
rect	190	43	191	44
rect	190	46	191	47
rect	190	49	191	50
rect	190	52	191	53
rect	190	55	191	56
rect	190	58	191	59
rect	190	61	191	62
rect	190	64	191	65
rect	190	67	191	68
rect	190	70	191	71
rect	190	73	191	74
rect	190	76	191	77
rect	190	79	191	80
rect	190	82	191	83
rect	190	85	191	86
rect	190	88	191	89
rect	190	91	191	92
rect	190	94	191	95
rect	190	97	191	98
rect	190	100	191	101
rect	190	103	191	104
rect	190	106	191	107
rect	190	109	191	110
rect	190	112	191	113
rect	190	115	191	116
rect	190	118	191	119
rect	190	121	191	122
rect	190	124	191	125
rect	190	127	191	128
rect	190	130	191	131
rect	190	133	191	134
rect	190	136	191	137
rect	190	139	191	140
rect	190	142	191	143
rect	190	145	191	146
rect	190	148	191	149
rect	190	151	191	152
rect	190	154	191	155
rect	190	157	191	158
rect	190	160	191	161
rect	190	163	191	164
rect	190	166	191	167
rect	190	169	191	170
rect	190	172	191	173
rect	190	175	191	176
rect	190	178	191	179
rect	190	181	191	182
rect	190	184	191	185
rect	190	187	191	188
rect	190	190	191	191
rect	190	193	191	194
rect	190	196	191	197
rect	190	199	191	200
rect	190	202	191	203
rect	190	205	191	206
rect	190	208	191	209
rect	190	211	191	212
rect	190	214	191	215
rect	190	217	191	218
rect	190	220	191	221
rect	190	223	191	224
rect	190	226	191	227
rect	190	229	191	230
rect	190	232	191	233
rect	190	235	191	236
rect	190	238	191	239
rect	190	241	191	242
rect	190	244	191	245
rect	190	247	191	248
rect	190	250	191	251
rect	190	253	191	254
rect	190	256	191	257
rect	190	259	191	260
rect	190	262	191	263
rect	190	265	191	266
rect	190	268	191	269
rect	190	271	191	272
rect	190	274	191	275
rect	190	277	191	278
rect	190	280	191	281
rect	190	283	191	284
rect	190	286	191	287
rect	190	289	191	290
rect	190	292	191	293
rect	190	295	191	296
rect	190	298	191	299
rect	190	301	191	302
rect	190	307	191	308
rect	190	310	191	311
rect	190	313	191	314
rect	190	316	191	317
rect	190	322	191	323
rect	190	325	191	326
rect	190	331	191	332
rect	190	334	191	335
rect	190	346	191	347
rect	190	349	191	350
rect	190	355	191	356
rect	190	358	191	359
rect	190	364	191	365
rect	191	4	192	5
rect	191	7	192	8
rect	191	10	192	11
rect	191	13	192	14
rect	191	16	192	17
rect	191	19	192	20
rect	191	22	192	23
rect	191	25	192	26
rect	191	28	192	29
rect	191	31	192	32
rect	191	34	192	35
rect	191	37	192	38
rect	191	40	192	41
rect	191	43	192	44
rect	191	46	192	47
rect	191	49	192	50
rect	191	52	192	53
rect	191	55	192	56
rect	191	58	192	59
rect	191	61	192	62
rect	191	64	192	65
rect	191	67	192	68
rect	191	70	192	71
rect	191	73	192	74
rect	191	76	192	77
rect	191	79	192	80
rect	191	82	192	83
rect	191	85	192	86
rect	191	88	192	89
rect	191	91	192	92
rect	191	94	192	95
rect	191	97	192	98
rect	191	100	192	101
rect	191	103	192	104
rect	191	106	192	107
rect	191	109	192	110
rect	191	112	192	113
rect	191	115	192	116
rect	191	118	192	119
rect	191	121	192	122
rect	191	124	192	125
rect	191	127	192	128
rect	191	130	192	131
rect	191	133	192	134
rect	191	136	192	137
rect	191	139	192	140
rect	191	142	192	143
rect	191	145	192	146
rect	191	148	192	149
rect	191	151	192	152
rect	191	154	192	155
rect	191	157	192	158
rect	191	160	192	161
rect	191	163	192	164
rect	191	166	192	167
rect	191	169	192	170
rect	191	172	192	173
rect	191	175	192	176
rect	191	178	192	179
rect	191	181	192	182
rect	191	184	192	185
rect	191	187	192	188
rect	191	190	192	191
rect	191	193	192	194
rect	191	196	192	197
rect	191	199	192	200
rect	191	202	192	203
rect	191	205	192	206
rect	191	208	192	209
rect	191	211	192	212
rect	191	214	192	215
rect	191	217	192	218
rect	191	220	192	221
rect	191	223	192	224
rect	191	226	192	227
rect	191	229	192	230
rect	191	232	192	233
rect	191	235	192	236
rect	191	238	192	239
rect	191	241	192	242
rect	191	244	192	245
rect	191	247	192	248
rect	191	250	192	251
rect	191	253	192	254
rect	191	256	192	257
rect	191	259	192	260
rect	191	262	192	263
rect	191	265	192	266
rect	191	268	192	269
rect	191	271	192	272
rect	191	274	192	275
rect	191	277	192	278
rect	191	280	192	281
rect	191	283	192	284
rect	191	286	192	287
rect	191	289	192	290
rect	191	292	192	293
rect	191	295	192	296
rect	191	298	192	299
rect	191	301	192	302
rect	191	307	192	308
rect	191	310	192	311
rect	191	313	192	314
rect	191	316	192	317
rect	191	322	192	323
rect	191	325	192	326
rect	191	331	192	332
rect	191	334	192	335
rect	191	346	192	347
rect	191	349	192	350
rect	191	355	192	356
rect	191	358	192	359
rect	191	364	192	365
rect	191	367	192	368
rect	192	4	193	5
rect	192	7	193	8
rect	192	10	193	11
rect	192	13	193	14
rect	192	16	193	17
rect	192	19	193	20
rect	192	22	193	23
rect	192	25	193	26
rect	192	28	193	29
rect	192	31	193	32
rect	192	34	193	35
rect	192	37	193	38
rect	192	40	193	41
rect	192	43	193	44
rect	192	46	193	47
rect	192	49	193	50
rect	192	52	193	53
rect	192	55	193	56
rect	192	58	193	59
rect	192	61	193	62
rect	192	64	193	65
rect	192	67	193	68
rect	192	70	193	71
rect	192	73	193	74
rect	192	76	193	77
rect	192	79	193	80
rect	192	82	193	83
rect	192	85	193	86
rect	192	88	193	89
rect	192	91	193	92
rect	192	94	193	95
rect	192	97	193	98
rect	192	100	193	101
rect	192	103	193	104
rect	192	106	193	107
rect	192	109	193	110
rect	192	112	193	113
rect	192	115	193	116
rect	192	118	193	119
rect	192	121	193	122
rect	192	124	193	125
rect	192	127	193	128
rect	192	130	193	131
rect	192	133	193	134
rect	192	136	193	137
rect	192	139	193	140
rect	192	142	193	143
rect	192	145	193	146
rect	192	148	193	149
rect	192	151	193	152
rect	192	154	193	155
rect	192	157	193	158
rect	192	160	193	161
rect	192	163	193	164
rect	192	166	193	167
rect	192	169	193	170
rect	192	172	193	173
rect	192	175	193	176
rect	192	178	193	179
rect	192	181	193	182
rect	192	184	193	185
rect	192	187	193	188
rect	192	190	193	191
rect	192	193	193	194
rect	192	196	193	197
rect	192	199	193	200
rect	192	202	193	203
rect	192	205	193	206
rect	192	208	193	209
rect	192	211	193	212
rect	192	214	193	215
rect	192	217	193	218
rect	192	220	193	221
rect	192	223	193	224
rect	192	226	193	227
rect	192	229	193	230
rect	192	232	193	233
rect	192	235	193	236
rect	192	238	193	239
rect	192	241	193	242
rect	192	244	193	245
rect	192	247	193	248
rect	192	250	193	251
rect	192	253	193	254
rect	192	256	193	257
rect	192	259	193	260
rect	192	265	193	266
rect	192	268	193	269
rect	192	271	193	272
rect	192	274	193	275
rect	192	277	193	278
rect	192	280	193	281
rect	192	283	193	284
rect	192	286	193	287
rect	192	289	193	290
rect	192	292	193	293
rect	192	295	193	296
rect	192	298	193	299
rect	192	301	193	302
rect	192	307	193	308
rect	192	310	193	311
rect	192	313	193	314
rect	192	316	193	317
rect	192	331	193	332
rect	192	334	193	335
rect	192	346	193	347
rect	193	4	194	5
rect	193	7	194	8
rect	193	10	194	11
rect	193	13	194	14
rect	193	16	194	17
rect	193	19	194	20
rect	193	22	194	23
rect	193	25	194	26
rect	193	28	194	29
rect	193	31	194	32
rect	193	34	194	35
rect	193	37	194	38
rect	193	40	194	41
rect	193	43	194	44
rect	193	46	194	47
rect	193	49	194	50
rect	193	52	194	53
rect	193	55	194	56
rect	193	58	194	59
rect	193	61	194	62
rect	193	64	194	65
rect	193	67	194	68
rect	193	70	194	71
rect	193	73	194	74
rect	193	76	194	77
rect	193	79	194	80
rect	193	82	194	83
rect	193	85	194	86
rect	193	88	194	89
rect	193	91	194	92
rect	193	94	194	95
rect	193	97	194	98
rect	193	100	194	101
rect	193	103	194	104
rect	193	106	194	107
rect	193	109	194	110
rect	193	112	194	113
rect	193	115	194	116
rect	193	118	194	119
rect	193	121	194	122
rect	193	124	194	125
rect	193	127	194	128
rect	193	130	194	131
rect	193	133	194	134
rect	193	136	194	137
rect	193	139	194	140
rect	193	142	194	143
rect	193	145	194	146
rect	193	148	194	149
rect	193	151	194	152
rect	193	154	194	155
rect	193	157	194	158
rect	193	160	194	161
rect	193	163	194	164
rect	193	166	194	167
rect	193	169	194	170
rect	193	172	194	173
rect	193	175	194	176
rect	193	178	194	179
rect	193	181	194	182
rect	193	184	194	185
rect	193	187	194	188
rect	193	190	194	191
rect	193	193	194	194
rect	193	196	194	197
rect	193	199	194	200
rect	193	202	194	203
rect	193	205	194	206
rect	193	208	194	209
rect	193	211	194	212
rect	193	214	194	215
rect	193	217	194	218
rect	193	220	194	221
rect	193	223	194	224
rect	193	226	194	227
rect	193	229	194	230
rect	193	232	194	233
rect	193	235	194	236
rect	193	238	194	239
rect	193	241	194	242
rect	193	244	194	245
rect	193	247	194	248
rect	193	250	194	251
rect	193	253	194	254
rect	193	256	194	257
rect	193	259	194	260
rect	193	265	194	266
rect	193	268	194	269
rect	193	271	194	272
rect	193	274	194	275
rect	193	277	194	278
rect	193	280	194	281
rect	193	283	194	284
rect	193	286	194	287
rect	193	289	194	290
rect	193	292	194	293
rect	193	295	194	296
rect	193	298	194	299
rect	193	301	194	302
rect	193	307	194	308
rect	193	310	194	311
rect	193	313	194	314
rect	193	316	194	317
rect	193	331	194	332
rect	193	334	194	335
rect	193	346	194	347
rect	194	4	195	5
rect	194	7	195	8
rect	194	10	195	11
rect	194	13	195	14
rect	194	16	195	17
rect	194	19	195	20
rect	194	22	195	23
rect	194	25	195	26
rect	194	28	195	29
rect	194	31	195	32
rect	194	34	195	35
rect	194	37	195	38
rect	194	40	195	41
rect	194	43	195	44
rect	194	46	195	47
rect	194	49	195	50
rect	194	52	195	53
rect	194	55	195	56
rect	194	58	195	59
rect	194	61	195	62
rect	194	64	195	65
rect	194	67	195	68
rect	194	70	195	71
rect	194	73	195	74
rect	194	76	195	77
rect	194	79	195	80
rect	194	82	195	83
rect	194	85	195	86
rect	194	88	195	89
rect	194	91	195	92
rect	194	94	195	95
rect	194	97	195	98
rect	194	100	195	101
rect	194	103	195	104
rect	194	106	195	107
rect	194	109	195	110
rect	194	112	195	113
rect	194	115	195	116
rect	194	118	195	119
rect	194	121	195	122
rect	194	124	195	125
rect	194	127	195	128
rect	194	130	195	131
rect	194	133	195	134
rect	194	136	195	137
rect	194	139	195	140
rect	194	142	195	143
rect	194	145	195	146
rect	194	148	195	149
rect	194	151	195	152
rect	194	154	195	155
rect	194	157	195	158
rect	194	160	195	161
rect	194	163	195	164
rect	194	166	195	167
rect	194	169	195	170
rect	194	172	195	173
rect	194	175	195	176
rect	194	178	195	179
rect	194	181	195	182
rect	194	184	195	185
rect	194	187	195	188
rect	194	190	195	191
rect	194	193	195	194
rect	194	196	195	197
rect	194	199	195	200
rect	194	202	195	203
rect	194	205	195	206
rect	194	208	195	209
rect	194	211	195	212
rect	194	214	195	215
rect	194	217	195	218
rect	194	220	195	221
rect	194	223	195	224
rect	194	226	195	227
rect	194	229	195	230
rect	194	232	195	233
rect	194	235	195	236
rect	194	238	195	239
rect	194	241	195	242
rect	194	244	195	245
rect	194	247	195	248
rect	194	250	195	251
rect	194	253	195	254
rect	194	256	195	257
rect	194	259	195	260
rect	194	265	195	266
rect	194	268	195	269
rect	194	271	195	272
rect	194	274	195	275
rect	194	277	195	278
rect	194	280	195	281
rect	194	283	195	284
rect	194	286	195	287
rect	194	289	195	290
rect	194	292	195	293
rect	194	295	195	296
rect	194	298	195	299
rect	194	301	195	302
rect	194	307	195	308
rect	194	310	195	311
rect	194	313	195	314
rect	194	316	195	317
rect	194	331	195	332
rect	194	334	195	335
rect	194	346	195	347
rect	195	4	196	5
rect	195	7	196	8
rect	195	10	196	11
rect	195	13	196	14
rect	195	16	196	17
rect	195	19	196	20
rect	195	22	196	23
rect	195	25	196	26
rect	195	28	196	29
rect	195	31	196	32
rect	195	34	196	35
rect	195	37	196	38
rect	195	40	196	41
rect	195	43	196	44
rect	195	46	196	47
rect	195	49	196	50
rect	195	52	196	53
rect	195	55	196	56
rect	195	58	196	59
rect	195	61	196	62
rect	195	64	196	65
rect	195	67	196	68
rect	195	70	196	71
rect	195	73	196	74
rect	195	76	196	77
rect	195	79	196	80
rect	195	82	196	83
rect	195	85	196	86
rect	195	88	196	89
rect	195	91	196	92
rect	195	94	196	95
rect	195	97	196	98
rect	195	100	196	101
rect	195	103	196	104
rect	195	106	196	107
rect	195	109	196	110
rect	195	112	196	113
rect	195	115	196	116
rect	195	118	196	119
rect	195	121	196	122
rect	195	124	196	125
rect	195	127	196	128
rect	195	130	196	131
rect	195	133	196	134
rect	195	136	196	137
rect	195	139	196	140
rect	195	142	196	143
rect	195	145	196	146
rect	195	148	196	149
rect	195	151	196	152
rect	195	154	196	155
rect	195	157	196	158
rect	195	160	196	161
rect	195	163	196	164
rect	195	166	196	167
rect	195	169	196	170
rect	195	172	196	173
rect	195	175	196	176
rect	195	178	196	179
rect	195	181	196	182
rect	195	184	196	185
rect	195	187	196	188
rect	195	190	196	191
rect	195	193	196	194
rect	195	196	196	197
rect	195	199	196	200
rect	195	202	196	203
rect	195	205	196	206
rect	195	208	196	209
rect	195	211	196	212
rect	195	214	196	215
rect	195	217	196	218
rect	195	220	196	221
rect	195	223	196	224
rect	195	226	196	227
rect	195	229	196	230
rect	195	232	196	233
rect	195	235	196	236
rect	195	238	196	239
rect	195	241	196	242
rect	195	244	196	245
rect	195	247	196	248
rect	195	250	196	251
rect	195	253	196	254
rect	195	256	196	257
rect	195	259	196	260
rect	195	265	196	266
rect	195	268	196	269
rect	195	271	196	272
rect	195	274	196	275
rect	195	277	196	278
rect	195	280	196	281
rect	195	283	196	284
rect	195	286	196	287
rect	195	289	196	290
rect	195	292	196	293
rect	195	295	196	296
rect	195	298	196	299
rect	195	301	196	302
rect	195	307	196	308
rect	195	310	196	311
rect	195	313	196	314
rect	195	316	196	317
rect	195	331	196	332
rect	195	334	196	335
rect	195	346	196	347
rect	196	4	197	5
rect	196	7	197	8
rect	196	10	197	11
rect	196	13	197	14
rect	196	16	197	17
rect	196	19	197	20
rect	196	22	197	23
rect	196	25	197	26
rect	196	28	197	29
rect	196	31	197	32
rect	196	34	197	35
rect	196	37	197	38
rect	196	40	197	41
rect	196	43	197	44
rect	196	46	197	47
rect	196	49	197	50
rect	196	52	197	53
rect	196	55	197	56
rect	196	58	197	59
rect	196	61	197	62
rect	196	64	197	65
rect	196	67	197	68
rect	196	70	197	71
rect	196	73	197	74
rect	196	76	197	77
rect	196	79	197	80
rect	196	82	197	83
rect	196	85	197	86
rect	196	88	197	89
rect	196	91	197	92
rect	196	94	197	95
rect	196	97	197	98
rect	196	100	197	101
rect	196	103	197	104
rect	196	106	197	107
rect	196	109	197	110
rect	196	112	197	113
rect	196	115	197	116
rect	196	118	197	119
rect	196	121	197	122
rect	196	124	197	125
rect	196	127	197	128
rect	196	130	197	131
rect	196	133	197	134
rect	196	136	197	137
rect	196	139	197	140
rect	196	142	197	143
rect	196	145	197	146
rect	196	148	197	149
rect	196	151	197	152
rect	196	154	197	155
rect	196	157	197	158
rect	196	160	197	161
rect	196	163	197	164
rect	196	166	197	167
rect	196	169	197	170
rect	196	172	197	173
rect	196	175	197	176
rect	196	178	197	179
rect	196	181	197	182
rect	196	184	197	185
rect	196	187	197	188
rect	196	190	197	191
rect	196	193	197	194
rect	196	196	197	197
rect	196	199	197	200
rect	196	202	197	203
rect	196	205	197	206
rect	196	208	197	209
rect	196	211	197	212
rect	196	214	197	215
rect	196	217	197	218
rect	196	220	197	221
rect	196	223	197	224
rect	196	226	197	227
rect	196	229	197	230
rect	196	232	197	233
rect	196	235	197	236
rect	196	238	197	239
rect	196	241	197	242
rect	196	244	197	245
rect	196	247	197	248
rect	196	250	197	251
rect	196	253	197	254
rect	196	256	197	257
rect	196	259	197	260
rect	196	265	197	266
rect	196	268	197	269
rect	196	271	197	272
rect	196	274	197	275
rect	196	277	197	278
rect	196	280	197	281
rect	196	283	197	284
rect	196	286	197	287
rect	196	289	197	290
rect	196	292	197	293
rect	196	295	197	296
rect	196	298	197	299
rect	196	301	197	302
rect	196	307	197	308
rect	196	310	197	311
rect	196	313	197	314
rect	196	316	197	317
rect	196	331	197	332
rect	196	334	197	335
rect	196	346	197	347
rect	197	4	198	5
rect	197	7	198	8
rect	197	10	198	11
rect	197	13	198	14
rect	197	16	198	17
rect	197	19	198	20
rect	197	22	198	23
rect	197	25	198	26
rect	197	28	198	29
rect	197	31	198	32
rect	197	34	198	35
rect	197	37	198	38
rect	197	40	198	41
rect	197	43	198	44
rect	197	46	198	47
rect	197	49	198	50
rect	197	52	198	53
rect	197	55	198	56
rect	197	58	198	59
rect	197	61	198	62
rect	197	64	198	65
rect	197	67	198	68
rect	197	70	198	71
rect	197	73	198	74
rect	197	76	198	77
rect	197	79	198	80
rect	197	82	198	83
rect	197	85	198	86
rect	197	88	198	89
rect	197	91	198	92
rect	197	94	198	95
rect	197	97	198	98
rect	197	100	198	101
rect	197	103	198	104
rect	197	106	198	107
rect	197	109	198	110
rect	197	112	198	113
rect	197	115	198	116
rect	197	118	198	119
rect	197	121	198	122
rect	197	124	198	125
rect	197	127	198	128
rect	197	130	198	131
rect	197	133	198	134
rect	197	136	198	137
rect	197	139	198	140
rect	197	142	198	143
rect	197	145	198	146
rect	197	148	198	149
rect	197	151	198	152
rect	197	154	198	155
rect	197	157	198	158
rect	197	160	198	161
rect	197	163	198	164
rect	197	166	198	167
rect	197	169	198	170
rect	197	172	198	173
rect	197	175	198	176
rect	197	178	198	179
rect	197	181	198	182
rect	197	184	198	185
rect	197	187	198	188
rect	197	190	198	191
rect	197	193	198	194
rect	197	196	198	197
rect	197	199	198	200
rect	197	202	198	203
rect	197	205	198	206
rect	197	208	198	209
rect	197	211	198	212
rect	197	214	198	215
rect	197	217	198	218
rect	197	220	198	221
rect	197	223	198	224
rect	197	226	198	227
rect	197	229	198	230
rect	197	232	198	233
rect	197	235	198	236
rect	197	238	198	239
rect	197	241	198	242
rect	197	244	198	245
rect	197	247	198	248
rect	197	250	198	251
rect	197	253	198	254
rect	197	256	198	257
rect	197	259	198	260
rect	197	265	198	266
rect	197	268	198	269
rect	197	271	198	272
rect	197	274	198	275
rect	197	277	198	278
rect	197	280	198	281
rect	197	283	198	284
rect	197	286	198	287
rect	197	289	198	290
rect	197	292	198	293
rect	197	295	198	296
rect	197	298	198	299
rect	197	301	198	302
rect	197	307	198	308
rect	197	310	198	311
rect	197	313	198	314
rect	197	316	198	317
rect	197	331	198	332
rect	197	334	198	335
rect	197	346	198	347
rect	198	4	199	5
rect	198	7	199	8
rect	198	10	199	11
rect	198	13	199	14
rect	198	16	199	17
rect	198	19	199	20
rect	198	22	199	23
rect	198	25	199	26
rect	198	28	199	29
rect	198	31	199	32
rect	198	34	199	35
rect	198	37	199	38
rect	198	40	199	41
rect	198	43	199	44
rect	198	46	199	47
rect	198	49	199	50
rect	198	52	199	53
rect	198	55	199	56
rect	198	58	199	59
rect	198	61	199	62
rect	198	64	199	65
rect	198	67	199	68
rect	198	70	199	71
rect	198	73	199	74
rect	198	76	199	77
rect	198	79	199	80
rect	198	82	199	83
rect	198	85	199	86
rect	198	88	199	89
rect	198	91	199	92
rect	198	94	199	95
rect	198	97	199	98
rect	198	100	199	101
rect	198	103	199	104
rect	198	106	199	107
rect	198	109	199	110
rect	198	112	199	113
rect	198	115	199	116
rect	198	118	199	119
rect	198	121	199	122
rect	198	124	199	125
rect	198	127	199	128
rect	198	130	199	131
rect	198	133	199	134
rect	198	136	199	137
rect	198	139	199	140
rect	198	142	199	143
rect	198	145	199	146
rect	198	148	199	149
rect	198	151	199	152
rect	198	154	199	155
rect	198	157	199	158
rect	198	160	199	161
rect	198	163	199	164
rect	198	166	199	167
rect	198	169	199	170
rect	198	172	199	173
rect	198	175	199	176
rect	198	178	199	179
rect	198	181	199	182
rect	198	184	199	185
rect	198	187	199	188
rect	198	190	199	191
rect	198	193	199	194
rect	198	196	199	197
rect	198	199	199	200
rect	198	202	199	203
rect	198	205	199	206
rect	198	208	199	209
rect	198	211	199	212
rect	198	214	199	215
rect	198	217	199	218
rect	198	220	199	221
rect	198	223	199	224
rect	198	226	199	227
rect	198	229	199	230
rect	198	232	199	233
rect	198	235	199	236
rect	198	238	199	239
rect	198	241	199	242
rect	198	244	199	245
rect	198	247	199	248
rect	198	250	199	251
rect	198	253	199	254
rect	198	256	199	257
rect	198	259	199	260
rect	198	265	199	266
rect	198	268	199	269
rect	198	271	199	272
rect	198	274	199	275
rect	198	277	199	278
rect	198	280	199	281
rect	198	283	199	284
rect	198	286	199	287
rect	198	289	199	290
rect	198	292	199	293
rect	198	295	199	296
rect	198	298	199	299
rect	198	301	199	302
rect	198	307	199	308
rect	198	310	199	311
rect	198	313	199	314
rect	198	316	199	317
rect	198	331	199	332
rect	198	334	199	335
rect	198	346	199	347
rect	199	4	200	5
rect	199	7	200	8
rect	199	10	200	11
rect	199	13	200	14
rect	199	16	200	17
rect	199	19	200	20
rect	199	22	200	23
rect	199	25	200	26
rect	199	28	200	29
rect	199	31	200	32
rect	199	34	200	35
rect	199	37	200	38
rect	199	40	200	41
rect	199	43	200	44
rect	199	46	200	47
rect	199	49	200	50
rect	199	52	200	53
rect	199	55	200	56
rect	199	58	200	59
rect	199	61	200	62
rect	199	64	200	65
rect	199	67	200	68
rect	199	70	200	71
rect	199	73	200	74
rect	199	76	200	77
rect	199	79	200	80
rect	199	82	200	83
rect	199	85	200	86
rect	199	88	200	89
rect	199	91	200	92
rect	199	94	200	95
rect	199	97	200	98
rect	199	100	200	101
rect	199	103	200	104
rect	199	106	200	107
rect	199	109	200	110
rect	199	112	200	113
rect	199	115	200	116
rect	199	118	200	119
rect	199	121	200	122
rect	199	124	200	125
rect	199	127	200	128
rect	199	130	200	131
rect	199	133	200	134
rect	199	136	200	137
rect	199	139	200	140
rect	199	142	200	143
rect	199	145	200	146
rect	199	148	200	149
rect	199	151	200	152
rect	199	154	200	155
rect	199	157	200	158
rect	199	160	200	161
rect	199	163	200	164
rect	199	166	200	167
rect	199	169	200	170
rect	199	172	200	173
rect	199	175	200	176
rect	199	178	200	179
rect	199	181	200	182
rect	199	184	200	185
rect	199	187	200	188
rect	199	190	200	191
rect	199	193	200	194
rect	199	196	200	197
rect	199	199	200	200
rect	199	202	200	203
rect	199	205	200	206
rect	199	208	200	209
rect	199	211	200	212
rect	199	214	200	215
rect	199	217	200	218
rect	199	220	200	221
rect	199	223	200	224
rect	199	226	200	227
rect	199	229	200	230
rect	199	232	200	233
rect	199	235	200	236
rect	199	238	200	239
rect	199	241	200	242
rect	199	244	200	245
rect	199	247	200	248
rect	199	250	200	251
rect	199	253	200	254
rect	199	256	200	257
rect	199	259	200	260
rect	199	265	200	266
rect	199	268	200	269
rect	199	271	200	272
rect	199	274	200	275
rect	199	277	200	278
rect	199	280	200	281
rect	199	283	200	284
rect	199	286	200	287
rect	199	289	200	290
rect	199	292	200	293
rect	199	295	200	296
rect	199	298	200	299
rect	199	301	200	302
rect	199	307	200	308
rect	199	310	200	311
rect	199	313	200	314
rect	199	316	200	317
rect	199	331	200	332
rect	199	334	200	335
rect	199	346	200	347
rect	200	4	201	5
rect	200	7	201	8
rect	200	10	201	11
rect	200	13	201	14
rect	200	16	201	17
rect	200	19	201	20
rect	200	22	201	23
rect	200	25	201	26
rect	200	28	201	29
rect	200	31	201	32
rect	200	34	201	35
rect	200	37	201	38
rect	200	40	201	41
rect	200	43	201	44
rect	200	46	201	47
rect	200	49	201	50
rect	200	52	201	53
rect	200	55	201	56
rect	200	58	201	59
rect	200	61	201	62
rect	200	64	201	65
rect	200	67	201	68
rect	200	70	201	71
rect	200	73	201	74
rect	200	76	201	77
rect	200	79	201	80
rect	200	82	201	83
rect	200	85	201	86
rect	200	88	201	89
rect	200	91	201	92
rect	200	94	201	95
rect	200	97	201	98
rect	200	100	201	101
rect	200	103	201	104
rect	200	106	201	107
rect	200	109	201	110
rect	200	112	201	113
rect	200	115	201	116
rect	200	118	201	119
rect	200	121	201	122
rect	200	124	201	125
rect	200	127	201	128
rect	200	130	201	131
rect	200	133	201	134
rect	200	136	201	137
rect	200	139	201	140
rect	200	142	201	143
rect	200	145	201	146
rect	200	148	201	149
rect	200	151	201	152
rect	200	154	201	155
rect	200	157	201	158
rect	200	160	201	161
rect	200	163	201	164
rect	200	166	201	167
rect	200	169	201	170
rect	200	172	201	173
rect	200	175	201	176
rect	200	178	201	179
rect	200	181	201	182
rect	200	184	201	185
rect	200	187	201	188
rect	200	190	201	191
rect	200	193	201	194
rect	200	196	201	197
rect	200	199	201	200
rect	200	202	201	203
rect	200	205	201	206
rect	200	208	201	209
rect	200	211	201	212
rect	200	214	201	215
rect	200	217	201	218
rect	200	220	201	221
rect	200	223	201	224
rect	200	226	201	227
rect	200	229	201	230
rect	200	232	201	233
rect	200	235	201	236
rect	200	238	201	239
rect	200	241	201	242
rect	200	244	201	245
rect	200	247	201	248
rect	200	250	201	251
rect	200	253	201	254
rect	200	256	201	257
rect	200	259	201	260
rect	200	265	201	266
rect	200	268	201	269
rect	200	271	201	272
rect	200	274	201	275
rect	200	277	201	278
rect	200	280	201	281
rect	200	283	201	284
rect	200	286	201	287
rect	200	289	201	290
rect	200	292	201	293
rect	200	295	201	296
rect	200	298	201	299
rect	200	301	201	302
rect	200	304	201	305
rect	200	307	201	308
rect	200	310	201	311
rect	200	313	201	314
rect	200	316	201	317
rect	200	331	201	332
rect	200	334	201	335
rect	200	346	201	347
rect	201	4	202	5
rect	201	7	202	8
rect	201	10	202	11
rect	201	13	202	14
rect	201	16	202	17
rect	201	19	202	20
rect	201	22	202	23
rect	201	25	202	26
rect	201	28	202	29
rect	201	31	202	32
rect	201	34	202	35
rect	201	37	202	38
rect	201	40	202	41
rect	201	43	202	44
rect	201	46	202	47
rect	201	49	202	50
rect	201	52	202	53
rect	201	55	202	56
rect	201	58	202	59
rect	201	61	202	62
rect	201	64	202	65
rect	201	67	202	68
rect	201	70	202	71
rect	201	73	202	74
rect	201	76	202	77
rect	201	79	202	80
rect	201	82	202	83
rect	201	85	202	86
rect	201	88	202	89
rect	201	91	202	92
rect	201	94	202	95
rect	201	97	202	98
rect	201	100	202	101
rect	201	103	202	104
rect	201	106	202	107
rect	201	109	202	110
rect	201	112	202	113
rect	201	115	202	116
rect	201	118	202	119
rect	201	121	202	122
rect	201	124	202	125
rect	201	127	202	128
rect	201	130	202	131
rect	201	133	202	134
rect	201	136	202	137
rect	201	139	202	140
rect	201	142	202	143
rect	201	145	202	146
rect	201	148	202	149
rect	201	151	202	152
rect	201	154	202	155
rect	201	157	202	158
rect	201	160	202	161
rect	201	163	202	164
rect	201	166	202	167
rect	201	169	202	170
rect	201	172	202	173
rect	201	175	202	176
rect	201	178	202	179
rect	201	181	202	182
rect	201	184	202	185
rect	201	187	202	188
rect	201	190	202	191
rect	201	193	202	194
rect	201	196	202	197
rect	201	199	202	200
rect	201	202	202	203
rect	201	205	202	206
rect	201	208	202	209
rect	201	211	202	212
rect	201	214	202	215
rect	201	217	202	218
rect	201	220	202	221
rect	201	223	202	224
rect	201	226	202	227
rect	201	229	202	230
rect	201	232	202	233
rect	201	235	202	236
rect	201	238	202	239
rect	201	241	202	242
rect	201	244	202	245
rect	201	247	202	248
rect	201	250	202	251
rect	201	256	202	257
rect	201	259	202	260
rect	201	265	202	266
rect	201	268	202	269
rect	201	271	202	272
rect	201	274	202	275
rect	201	277	202	278
rect	201	280	202	281
rect	201	283	202	284
rect	201	286	202	287
rect	201	289	202	290
rect	201	292	202	293
rect	201	295	202	296
rect	201	298	202	299
rect	201	301	202	302
rect	201	304	202	305
rect	201	307	202	308
rect	201	310	202	311
rect	201	313	202	314
rect	201	316	202	317
rect	201	331	202	332
rect	201	334	202	335
rect	201	346	202	347
rect	202	4	203	5
rect	202	7	203	8
rect	202	10	203	11
rect	202	13	203	14
rect	202	16	203	17
rect	202	19	203	20
rect	202	22	203	23
rect	202	25	203	26
rect	202	28	203	29
rect	202	31	203	32
rect	202	34	203	35
rect	202	37	203	38
rect	202	40	203	41
rect	202	43	203	44
rect	202	46	203	47
rect	202	49	203	50
rect	202	52	203	53
rect	202	55	203	56
rect	202	58	203	59
rect	202	61	203	62
rect	202	64	203	65
rect	202	67	203	68
rect	202	70	203	71
rect	202	73	203	74
rect	202	76	203	77
rect	202	79	203	80
rect	202	82	203	83
rect	202	85	203	86
rect	202	88	203	89
rect	202	91	203	92
rect	202	94	203	95
rect	202	97	203	98
rect	202	100	203	101
rect	202	103	203	104
rect	202	106	203	107
rect	202	109	203	110
rect	202	112	203	113
rect	202	115	203	116
rect	202	118	203	119
rect	202	121	203	122
rect	202	124	203	125
rect	202	127	203	128
rect	202	130	203	131
rect	202	133	203	134
rect	202	136	203	137
rect	202	139	203	140
rect	202	142	203	143
rect	202	145	203	146
rect	202	148	203	149
rect	202	151	203	152
rect	202	154	203	155
rect	202	157	203	158
rect	202	160	203	161
rect	202	163	203	164
rect	202	166	203	167
rect	202	169	203	170
rect	202	172	203	173
rect	202	175	203	176
rect	202	178	203	179
rect	202	181	203	182
rect	202	184	203	185
rect	202	187	203	188
rect	202	190	203	191
rect	202	193	203	194
rect	202	196	203	197
rect	202	199	203	200
rect	202	202	203	203
rect	202	205	203	206
rect	202	208	203	209
rect	202	211	203	212
rect	202	214	203	215
rect	202	217	203	218
rect	202	220	203	221
rect	202	223	203	224
rect	202	226	203	227
rect	202	229	203	230
rect	202	232	203	233
rect	202	235	203	236
rect	202	238	203	239
rect	202	241	203	242
rect	202	244	203	245
rect	202	247	203	248
rect	202	250	203	251
rect	202	253	203	254
rect	202	256	203	257
rect	202	259	203	260
rect	202	265	203	266
rect	202	268	203	269
rect	202	271	203	272
rect	202	274	203	275
rect	202	277	203	278
rect	202	280	203	281
rect	202	283	203	284
rect	202	286	203	287
rect	202	289	203	290
rect	202	292	203	293
rect	202	295	203	296
rect	202	298	203	299
rect	202	301	203	302
rect	202	304	203	305
rect	202	307	203	308
rect	202	310	203	311
rect	202	313	203	314
rect	202	316	203	317
rect	202	331	203	332
rect	202	334	203	335
rect	202	343	203	344
rect	202	346	203	347
rect	203	4	204	5
rect	203	7	204	8
rect	203	10	204	11
rect	203	13	204	14
rect	203	16	204	17
rect	203	19	204	20
rect	203	22	204	23
rect	203	25	204	26
rect	203	28	204	29
rect	203	31	204	32
rect	203	34	204	35
rect	203	37	204	38
rect	203	40	204	41
rect	203	43	204	44
rect	203	46	204	47
rect	203	49	204	50
rect	203	52	204	53
rect	203	55	204	56
rect	203	58	204	59
rect	203	61	204	62
rect	203	64	204	65
rect	203	67	204	68
rect	203	70	204	71
rect	203	73	204	74
rect	203	76	204	77
rect	203	79	204	80
rect	203	82	204	83
rect	203	85	204	86
rect	203	88	204	89
rect	203	91	204	92
rect	203	94	204	95
rect	203	97	204	98
rect	203	103	204	104
rect	203	106	204	107
rect	203	109	204	110
rect	203	115	204	116
rect	203	118	204	119
rect	203	121	204	122
rect	203	124	204	125
rect	203	127	204	128
rect	203	130	204	131
rect	203	133	204	134
rect	203	136	204	137
rect	203	139	204	140
rect	203	142	204	143
rect	203	145	204	146
rect	203	148	204	149
rect	203	151	204	152
rect	203	154	204	155
rect	203	157	204	158
rect	203	160	204	161
rect	203	163	204	164
rect	203	166	204	167
rect	203	169	204	170
rect	203	172	204	173
rect	203	175	204	176
rect	203	178	204	179
rect	203	181	204	182
rect	203	184	204	185
rect	203	187	204	188
rect	203	193	204	194
rect	203	196	204	197
rect	203	199	204	200
rect	203	202	204	203
rect	203	205	204	206
rect	203	208	204	209
rect	203	211	204	212
rect	203	214	204	215
rect	203	217	204	218
rect	203	220	204	221
rect	203	223	204	224
rect	203	226	204	227
rect	203	229	204	230
rect	203	232	204	233
rect	203	235	204	236
rect	203	238	204	239
rect	203	241	204	242
rect	203	244	204	245
rect	203	247	204	248
rect	203	250	204	251
rect	203	253	204	254
rect	203	256	204	257
rect	203	259	204	260
rect	203	265	204	266
rect	203	268	204	269
rect	203	271	204	272
rect	203	274	204	275
rect	203	277	204	278
rect	203	280	204	281
rect	203	283	204	284
rect	203	286	204	287
rect	203	289	204	290
rect	203	292	204	293
rect	203	295	204	296
rect	203	298	204	299
rect	203	301	204	302
rect	203	304	204	305
rect	203	307	204	308
rect	203	310	204	311
rect	203	313	204	314
rect	203	316	204	317
rect	203	331	204	332
rect	203	334	204	335
rect	203	343	204	344
rect	204	7	205	8
rect	204	10	205	11
rect	204	13	205	14
rect	204	16	205	17
rect	204	19	205	20
rect	204	22	205	23
rect	204	25	205	26
rect	204	28	205	29
rect	204	31	205	32
rect	204	34	205	35
rect	204	37	205	38
rect	204	40	205	41
rect	204	43	205	44
rect	204	46	205	47
rect	204	49	205	50
rect	204	52	205	53
rect	204	55	205	56
rect	204	58	205	59
rect	204	61	205	62
rect	204	64	205	65
rect	204	67	205	68
rect	204	70	205	71
rect	204	73	205	74
rect	204	76	205	77
rect	204	79	205	80
rect	204	82	205	83
rect	204	85	205	86
rect	204	88	205	89
rect	204	91	205	92
rect	204	94	205	95
rect	204	97	205	98
rect	204	100	205	101
rect	204	103	205	104
rect	204	106	205	107
rect	204	109	205	110
rect	204	112	205	113
rect	204	115	205	116
rect	204	118	205	119
rect	204	121	205	122
rect	204	124	205	125
rect	204	127	205	128
rect	204	130	205	131
rect	204	133	205	134
rect	204	136	205	137
rect	204	139	205	140
rect	204	142	205	143
rect	204	145	205	146
rect	204	148	205	149
rect	204	151	205	152
rect	204	154	205	155
rect	204	157	205	158
rect	204	160	205	161
rect	204	163	205	164
rect	204	166	205	167
rect	204	169	205	170
rect	204	172	205	173
rect	204	175	205	176
rect	204	178	205	179
rect	204	181	205	182
rect	204	184	205	185
rect	204	187	205	188
rect	204	190	205	191
rect	204	193	205	194
rect	204	196	205	197
rect	204	199	205	200
rect	204	202	205	203
rect	204	205	205	206
rect	204	208	205	209
rect	204	211	205	212
rect	204	214	205	215
rect	204	217	205	218
rect	204	220	205	221
rect	204	223	205	224
rect	204	226	205	227
rect	204	229	205	230
rect	204	232	205	233
rect	204	235	205	236
rect	204	238	205	239
rect	204	241	205	242
rect	204	244	205	245
rect	204	247	205	248
rect	204	250	205	251
rect	204	253	205	254
rect	204	256	205	257
rect	204	259	205	260
rect	204	265	205	266
rect	204	268	205	269
rect	204	271	205	272
rect	204	274	205	275
rect	204	277	205	278
rect	204	280	205	281
rect	204	283	205	284
rect	204	286	205	287
rect	204	292	205	293
rect	204	295	205	296
rect	204	298	205	299
rect	204	301	205	302
rect	204	307	205	308
rect	204	310	205	311
rect	204	316	205	317
rect	204	331	205	332
rect	204	343	205	344
rect	204	346	205	347
rect	205	7	206	8
rect	205	10	206	11
rect	205	13	206	14
rect	205	16	206	17
rect	205	19	206	20
rect	205	22	206	23
rect	205	25	206	26
rect	205	28	206	29
rect	205	31	206	32
rect	205	34	206	35
rect	205	37	206	38
rect	205	40	206	41
rect	205	43	206	44
rect	205	46	206	47
rect	205	49	206	50
rect	205	52	206	53
rect	205	55	206	56
rect	205	58	206	59
rect	205	61	206	62
rect	205	64	206	65
rect	205	67	206	68
rect	205	70	206	71
rect	205	73	206	74
rect	205	76	206	77
rect	205	79	206	80
rect	205	82	206	83
rect	205	85	206	86
rect	205	88	206	89
rect	205	91	206	92
rect	205	94	206	95
rect	205	97	206	98
rect	205	100	206	101
rect	205	103	206	104
rect	205	106	206	107
rect	205	109	206	110
rect	205	112	206	113
rect	205	115	206	116
rect	205	118	206	119
rect	205	121	206	122
rect	205	124	206	125
rect	205	127	206	128
rect	205	130	206	131
rect	205	133	206	134
rect	205	136	206	137
rect	205	139	206	140
rect	205	142	206	143
rect	205	145	206	146
rect	205	148	206	149
rect	205	151	206	152
rect	205	154	206	155
rect	205	157	206	158
rect	205	160	206	161
rect	205	163	206	164
rect	205	166	206	167
rect	205	169	206	170
rect	205	172	206	173
rect	205	175	206	176
rect	205	178	206	179
rect	205	181	206	182
rect	205	184	206	185
rect	205	187	206	188
rect	205	190	206	191
rect	205	193	206	194
rect	205	196	206	197
rect	205	199	206	200
rect	205	202	206	203
rect	205	205	206	206
rect	205	208	206	209
rect	205	211	206	212
rect	205	214	206	215
rect	205	217	206	218
rect	205	220	206	221
rect	205	223	206	224
rect	205	226	206	227
rect	205	229	206	230
rect	205	232	206	233
rect	205	235	206	236
rect	205	238	206	239
rect	205	241	206	242
rect	205	244	206	245
rect	205	247	206	248
rect	205	250	206	251
rect	205	253	206	254
rect	205	256	206	257
rect	205	259	206	260
rect	205	265	206	266
rect	205	268	206	269
rect	205	271	206	272
rect	205	274	206	275
rect	205	277	206	278
rect	205	280	206	281
rect	205	283	206	284
rect	205	286	206	287
rect	205	292	206	293
rect	205	295	206	296
rect	205	298	206	299
rect	205	301	206	302
rect	205	310	206	311
rect	205	316	206	317
rect	205	331	206	332
rect	205	343	206	344
rect	205	346	206	347
rect	206	7	207	8
rect	206	10	207	11
rect	206	13	207	14
rect	206	16	207	17
rect	206	19	207	20
rect	206	22	207	23
rect	206	25	207	26
rect	206	28	207	29
rect	206	31	207	32
rect	206	34	207	35
rect	206	37	207	38
rect	206	40	207	41
rect	206	43	207	44
rect	206	46	207	47
rect	206	49	207	50
rect	206	52	207	53
rect	206	55	207	56
rect	206	58	207	59
rect	206	61	207	62
rect	206	64	207	65
rect	206	67	207	68
rect	206	70	207	71
rect	206	73	207	74
rect	206	76	207	77
rect	206	79	207	80
rect	206	82	207	83
rect	206	85	207	86
rect	206	88	207	89
rect	206	91	207	92
rect	206	94	207	95
rect	206	97	207	98
rect	206	100	207	101
rect	206	103	207	104
rect	206	106	207	107
rect	206	109	207	110
rect	206	112	207	113
rect	206	115	207	116
rect	206	118	207	119
rect	206	121	207	122
rect	206	124	207	125
rect	206	127	207	128
rect	206	130	207	131
rect	206	133	207	134
rect	206	136	207	137
rect	206	139	207	140
rect	206	142	207	143
rect	206	145	207	146
rect	206	148	207	149
rect	206	151	207	152
rect	206	154	207	155
rect	206	157	207	158
rect	206	160	207	161
rect	206	163	207	164
rect	206	166	207	167
rect	206	169	207	170
rect	206	172	207	173
rect	206	175	207	176
rect	206	178	207	179
rect	206	181	207	182
rect	206	184	207	185
rect	206	187	207	188
rect	206	190	207	191
rect	206	193	207	194
rect	206	196	207	197
rect	206	199	207	200
rect	206	202	207	203
rect	206	205	207	206
rect	206	208	207	209
rect	206	211	207	212
rect	206	214	207	215
rect	206	217	207	218
rect	206	220	207	221
rect	206	223	207	224
rect	206	226	207	227
rect	206	229	207	230
rect	206	232	207	233
rect	206	235	207	236
rect	206	238	207	239
rect	206	241	207	242
rect	206	244	207	245
rect	206	247	207	248
rect	206	250	207	251
rect	206	253	207	254
rect	206	256	207	257
rect	206	259	207	260
rect	206	265	207	266
rect	206	268	207	269
rect	206	271	207	272
rect	206	274	207	275
rect	206	277	207	278
rect	206	280	207	281
rect	206	283	207	284
rect	206	286	207	287
rect	206	292	207	293
rect	206	295	207	296
rect	206	298	207	299
rect	206	301	207	302
rect	206	307	207	308
rect	206	310	207	311
rect	206	316	207	317
rect	206	331	207	332
rect	206	343	207	344
rect	206	346	207	347
rect	207	7	208	8
rect	207	10	208	11
rect	207	13	208	14
rect	207	16	208	17
rect	207	19	208	20
rect	207	22	208	23
rect	207	25	208	26
rect	207	28	208	29
rect	207	31	208	32
rect	207	34	208	35
rect	207	37	208	38
rect	207	40	208	41
rect	207	43	208	44
rect	207	46	208	47
rect	207	49	208	50
rect	207	52	208	53
rect	207	55	208	56
rect	207	58	208	59
rect	207	61	208	62
rect	207	64	208	65
rect	207	67	208	68
rect	207	70	208	71
rect	207	73	208	74
rect	207	76	208	77
rect	207	79	208	80
rect	207	82	208	83
rect	207	85	208	86
rect	207	88	208	89
rect	207	91	208	92
rect	207	94	208	95
rect	207	97	208	98
rect	207	100	208	101
rect	207	103	208	104
rect	207	106	208	107
rect	207	109	208	110
rect	207	112	208	113
rect	207	115	208	116
rect	207	118	208	119
rect	207	121	208	122
rect	207	124	208	125
rect	207	127	208	128
rect	207	130	208	131
rect	207	133	208	134
rect	207	136	208	137
rect	207	139	208	140
rect	207	142	208	143
rect	207	145	208	146
rect	207	148	208	149
rect	207	151	208	152
rect	207	154	208	155
rect	207	157	208	158
rect	207	160	208	161
rect	207	163	208	164
rect	207	166	208	167
rect	207	169	208	170
rect	207	172	208	173
rect	207	175	208	176
rect	207	178	208	179
rect	207	181	208	182
rect	207	184	208	185
rect	207	187	208	188
rect	207	190	208	191
rect	207	193	208	194
rect	207	196	208	197
rect	207	199	208	200
rect	207	202	208	203
rect	207	205	208	206
rect	207	208	208	209
rect	207	211	208	212
rect	207	214	208	215
rect	207	217	208	218
rect	207	220	208	221
rect	207	223	208	224
rect	207	226	208	227
rect	207	229	208	230
rect	207	232	208	233
rect	207	235	208	236
rect	207	238	208	239
rect	207	241	208	242
rect	207	244	208	245
rect	207	247	208	248
rect	207	250	208	251
rect	207	253	208	254
rect	207	256	208	257
rect	207	259	208	260
rect	207	265	208	266
rect	207	268	208	269
rect	207	271	208	272
rect	207	274	208	275
rect	207	277	208	278
rect	207	280	208	281
rect	207	283	208	284
rect	207	286	208	287
rect	207	292	208	293
rect	207	295	208	296
rect	207	298	208	299
rect	207	301	208	302
rect	207	307	208	308
rect	207	310	208	311
rect	207	316	208	317
rect	207	331	208	332
rect	207	343	208	344
rect	207	346	208	347
rect	208	4	209	5
rect	208	7	209	8
rect	208	10	209	11
rect	208	13	209	14
rect	208	16	209	17
rect	208	19	209	20
rect	208	22	209	23
rect	208	25	209	26
rect	208	28	209	29
rect	208	31	209	32
rect	208	34	209	35
rect	208	37	209	38
rect	208	40	209	41
rect	208	43	209	44
rect	208	46	209	47
rect	208	49	209	50
rect	208	52	209	53
rect	208	55	209	56
rect	208	58	209	59
rect	208	61	209	62
rect	208	64	209	65
rect	208	67	209	68
rect	208	70	209	71
rect	208	73	209	74
rect	208	76	209	77
rect	208	79	209	80
rect	208	82	209	83
rect	208	85	209	86
rect	208	88	209	89
rect	208	91	209	92
rect	208	94	209	95
rect	208	97	209	98
rect	208	100	209	101
rect	208	103	209	104
rect	208	106	209	107
rect	208	109	209	110
rect	208	112	209	113
rect	208	115	209	116
rect	208	118	209	119
rect	208	121	209	122
rect	208	124	209	125
rect	208	127	209	128
rect	208	130	209	131
rect	208	133	209	134
rect	208	136	209	137
rect	208	139	209	140
rect	208	142	209	143
rect	208	145	209	146
rect	208	148	209	149
rect	208	151	209	152
rect	208	154	209	155
rect	208	157	209	158
rect	208	160	209	161
rect	208	163	209	164
rect	208	166	209	167
rect	208	169	209	170
rect	208	172	209	173
rect	208	175	209	176
rect	208	178	209	179
rect	208	181	209	182
rect	208	184	209	185
rect	208	187	209	188
rect	208	190	209	191
rect	208	193	209	194
rect	208	196	209	197
rect	208	199	209	200
rect	208	202	209	203
rect	208	205	209	206
rect	208	208	209	209
rect	208	211	209	212
rect	208	214	209	215
rect	208	217	209	218
rect	208	220	209	221
rect	208	223	209	224
rect	208	226	209	227
rect	208	229	209	230
rect	208	232	209	233
rect	208	235	209	236
rect	208	238	209	239
rect	208	241	209	242
rect	208	244	209	245
rect	208	247	209	248
rect	208	250	209	251
rect	208	253	209	254
rect	208	256	209	257
rect	208	259	209	260
rect	208	265	209	266
rect	208	268	209	269
rect	208	271	209	272
rect	208	274	209	275
rect	208	277	209	278
rect	208	280	209	281
rect	208	283	209	284
rect	208	286	209	287
rect	208	292	209	293
rect	208	295	209	296
rect	208	298	209	299
rect	208	301	209	302
rect	208	307	209	308
rect	208	310	209	311
rect	208	313	209	314
rect	208	316	209	317
rect	208	331	209	332
rect	208	343	209	344
rect	208	346	209	347
rect	209	7	210	8
rect	209	10	210	11
rect	209	13	210	14
rect	209	16	210	17
rect	209	19	210	20
rect	209	22	210	23
rect	209	25	210	26
rect	209	28	210	29
rect	209	31	210	32
rect	209	34	210	35
rect	209	37	210	38
rect	209	40	210	41
rect	209	43	210	44
rect	209	46	210	47
rect	209	49	210	50
rect	209	52	210	53
rect	209	55	210	56
rect	209	58	210	59
rect	209	61	210	62
rect	209	64	210	65
rect	209	67	210	68
rect	209	70	210	71
rect	209	73	210	74
rect	209	76	210	77
rect	209	79	210	80
rect	209	82	210	83
rect	209	85	210	86
rect	209	88	210	89
rect	209	91	210	92
rect	209	94	210	95
rect	209	97	210	98
rect	209	100	210	101
rect	209	103	210	104
rect	209	106	210	107
rect	209	109	210	110
rect	209	112	210	113
rect	209	115	210	116
rect	209	118	210	119
rect	209	121	210	122
rect	209	124	210	125
rect	209	127	210	128
rect	209	130	210	131
rect	209	133	210	134
rect	209	136	210	137
rect	209	139	210	140
rect	209	142	210	143
rect	209	145	210	146
rect	209	148	210	149
rect	209	151	210	152
rect	209	154	210	155
rect	209	157	210	158
rect	209	160	210	161
rect	209	163	210	164
rect	209	166	210	167
rect	209	169	210	170
rect	209	172	210	173
rect	209	175	210	176
rect	209	178	210	179
rect	209	181	210	182
rect	209	184	210	185
rect	209	187	210	188
rect	209	190	210	191
rect	209	193	210	194
rect	209	196	210	197
rect	209	199	210	200
rect	209	202	210	203
rect	209	205	210	206
rect	209	208	210	209
rect	209	211	210	212
rect	209	214	210	215
rect	209	217	210	218
rect	209	220	210	221
rect	209	223	210	224
rect	209	226	210	227
rect	209	229	210	230
rect	209	232	210	233
rect	209	235	210	236
rect	209	238	210	239
rect	209	241	210	242
rect	209	244	210	245
rect	209	247	210	248
rect	209	250	210	251
rect	209	256	210	257
rect	209	259	210	260
rect	209	265	210	266
rect	209	268	210	269
rect	209	271	210	272
rect	209	274	210	275
rect	209	277	210	278
rect	209	283	210	284
rect	209	286	210	287
rect	209	292	210	293
rect	209	307	210	308
rect	209	310	210	311
rect	209	316	210	317
rect	210	7	211	8
rect	210	10	211	11
rect	210	13	211	14
rect	210	16	211	17
rect	210	19	211	20
rect	210	22	211	23
rect	210	25	211	26
rect	210	28	211	29
rect	210	31	211	32
rect	210	34	211	35
rect	210	37	211	38
rect	210	40	211	41
rect	210	43	211	44
rect	210	46	211	47
rect	210	49	211	50
rect	210	52	211	53
rect	210	55	211	56
rect	210	58	211	59
rect	210	61	211	62
rect	210	64	211	65
rect	210	67	211	68
rect	210	70	211	71
rect	210	73	211	74
rect	210	76	211	77
rect	210	79	211	80
rect	210	82	211	83
rect	210	85	211	86
rect	210	88	211	89
rect	210	91	211	92
rect	210	94	211	95
rect	210	97	211	98
rect	210	100	211	101
rect	210	103	211	104
rect	210	106	211	107
rect	210	109	211	110
rect	210	112	211	113
rect	210	115	211	116
rect	210	118	211	119
rect	210	121	211	122
rect	210	124	211	125
rect	210	127	211	128
rect	210	130	211	131
rect	210	133	211	134
rect	210	136	211	137
rect	210	139	211	140
rect	210	142	211	143
rect	210	145	211	146
rect	210	148	211	149
rect	210	151	211	152
rect	210	154	211	155
rect	210	157	211	158
rect	210	160	211	161
rect	210	163	211	164
rect	210	166	211	167
rect	210	169	211	170
rect	210	172	211	173
rect	210	175	211	176
rect	210	178	211	179
rect	210	181	211	182
rect	210	184	211	185
rect	210	187	211	188
rect	210	190	211	191
rect	210	193	211	194
rect	210	196	211	197
rect	210	199	211	200
rect	210	202	211	203
rect	210	205	211	206
rect	210	208	211	209
rect	210	211	211	212
rect	210	214	211	215
rect	210	217	211	218
rect	210	220	211	221
rect	210	223	211	224
rect	210	226	211	227
rect	210	229	211	230
rect	210	232	211	233
rect	210	235	211	236
rect	210	238	211	239
rect	210	241	211	242
rect	210	244	211	245
rect	210	247	211	248
rect	210	250	211	251
rect	210	256	211	257
rect	210	259	211	260
rect	210	265	211	266
rect	210	268	211	269
rect	210	271	211	272
rect	210	274	211	275
rect	210	277	211	278
rect	210	283	211	284
rect	210	286	211	287
rect	210	292	211	293
rect	210	307	211	308
rect	210	310	211	311
rect	210	316	211	317
rect	211	7	212	8
rect	211	10	212	11
rect	211	13	212	14
rect	211	16	212	17
rect	211	19	212	20
rect	211	22	212	23
rect	211	25	212	26
rect	211	28	212	29
rect	211	31	212	32
rect	211	34	212	35
rect	211	37	212	38
rect	211	40	212	41
rect	211	43	212	44
rect	211	46	212	47
rect	211	49	212	50
rect	211	52	212	53
rect	211	55	212	56
rect	211	58	212	59
rect	211	61	212	62
rect	211	64	212	65
rect	211	67	212	68
rect	211	70	212	71
rect	211	73	212	74
rect	211	76	212	77
rect	211	79	212	80
rect	211	82	212	83
rect	211	85	212	86
rect	211	88	212	89
rect	211	91	212	92
rect	211	94	212	95
rect	211	97	212	98
rect	211	100	212	101
rect	211	103	212	104
rect	211	106	212	107
rect	211	109	212	110
rect	211	112	212	113
rect	211	115	212	116
rect	211	118	212	119
rect	211	121	212	122
rect	211	124	212	125
rect	211	127	212	128
rect	211	130	212	131
rect	211	133	212	134
rect	211	136	212	137
rect	211	139	212	140
rect	211	142	212	143
rect	211	145	212	146
rect	211	148	212	149
rect	211	151	212	152
rect	211	154	212	155
rect	211	157	212	158
rect	211	160	212	161
rect	211	163	212	164
rect	211	166	212	167
rect	211	169	212	170
rect	211	172	212	173
rect	211	175	212	176
rect	211	178	212	179
rect	211	181	212	182
rect	211	184	212	185
rect	211	187	212	188
rect	211	190	212	191
rect	211	193	212	194
rect	211	196	212	197
rect	211	199	212	200
rect	211	202	212	203
rect	211	205	212	206
rect	211	208	212	209
rect	211	211	212	212
rect	211	214	212	215
rect	211	217	212	218
rect	211	220	212	221
rect	211	223	212	224
rect	211	226	212	227
rect	211	229	212	230
rect	211	232	212	233
rect	211	235	212	236
rect	211	238	212	239
rect	211	241	212	242
rect	211	244	212	245
rect	211	247	212	248
rect	211	250	212	251
rect	211	256	212	257
rect	211	259	212	260
rect	211	265	212	266
rect	211	268	212	269
rect	211	271	212	272
rect	211	274	212	275
rect	211	277	212	278
rect	211	283	212	284
rect	211	286	212	287
rect	211	292	212	293
rect	211	307	212	308
rect	211	310	212	311
rect	211	316	212	317
rect	212	7	213	8
rect	212	10	213	11
rect	212	13	213	14
rect	212	16	213	17
rect	212	19	213	20
rect	212	22	213	23
rect	212	25	213	26
rect	212	28	213	29
rect	212	31	213	32
rect	212	34	213	35
rect	212	37	213	38
rect	212	40	213	41
rect	212	43	213	44
rect	212	46	213	47
rect	212	49	213	50
rect	212	52	213	53
rect	212	55	213	56
rect	212	58	213	59
rect	212	61	213	62
rect	212	64	213	65
rect	212	67	213	68
rect	212	70	213	71
rect	212	73	213	74
rect	212	76	213	77
rect	212	79	213	80
rect	212	82	213	83
rect	212	85	213	86
rect	212	88	213	89
rect	212	91	213	92
rect	212	94	213	95
rect	212	97	213	98
rect	212	100	213	101
rect	212	103	213	104
rect	212	106	213	107
rect	212	109	213	110
rect	212	112	213	113
rect	212	115	213	116
rect	212	118	213	119
rect	212	121	213	122
rect	212	124	213	125
rect	212	127	213	128
rect	212	130	213	131
rect	212	133	213	134
rect	212	136	213	137
rect	212	139	213	140
rect	212	142	213	143
rect	212	145	213	146
rect	212	148	213	149
rect	212	151	213	152
rect	212	154	213	155
rect	212	157	213	158
rect	212	160	213	161
rect	212	163	213	164
rect	212	166	213	167
rect	212	169	213	170
rect	212	172	213	173
rect	212	175	213	176
rect	212	178	213	179
rect	212	181	213	182
rect	212	184	213	185
rect	212	187	213	188
rect	212	190	213	191
rect	212	193	213	194
rect	212	196	213	197
rect	212	199	213	200
rect	212	202	213	203
rect	212	205	213	206
rect	212	208	213	209
rect	212	211	213	212
rect	212	214	213	215
rect	212	217	213	218
rect	212	220	213	221
rect	212	223	213	224
rect	212	226	213	227
rect	212	229	213	230
rect	212	232	213	233
rect	212	235	213	236
rect	212	238	213	239
rect	212	241	213	242
rect	212	244	213	245
rect	212	247	213	248
rect	212	250	213	251
rect	212	256	213	257
rect	212	259	213	260
rect	212	265	213	266
rect	212	268	213	269
rect	212	271	213	272
rect	212	274	213	275
rect	212	277	213	278
rect	212	283	213	284
rect	212	286	213	287
rect	212	292	213	293
rect	212	307	213	308
rect	212	310	213	311
rect	212	316	213	317
rect	213	7	214	8
rect	213	10	214	11
rect	213	13	214	14
rect	213	16	214	17
rect	213	19	214	20
rect	213	22	214	23
rect	213	25	214	26
rect	213	28	214	29
rect	213	31	214	32
rect	213	34	214	35
rect	213	37	214	38
rect	213	40	214	41
rect	213	43	214	44
rect	213	46	214	47
rect	213	49	214	50
rect	213	52	214	53
rect	213	55	214	56
rect	213	58	214	59
rect	213	61	214	62
rect	213	64	214	65
rect	213	67	214	68
rect	213	70	214	71
rect	213	73	214	74
rect	213	76	214	77
rect	213	79	214	80
rect	213	82	214	83
rect	213	85	214	86
rect	213	88	214	89
rect	213	91	214	92
rect	213	94	214	95
rect	213	97	214	98
rect	213	100	214	101
rect	213	103	214	104
rect	213	106	214	107
rect	213	109	214	110
rect	213	112	214	113
rect	213	115	214	116
rect	213	118	214	119
rect	213	121	214	122
rect	213	124	214	125
rect	213	127	214	128
rect	213	130	214	131
rect	213	133	214	134
rect	213	136	214	137
rect	213	139	214	140
rect	213	142	214	143
rect	213	145	214	146
rect	213	148	214	149
rect	213	151	214	152
rect	213	154	214	155
rect	213	157	214	158
rect	213	160	214	161
rect	213	163	214	164
rect	213	166	214	167
rect	213	169	214	170
rect	213	172	214	173
rect	213	175	214	176
rect	213	178	214	179
rect	213	181	214	182
rect	213	184	214	185
rect	213	187	214	188
rect	213	190	214	191
rect	213	193	214	194
rect	213	196	214	197
rect	213	199	214	200
rect	213	202	214	203
rect	213	205	214	206
rect	213	208	214	209
rect	213	211	214	212
rect	213	214	214	215
rect	213	217	214	218
rect	213	220	214	221
rect	213	223	214	224
rect	213	226	214	227
rect	213	229	214	230
rect	213	232	214	233
rect	213	235	214	236
rect	213	238	214	239
rect	213	241	214	242
rect	213	244	214	245
rect	213	247	214	248
rect	213	250	214	251
rect	213	256	214	257
rect	213	259	214	260
rect	213	265	214	266
rect	213	268	214	269
rect	213	271	214	272
rect	213	274	214	275
rect	213	277	214	278
rect	213	283	214	284
rect	213	286	214	287
rect	213	292	214	293
rect	213	307	214	308
rect	213	310	214	311
rect	213	316	214	317
rect	214	7	215	8
rect	214	10	215	11
rect	214	13	215	14
rect	214	16	215	17
rect	214	19	215	20
rect	214	22	215	23
rect	214	25	215	26
rect	214	28	215	29
rect	214	31	215	32
rect	214	34	215	35
rect	214	37	215	38
rect	214	40	215	41
rect	214	43	215	44
rect	214	46	215	47
rect	214	49	215	50
rect	214	52	215	53
rect	214	55	215	56
rect	214	58	215	59
rect	214	61	215	62
rect	214	64	215	65
rect	214	67	215	68
rect	214	70	215	71
rect	214	73	215	74
rect	214	76	215	77
rect	214	79	215	80
rect	214	82	215	83
rect	214	85	215	86
rect	214	88	215	89
rect	214	91	215	92
rect	214	94	215	95
rect	214	97	215	98
rect	214	100	215	101
rect	214	103	215	104
rect	214	106	215	107
rect	214	109	215	110
rect	214	112	215	113
rect	214	115	215	116
rect	214	118	215	119
rect	214	121	215	122
rect	214	124	215	125
rect	214	127	215	128
rect	214	130	215	131
rect	214	133	215	134
rect	214	136	215	137
rect	214	139	215	140
rect	214	142	215	143
rect	214	145	215	146
rect	214	148	215	149
rect	214	151	215	152
rect	214	154	215	155
rect	214	157	215	158
rect	214	160	215	161
rect	214	163	215	164
rect	214	166	215	167
rect	214	169	215	170
rect	214	172	215	173
rect	214	175	215	176
rect	214	178	215	179
rect	214	181	215	182
rect	214	184	215	185
rect	214	187	215	188
rect	214	190	215	191
rect	214	193	215	194
rect	214	196	215	197
rect	214	199	215	200
rect	214	202	215	203
rect	214	205	215	206
rect	214	208	215	209
rect	214	211	215	212
rect	214	214	215	215
rect	214	217	215	218
rect	214	220	215	221
rect	214	223	215	224
rect	214	226	215	227
rect	214	229	215	230
rect	214	232	215	233
rect	214	235	215	236
rect	214	238	215	239
rect	214	241	215	242
rect	214	244	215	245
rect	214	247	215	248
rect	214	250	215	251
rect	214	256	215	257
rect	214	259	215	260
rect	214	265	215	266
rect	214	268	215	269
rect	214	271	215	272
rect	214	274	215	275
rect	214	277	215	278
rect	214	283	215	284
rect	214	286	215	287
rect	214	292	215	293
rect	214	307	215	308
rect	214	310	215	311
rect	214	316	215	317
rect	215	7	216	8
rect	215	10	216	11
rect	215	13	216	14
rect	215	16	216	17
rect	215	19	216	20
rect	215	22	216	23
rect	215	25	216	26
rect	215	28	216	29
rect	215	31	216	32
rect	215	34	216	35
rect	215	37	216	38
rect	215	40	216	41
rect	215	43	216	44
rect	215	46	216	47
rect	215	49	216	50
rect	215	52	216	53
rect	215	55	216	56
rect	215	58	216	59
rect	215	61	216	62
rect	215	64	216	65
rect	215	67	216	68
rect	215	70	216	71
rect	215	73	216	74
rect	215	76	216	77
rect	215	79	216	80
rect	215	82	216	83
rect	215	85	216	86
rect	215	88	216	89
rect	215	91	216	92
rect	215	94	216	95
rect	215	97	216	98
rect	215	100	216	101
rect	215	103	216	104
rect	215	106	216	107
rect	215	109	216	110
rect	215	112	216	113
rect	215	115	216	116
rect	215	118	216	119
rect	215	121	216	122
rect	215	124	216	125
rect	215	127	216	128
rect	215	130	216	131
rect	215	133	216	134
rect	215	136	216	137
rect	215	139	216	140
rect	215	142	216	143
rect	215	145	216	146
rect	215	148	216	149
rect	215	151	216	152
rect	215	154	216	155
rect	215	157	216	158
rect	215	160	216	161
rect	215	163	216	164
rect	215	166	216	167
rect	215	169	216	170
rect	215	172	216	173
rect	215	175	216	176
rect	215	178	216	179
rect	215	181	216	182
rect	215	184	216	185
rect	215	187	216	188
rect	215	190	216	191
rect	215	193	216	194
rect	215	196	216	197
rect	215	199	216	200
rect	215	202	216	203
rect	215	205	216	206
rect	215	208	216	209
rect	215	211	216	212
rect	215	214	216	215
rect	215	217	216	218
rect	215	220	216	221
rect	215	223	216	224
rect	215	226	216	227
rect	215	229	216	230
rect	215	232	216	233
rect	215	235	216	236
rect	215	238	216	239
rect	215	241	216	242
rect	215	244	216	245
rect	215	247	216	248
rect	215	250	216	251
rect	215	256	216	257
rect	215	259	216	260
rect	215	265	216	266
rect	215	268	216	269
rect	215	271	216	272
rect	215	274	216	275
rect	215	277	216	278
rect	215	292	216	293
rect	215	307	216	308
rect	216	7	217	8
rect	216	10	217	11
rect	216	13	217	14
rect	216	16	217	17
rect	216	19	217	20
rect	216	22	217	23
rect	216	25	217	26
rect	216	28	217	29
rect	216	31	217	32
rect	216	34	217	35
rect	216	37	217	38
rect	216	40	217	41
rect	216	43	217	44
rect	216	46	217	47
rect	216	49	217	50
rect	216	52	217	53
rect	216	55	217	56
rect	216	58	217	59
rect	216	61	217	62
rect	216	64	217	65
rect	216	67	217	68
rect	216	70	217	71
rect	216	73	217	74
rect	216	76	217	77
rect	216	79	217	80
rect	216	82	217	83
rect	216	85	217	86
rect	216	88	217	89
rect	216	91	217	92
rect	216	94	217	95
rect	216	97	217	98
rect	216	100	217	101
rect	216	103	217	104
rect	216	106	217	107
rect	216	109	217	110
rect	216	112	217	113
rect	216	115	217	116
rect	216	118	217	119
rect	216	121	217	122
rect	216	124	217	125
rect	216	127	217	128
rect	216	130	217	131
rect	216	133	217	134
rect	216	136	217	137
rect	216	139	217	140
rect	216	142	217	143
rect	216	145	217	146
rect	216	148	217	149
rect	216	151	217	152
rect	216	154	217	155
rect	216	157	217	158
rect	216	160	217	161
rect	216	163	217	164
rect	216	166	217	167
rect	216	169	217	170
rect	216	172	217	173
rect	216	175	217	176
rect	216	178	217	179
rect	216	181	217	182
rect	216	184	217	185
rect	216	187	217	188
rect	216	190	217	191
rect	216	193	217	194
rect	216	196	217	197
rect	216	199	217	200
rect	216	202	217	203
rect	216	205	217	206
rect	216	211	217	212
rect	216	214	217	215
rect	216	217	217	218
rect	216	220	217	221
rect	216	223	217	224
rect	216	226	217	227
rect	216	229	217	230
rect	216	232	217	233
rect	216	235	217	236
rect	216	238	217	239
rect	216	241	217	242
rect	216	244	217	245
rect	216	247	217	248
rect	216	250	217	251
rect	216	256	217	257
rect	216	259	217	260
rect	216	265	217	266
rect	216	268	217	269
rect	216	271	217	272
rect	216	274	217	275
rect	216	277	217	278
rect	216	292	217	293
rect	216	307	217	308
rect	217	4	218	5
rect	217	7	218	8
rect	217	10	218	11
rect	217	13	218	14
rect	217	16	218	17
rect	217	19	218	20
rect	217	22	218	23
rect	217	25	218	26
rect	217	28	218	29
rect	217	31	218	32
rect	217	34	218	35
rect	217	37	218	38
rect	217	40	218	41
rect	217	43	218	44
rect	217	46	218	47
rect	217	49	218	50
rect	217	52	218	53
rect	217	55	218	56
rect	217	58	218	59
rect	217	61	218	62
rect	217	64	218	65
rect	217	67	218	68
rect	217	70	218	71
rect	217	73	218	74
rect	217	76	218	77
rect	217	79	218	80
rect	217	82	218	83
rect	217	85	218	86
rect	217	88	218	89
rect	217	91	218	92
rect	217	94	218	95
rect	217	97	218	98
rect	217	100	218	101
rect	217	103	218	104
rect	217	106	218	107
rect	217	109	218	110
rect	217	112	218	113
rect	217	115	218	116
rect	217	118	218	119
rect	217	121	218	122
rect	217	124	218	125
rect	217	127	218	128
rect	217	130	218	131
rect	217	133	218	134
rect	217	136	218	137
rect	217	139	218	140
rect	217	142	218	143
rect	217	145	218	146
rect	217	148	218	149
rect	217	151	218	152
rect	217	154	218	155
rect	217	157	218	158
rect	217	160	218	161
rect	217	163	218	164
rect	217	166	218	167
rect	217	169	218	170
rect	217	172	218	173
rect	217	175	218	176
rect	217	178	218	179
rect	217	181	218	182
rect	217	184	218	185
rect	217	187	218	188
rect	217	190	218	191
rect	217	193	218	194
rect	217	196	218	197
rect	217	199	218	200
rect	217	202	218	203
rect	217	205	218	206
rect	217	208	218	209
rect	217	211	218	212
rect	217	214	218	215
rect	217	217	218	218
rect	217	220	218	221
rect	217	223	218	224
rect	217	226	218	227
rect	217	229	218	230
rect	217	232	218	233
rect	217	235	218	236
rect	217	238	218	239
rect	217	241	218	242
rect	217	244	218	245
rect	217	247	218	248
rect	217	250	218	251
rect	217	256	218	257
rect	217	259	218	260
rect	217	265	218	266
rect	217	268	218	269
rect	217	271	218	272
rect	217	274	218	275
rect	217	277	218	278
rect	217	292	218	293
rect	217	307	218	308
rect	218	4	219	5
rect	218	10	219	11
rect	218	13	219	14
rect	218	16	219	17
rect	218	19	219	20
rect	218	22	219	23
rect	218	25	219	26
rect	218	28	219	29
rect	218	31	219	32
rect	218	34	219	35
rect	218	37	219	38
rect	218	40	219	41
rect	218	43	219	44
rect	218	46	219	47
rect	218	49	219	50
rect	218	52	219	53
rect	218	55	219	56
rect	218	58	219	59
rect	218	61	219	62
rect	218	64	219	65
rect	218	67	219	68
rect	218	70	219	71
rect	218	73	219	74
rect	218	76	219	77
rect	218	79	219	80
rect	218	82	219	83
rect	218	85	219	86
rect	218	88	219	89
rect	218	91	219	92
rect	218	94	219	95
rect	218	97	219	98
rect	218	100	219	101
rect	218	103	219	104
rect	218	109	219	110
rect	218	112	219	113
rect	218	115	219	116
rect	218	118	219	119
rect	218	121	219	122
rect	218	124	219	125
rect	218	127	219	128
rect	218	133	219	134
rect	218	136	219	137
rect	218	142	219	143
rect	218	145	219	146
rect	218	148	219	149
rect	218	151	219	152
rect	218	154	219	155
rect	218	157	219	158
rect	218	160	219	161
rect	218	163	219	164
rect	218	166	219	167
rect	218	169	219	170
rect	218	172	219	173
rect	218	175	219	176
rect	218	178	219	179
rect	218	181	219	182
rect	218	184	219	185
rect	218	187	219	188
rect	218	190	219	191
rect	218	193	219	194
rect	218	196	219	197
rect	218	199	219	200
rect	218	202	219	203
rect	218	205	219	206
rect	218	208	219	209
rect	218	211	219	212
rect	218	214	219	215
rect	218	217	219	218
rect	218	220	219	221
rect	218	223	219	224
rect	218	226	219	227
rect	218	229	219	230
rect	218	232	219	233
rect	218	235	219	236
rect	218	241	219	242
rect	218	244	219	245
rect	218	247	219	248
rect	218	250	219	251
rect	218	256	219	257
rect	218	259	219	260
rect	218	265	219	266
rect	218	268	219	269
rect	218	271	219	272
rect	218	274	219	275
rect	218	277	219	278
rect	218	292	219	293
rect	218	307	219	308
rect	219	1	220	2
rect	219	4	220	5
rect	219	7	220	8
rect	219	10	220	11
rect	219	13	220	14
rect	219	16	220	17
rect	219	19	220	20
rect	219	22	220	23
rect	219	25	220	26
rect	219	28	220	29
rect	219	31	220	32
rect	219	34	220	35
rect	219	37	220	38
rect	219	40	220	41
rect	219	43	220	44
rect	219	46	220	47
rect	219	49	220	50
rect	219	52	220	53
rect	219	55	220	56
rect	219	58	220	59
rect	219	61	220	62
rect	219	64	220	65
rect	219	67	220	68
rect	219	70	220	71
rect	219	73	220	74
rect	219	76	220	77
rect	219	79	220	80
rect	219	82	220	83
rect	219	85	220	86
rect	219	88	220	89
rect	219	91	220	92
rect	219	94	220	95
rect	219	97	220	98
rect	219	100	220	101
rect	219	103	220	104
rect	219	106	220	107
rect	219	109	220	110
rect	219	112	220	113
rect	219	115	220	116
rect	219	118	220	119
rect	219	121	220	122
rect	219	124	220	125
rect	219	127	220	128
rect	219	130	220	131
rect	219	133	220	134
rect	219	136	220	137
rect	219	139	220	140
rect	219	142	220	143
rect	219	145	220	146
rect	219	148	220	149
rect	219	151	220	152
rect	219	154	220	155
rect	219	157	220	158
rect	219	160	220	161
rect	219	163	220	164
rect	219	166	220	167
rect	219	169	220	170
rect	219	172	220	173
rect	219	175	220	176
rect	219	178	220	179
rect	219	181	220	182
rect	219	184	220	185
rect	219	187	220	188
rect	219	190	220	191
rect	219	193	220	194
rect	219	196	220	197
rect	219	199	220	200
rect	219	202	220	203
rect	219	205	220	206
rect	219	208	220	209
rect	219	211	220	212
rect	219	214	220	215
rect	219	217	220	218
rect	219	220	220	221
rect	219	223	220	224
rect	219	226	220	227
rect	219	229	220	230
rect	219	232	220	233
rect	219	235	220	236
rect	219	238	220	239
rect	219	241	220	242
rect	219	244	220	245
rect	219	247	220	248
rect	219	250	220	251
rect	219	256	220	257
rect	219	259	220	260
rect	219	265	220	266
rect	219	268	220	269
rect	219	271	220	272
rect	219	274	220	275
rect	219	277	220	278
rect	219	283	220	284
rect	219	292	220	293
rect	219	307	220	308
rect	220	7	221	8
rect	220	10	221	11
rect	220	13	221	14
rect	220	16	221	17
rect	220	19	221	20
rect	220	22	221	23
rect	220	25	221	26
rect	220	28	221	29
rect	220	31	221	32
rect	220	34	221	35
rect	220	37	221	38
rect	220	40	221	41
rect	220	43	221	44
rect	220	46	221	47
rect	220	49	221	50
rect	220	52	221	53
rect	220	55	221	56
rect	220	58	221	59
rect	220	61	221	62
rect	220	64	221	65
rect	220	67	221	68
rect	220	70	221	71
rect	220	73	221	74
rect	220	76	221	77
rect	220	79	221	80
rect	220	82	221	83
rect	220	85	221	86
rect	220	88	221	89
rect	220	91	221	92
rect	220	94	221	95
rect	220	97	221	98
rect	220	100	221	101
rect	220	103	221	104
rect	220	106	221	107
rect	220	109	221	110
rect	220	112	221	113
rect	220	115	221	116
rect	220	118	221	119
rect	220	121	221	122
rect	220	124	221	125
rect	220	127	221	128
rect	220	130	221	131
rect	220	133	221	134
rect	220	136	221	137
rect	220	139	221	140
rect	220	142	221	143
rect	220	145	221	146
rect	220	148	221	149
rect	220	151	221	152
rect	220	154	221	155
rect	220	157	221	158
rect	220	160	221	161
rect	220	163	221	164
rect	220	166	221	167
rect	220	169	221	170
rect	220	172	221	173
rect	220	175	221	176
rect	220	178	221	179
rect	220	181	221	182
rect	220	184	221	185
rect	220	187	221	188
rect	220	190	221	191
rect	220	193	221	194
rect	220	196	221	197
rect	220	199	221	200
rect	220	202	221	203
rect	220	205	221	206
rect	220	208	221	209
rect	220	211	221	212
rect	220	214	221	215
rect	220	217	221	218
rect	220	220	221	221
rect	220	223	221	224
rect	220	226	221	227
rect	220	229	221	230
rect	220	232	221	233
rect	220	235	221	236
rect	220	238	221	239
rect	220	241	221	242
rect	220	244	221	245
rect	220	247	221	248
rect	220	250	221	251
rect	220	256	221	257
rect	220	259	221	260
rect	220	265	221	266
rect	220	274	221	275
rect	220	277	221	278
rect	221	7	222	8
rect	221	10	222	11
rect	221	13	222	14
rect	221	16	222	17
rect	221	19	222	20
rect	221	22	222	23
rect	221	25	222	26
rect	221	28	222	29
rect	221	31	222	32
rect	221	34	222	35
rect	221	37	222	38
rect	221	40	222	41
rect	221	43	222	44
rect	221	46	222	47
rect	221	49	222	50
rect	221	52	222	53
rect	221	55	222	56
rect	221	58	222	59
rect	221	61	222	62
rect	221	64	222	65
rect	221	67	222	68
rect	221	70	222	71
rect	221	73	222	74
rect	221	76	222	77
rect	221	79	222	80
rect	221	82	222	83
rect	221	85	222	86
rect	221	88	222	89
rect	221	91	222	92
rect	221	94	222	95
rect	221	97	222	98
rect	221	100	222	101
rect	221	103	222	104
rect	221	106	222	107
rect	221	109	222	110
rect	221	112	222	113
rect	221	115	222	116
rect	221	118	222	119
rect	221	121	222	122
rect	221	124	222	125
rect	221	127	222	128
rect	221	130	222	131
rect	221	133	222	134
rect	221	136	222	137
rect	221	139	222	140
rect	221	142	222	143
rect	221	145	222	146
rect	221	148	222	149
rect	221	151	222	152
rect	221	154	222	155
rect	221	157	222	158
rect	221	160	222	161
rect	221	163	222	164
rect	221	166	222	167
rect	221	169	222	170
rect	221	172	222	173
rect	221	175	222	176
rect	221	178	222	179
rect	221	181	222	182
rect	221	184	222	185
rect	221	187	222	188
rect	221	190	222	191
rect	221	193	222	194
rect	221	196	222	197
rect	221	199	222	200
rect	221	202	222	203
rect	221	205	222	206
rect	221	208	222	209
rect	221	211	222	212
rect	221	214	222	215
rect	221	217	222	218
rect	221	220	222	221
rect	221	223	222	224
rect	221	226	222	227
rect	221	229	222	230
rect	221	232	222	233
rect	221	235	222	236
rect	221	238	222	239
rect	221	241	222	242
rect	221	244	222	245
rect	221	247	222	248
rect	221	250	222	251
rect	221	256	222	257
rect	221	259	222	260
rect	221	265	222	266
rect	221	274	222	275
rect	221	277	222	278
rect	222	7	223	8
rect	222	10	223	11
rect	222	13	223	14
rect	222	16	223	17
rect	222	19	223	20
rect	222	22	223	23
rect	222	25	223	26
rect	222	28	223	29
rect	222	31	223	32
rect	222	34	223	35
rect	222	37	223	38
rect	222	40	223	41
rect	222	43	223	44
rect	222	46	223	47
rect	222	49	223	50
rect	222	52	223	53
rect	222	55	223	56
rect	222	58	223	59
rect	222	61	223	62
rect	222	64	223	65
rect	222	67	223	68
rect	222	70	223	71
rect	222	73	223	74
rect	222	76	223	77
rect	222	79	223	80
rect	222	82	223	83
rect	222	85	223	86
rect	222	88	223	89
rect	222	91	223	92
rect	222	94	223	95
rect	222	97	223	98
rect	222	100	223	101
rect	222	103	223	104
rect	222	106	223	107
rect	222	109	223	110
rect	222	112	223	113
rect	222	115	223	116
rect	222	118	223	119
rect	222	121	223	122
rect	222	124	223	125
rect	222	127	223	128
rect	222	130	223	131
rect	222	133	223	134
rect	222	136	223	137
rect	222	139	223	140
rect	222	142	223	143
rect	222	145	223	146
rect	222	148	223	149
rect	222	151	223	152
rect	222	154	223	155
rect	222	157	223	158
rect	222	160	223	161
rect	222	163	223	164
rect	222	166	223	167
rect	222	169	223	170
rect	222	172	223	173
rect	222	175	223	176
rect	222	178	223	179
rect	222	181	223	182
rect	222	184	223	185
rect	222	187	223	188
rect	222	190	223	191
rect	222	193	223	194
rect	222	196	223	197
rect	222	199	223	200
rect	222	202	223	203
rect	222	205	223	206
rect	222	208	223	209
rect	222	211	223	212
rect	222	214	223	215
rect	222	217	223	218
rect	222	220	223	221
rect	222	223	223	224
rect	222	226	223	227
rect	222	229	223	230
rect	222	232	223	233
rect	222	235	223	236
rect	222	238	223	239
rect	222	241	223	242
rect	222	244	223	245
rect	222	247	223	248
rect	222	250	223	251
rect	222	256	223	257
rect	222	259	223	260
rect	222	265	223	266
rect	222	274	223	275
rect	222	277	223	278
rect	223	7	224	8
rect	223	10	224	11
rect	223	13	224	14
rect	223	16	224	17
rect	223	19	224	20
rect	223	22	224	23
rect	223	25	224	26
rect	223	28	224	29
rect	223	31	224	32
rect	223	34	224	35
rect	223	37	224	38
rect	223	40	224	41
rect	223	43	224	44
rect	223	46	224	47
rect	223	49	224	50
rect	223	52	224	53
rect	223	55	224	56
rect	223	58	224	59
rect	223	61	224	62
rect	223	64	224	65
rect	223	67	224	68
rect	223	70	224	71
rect	223	73	224	74
rect	223	76	224	77
rect	223	79	224	80
rect	223	82	224	83
rect	223	85	224	86
rect	223	88	224	89
rect	223	91	224	92
rect	223	94	224	95
rect	223	97	224	98
rect	223	100	224	101
rect	223	103	224	104
rect	223	106	224	107
rect	223	109	224	110
rect	223	112	224	113
rect	223	115	224	116
rect	223	118	224	119
rect	223	121	224	122
rect	223	124	224	125
rect	223	127	224	128
rect	223	130	224	131
rect	223	133	224	134
rect	223	136	224	137
rect	223	139	224	140
rect	223	142	224	143
rect	223	145	224	146
rect	223	148	224	149
rect	223	151	224	152
rect	223	154	224	155
rect	223	157	224	158
rect	223	160	224	161
rect	223	163	224	164
rect	223	166	224	167
rect	223	169	224	170
rect	223	172	224	173
rect	223	175	224	176
rect	223	178	224	179
rect	223	181	224	182
rect	223	184	224	185
rect	223	187	224	188
rect	223	190	224	191
rect	223	193	224	194
rect	223	196	224	197
rect	223	199	224	200
rect	223	202	224	203
rect	223	205	224	206
rect	223	208	224	209
rect	223	211	224	212
rect	223	214	224	215
rect	223	217	224	218
rect	223	220	224	221
rect	223	223	224	224
rect	223	226	224	227
rect	223	229	224	230
rect	223	232	224	233
rect	223	235	224	236
rect	223	238	224	239
rect	223	241	224	242
rect	223	244	224	245
rect	223	247	224	248
rect	223	250	224	251
rect	223	256	224	257
rect	223	259	224	260
rect	223	265	224	266
rect	223	274	224	275
rect	223	277	224	278
rect	224	7	225	8
rect	224	10	225	11
rect	224	13	225	14
rect	224	16	225	17
rect	224	19	225	20
rect	224	22	225	23
rect	224	25	225	26
rect	224	28	225	29
rect	224	31	225	32
rect	224	34	225	35
rect	224	37	225	38
rect	224	40	225	41
rect	224	43	225	44
rect	224	46	225	47
rect	224	49	225	50
rect	224	52	225	53
rect	224	55	225	56
rect	224	58	225	59
rect	224	61	225	62
rect	224	64	225	65
rect	224	67	225	68
rect	224	70	225	71
rect	224	73	225	74
rect	224	76	225	77
rect	224	79	225	80
rect	224	82	225	83
rect	224	85	225	86
rect	224	88	225	89
rect	224	91	225	92
rect	224	94	225	95
rect	224	97	225	98
rect	224	100	225	101
rect	224	103	225	104
rect	224	106	225	107
rect	224	109	225	110
rect	224	112	225	113
rect	224	115	225	116
rect	224	118	225	119
rect	224	121	225	122
rect	224	124	225	125
rect	224	127	225	128
rect	224	130	225	131
rect	224	133	225	134
rect	224	136	225	137
rect	224	139	225	140
rect	224	142	225	143
rect	224	145	225	146
rect	224	148	225	149
rect	224	151	225	152
rect	224	154	225	155
rect	224	157	225	158
rect	224	160	225	161
rect	224	163	225	164
rect	224	166	225	167
rect	224	169	225	170
rect	224	172	225	173
rect	224	175	225	176
rect	224	178	225	179
rect	224	181	225	182
rect	224	184	225	185
rect	224	187	225	188
rect	224	190	225	191
rect	224	193	225	194
rect	224	196	225	197
rect	224	199	225	200
rect	224	202	225	203
rect	224	205	225	206
rect	224	208	225	209
rect	224	211	225	212
rect	224	214	225	215
rect	224	217	225	218
rect	224	220	225	221
rect	224	223	225	224
rect	224	226	225	227
rect	224	229	225	230
rect	224	232	225	233
rect	224	235	225	236
rect	224	238	225	239
rect	224	241	225	242
rect	224	244	225	245
rect	224	247	225	248
rect	224	250	225	251
rect	224	256	225	257
rect	224	259	225	260
rect	224	265	225	266
rect	224	274	225	275
rect	224	277	225	278
rect	225	7	226	8
rect	225	10	226	11
rect	225	13	226	14
rect	225	16	226	17
rect	225	19	226	20
rect	225	22	226	23
rect	225	25	226	26
rect	225	28	226	29
rect	225	31	226	32
rect	225	34	226	35
rect	225	37	226	38
rect	225	40	226	41
rect	225	43	226	44
rect	225	46	226	47
rect	225	49	226	50
rect	225	52	226	53
rect	225	55	226	56
rect	225	58	226	59
rect	225	61	226	62
rect	225	64	226	65
rect	225	67	226	68
rect	225	70	226	71
rect	225	73	226	74
rect	225	76	226	77
rect	225	79	226	80
rect	225	82	226	83
rect	225	85	226	86
rect	225	88	226	89
rect	225	91	226	92
rect	225	94	226	95
rect	225	97	226	98
rect	225	100	226	101
rect	225	103	226	104
rect	225	106	226	107
rect	225	109	226	110
rect	225	112	226	113
rect	225	115	226	116
rect	225	118	226	119
rect	225	121	226	122
rect	225	124	226	125
rect	225	127	226	128
rect	225	130	226	131
rect	225	133	226	134
rect	225	136	226	137
rect	225	139	226	140
rect	225	142	226	143
rect	225	145	226	146
rect	225	148	226	149
rect	225	151	226	152
rect	225	154	226	155
rect	225	157	226	158
rect	225	160	226	161
rect	225	163	226	164
rect	225	166	226	167
rect	225	169	226	170
rect	225	172	226	173
rect	225	175	226	176
rect	225	178	226	179
rect	225	181	226	182
rect	225	184	226	185
rect	225	187	226	188
rect	225	190	226	191
rect	225	193	226	194
rect	225	196	226	197
rect	225	199	226	200
rect	225	202	226	203
rect	225	205	226	206
rect	225	208	226	209
rect	225	211	226	212
rect	225	214	226	215
rect	225	217	226	218
rect	225	220	226	221
rect	225	223	226	224
rect	225	226	226	227
rect	225	229	226	230
rect	225	232	226	233
rect	225	235	226	236
rect	225	238	226	239
rect	225	241	226	242
rect	225	244	226	245
rect	225	247	226	248
rect	225	250	226	251
rect	225	256	226	257
rect	225	259	226	260
rect	225	265	226	266
rect	225	274	226	275
rect	225	277	226	278
rect	226	7	227	8
rect	226	10	227	11
rect	226	13	227	14
rect	226	16	227	17
rect	226	19	227	20
rect	226	22	227	23
rect	226	25	227	26
rect	226	28	227	29
rect	226	31	227	32
rect	226	34	227	35
rect	226	37	227	38
rect	226	40	227	41
rect	226	43	227	44
rect	226	46	227	47
rect	226	49	227	50
rect	226	52	227	53
rect	226	55	227	56
rect	226	58	227	59
rect	226	61	227	62
rect	226	64	227	65
rect	226	67	227	68
rect	226	70	227	71
rect	226	73	227	74
rect	226	76	227	77
rect	226	79	227	80
rect	226	82	227	83
rect	226	85	227	86
rect	226	88	227	89
rect	226	91	227	92
rect	226	94	227	95
rect	226	97	227	98
rect	226	100	227	101
rect	226	103	227	104
rect	226	106	227	107
rect	226	109	227	110
rect	226	112	227	113
rect	226	115	227	116
rect	226	118	227	119
rect	226	121	227	122
rect	226	124	227	125
rect	226	127	227	128
rect	226	130	227	131
rect	226	133	227	134
rect	226	136	227	137
rect	226	139	227	140
rect	226	142	227	143
rect	226	145	227	146
rect	226	148	227	149
rect	226	151	227	152
rect	226	154	227	155
rect	226	157	227	158
rect	226	160	227	161
rect	226	163	227	164
rect	226	166	227	167
rect	226	169	227	170
rect	226	172	227	173
rect	226	175	227	176
rect	226	178	227	179
rect	226	181	227	182
rect	226	184	227	185
rect	226	187	227	188
rect	226	190	227	191
rect	226	193	227	194
rect	226	196	227	197
rect	226	199	227	200
rect	226	202	227	203
rect	226	205	227	206
rect	226	208	227	209
rect	226	211	227	212
rect	226	214	227	215
rect	226	217	227	218
rect	226	220	227	221
rect	226	223	227	224
rect	226	226	227	227
rect	226	229	227	230
rect	226	232	227	233
rect	226	235	227	236
rect	226	238	227	239
rect	226	241	227	242
rect	226	244	227	245
rect	226	247	227	248
rect	226	250	227	251
rect	226	256	227	257
rect	226	259	227	260
rect	226	265	227	266
rect	226	274	227	275
rect	226	277	227	278
rect	227	7	228	8
rect	227	10	228	11
rect	227	13	228	14
rect	227	16	228	17
rect	227	19	228	20
rect	227	22	228	23
rect	227	25	228	26
rect	227	28	228	29
rect	227	31	228	32
rect	227	34	228	35
rect	227	37	228	38
rect	227	40	228	41
rect	227	43	228	44
rect	227	46	228	47
rect	227	49	228	50
rect	227	52	228	53
rect	227	55	228	56
rect	227	58	228	59
rect	227	61	228	62
rect	227	64	228	65
rect	227	67	228	68
rect	227	70	228	71
rect	227	73	228	74
rect	227	76	228	77
rect	227	79	228	80
rect	227	82	228	83
rect	227	85	228	86
rect	227	88	228	89
rect	227	91	228	92
rect	227	94	228	95
rect	227	97	228	98
rect	227	100	228	101
rect	227	103	228	104
rect	227	106	228	107
rect	227	109	228	110
rect	227	112	228	113
rect	227	115	228	116
rect	227	118	228	119
rect	227	121	228	122
rect	227	124	228	125
rect	227	127	228	128
rect	227	130	228	131
rect	227	133	228	134
rect	227	136	228	137
rect	227	139	228	140
rect	227	142	228	143
rect	227	145	228	146
rect	227	148	228	149
rect	227	151	228	152
rect	227	154	228	155
rect	227	157	228	158
rect	227	160	228	161
rect	227	163	228	164
rect	227	166	228	167
rect	227	169	228	170
rect	227	172	228	173
rect	227	175	228	176
rect	227	178	228	179
rect	227	181	228	182
rect	227	184	228	185
rect	227	187	228	188
rect	227	190	228	191
rect	227	193	228	194
rect	227	196	228	197
rect	227	202	228	203
rect	227	205	228	206
rect	227	211	228	212
rect	227	214	228	215
rect	227	217	228	218
rect	227	220	228	221
rect	227	223	228	224
rect	227	226	228	227
rect	227	229	228	230
rect	227	232	228	233
rect	227	235	228	236
rect	227	238	228	239
rect	227	241	228	242
rect	227	244	228	245
rect	227	247	228	248
rect	227	250	228	251
rect	227	256	228	257
rect	227	259	228	260
rect	227	265	228	266
rect	227	274	228	275
rect	227	277	228	278
rect	228	7	229	8
rect	228	10	229	11
rect	228	13	229	14
rect	228	16	229	17
rect	228	19	229	20
rect	228	22	229	23
rect	228	25	229	26
rect	228	28	229	29
rect	228	31	229	32
rect	228	34	229	35
rect	228	37	229	38
rect	228	40	229	41
rect	228	43	229	44
rect	228	46	229	47
rect	228	49	229	50
rect	228	52	229	53
rect	228	55	229	56
rect	228	58	229	59
rect	228	61	229	62
rect	228	64	229	65
rect	228	67	229	68
rect	228	70	229	71
rect	228	73	229	74
rect	228	76	229	77
rect	228	79	229	80
rect	228	82	229	83
rect	228	85	229	86
rect	228	88	229	89
rect	228	91	229	92
rect	228	94	229	95
rect	228	97	229	98
rect	228	100	229	101
rect	228	103	229	104
rect	228	106	229	107
rect	228	109	229	110
rect	228	112	229	113
rect	228	115	229	116
rect	228	118	229	119
rect	228	121	229	122
rect	228	124	229	125
rect	228	127	229	128
rect	228	130	229	131
rect	228	133	229	134
rect	228	136	229	137
rect	228	139	229	140
rect	228	142	229	143
rect	228	145	229	146
rect	228	148	229	149
rect	228	151	229	152
rect	228	154	229	155
rect	228	157	229	158
rect	228	160	229	161
rect	228	163	229	164
rect	228	166	229	167
rect	228	169	229	170
rect	228	172	229	173
rect	228	175	229	176
rect	228	178	229	179
rect	228	181	229	182
rect	228	184	229	185
rect	228	187	229	188
rect	228	190	229	191
rect	228	193	229	194
rect	228	196	229	197
rect	228	199	229	200
rect	228	202	229	203
rect	228	205	229	206
rect	228	208	229	209
rect	228	211	229	212
rect	228	214	229	215
rect	228	217	229	218
rect	228	220	229	221
rect	228	223	229	224
rect	228	226	229	227
rect	228	229	229	230
rect	228	232	229	233
rect	228	235	229	236
rect	228	238	229	239
rect	228	241	229	242
rect	228	244	229	245
rect	228	247	229	248
rect	228	250	229	251
rect	228	256	229	257
rect	228	259	229	260
rect	228	265	229	266
rect	228	274	229	275
rect	228	277	229	278
rect	229	7	230	8
rect	229	10	230	11
rect	229	13	230	14
rect	229	16	230	17
rect	229	19	230	20
rect	229	22	230	23
rect	229	25	230	26
rect	229	28	230	29
rect	229	31	230	32
rect	229	34	230	35
rect	229	37	230	38
rect	229	40	230	41
rect	229	43	230	44
rect	229	46	230	47
rect	229	49	230	50
rect	229	52	230	53
rect	229	55	230	56
rect	229	58	230	59
rect	229	61	230	62
rect	229	64	230	65
rect	229	67	230	68
rect	229	70	230	71
rect	229	73	230	74
rect	229	76	230	77
rect	229	79	230	80
rect	229	82	230	83
rect	229	85	230	86
rect	229	88	230	89
rect	229	91	230	92
rect	229	94	230	95
rect	229	97	230	98
rect	229	100	230	101
rect	229	103	230	104
rect	229	106	230	107
rect	229	109	230	110
rect	229	112	230	113
rect	229	115	230	116
rect	229	118	230	119
rect	229	121	230	122
rect	229	124	230	125
rect	229	127	230	128
rect	229	130	230	131
rect	229	133	230	134
rect	229	136	230	137
rect	229	139	230	140
rect	229	142	230	143
rect	229	145	230	146
rect	229	148	230	149
rect	229	151	230	152
rect	229	154	230	155
rect	229	157	230	158
rect	229	160	230	161
rect	229	163	230	164
rect	229	166	230	167
rect	229	169	230	170
rect	229	172	230	173
rect	229	175	230	176
rect	229	178	230	179
rect	229	181	230	182
rect	229	184	230	185
rect	229	187	230	188
rect	229	190	230	191
rect	229	193	230	194
rect	229	196	230	197
rect	229	199	230	200
rect	229	205	230	206
rect	229	211	230	212
rect	229	214	230	215
rect	229	217	230	218
rect	229	220	230	221
rect	229	223	230	224
rect	229	226	230	227
rect	229	229	230	230
rect	229	232	230	233
rect	229	235	230	236
rect	229	238	230	239
rect	229	241	230	242
rect	229	244	230	245
rect	229	247	230	248
rect	229	250	230	251
rect	229	256	230	257
rect	229	259	230	260
rect	229	265	230	266
rect	229	274	230	275
rect	229	277	230	278
rect	230	7	231	8
rect	230	10	231	11
rect	230	13	231	14
rect	230	16	231	17
rect	230	19	231	20
rect	230	22	231	23
rect	230	25	231	26
rect	230	28	231	29
rect	230	31	231	32
rect	230	34	231	35
rect	230	37	231	38
rect	230	40	231	41
rect	230	43	231	44
rect	230	46	231	47
rect	230	49	231	50
rect	230	52	231	53
rect	230	55	231	56
rect	230	58	231	59
rect	230	61	231	62
rect	230	64	231	65
rect	230	67	231	68
rect	230	70	231	71
rect	230	73	231	74
rect	230	76	231	77
rect	230	79	231	80
rect	230	82	231	83
rect	230	85	231	86
rect	230	88	231	89
rect	230	91	231	92
rect	230	94	231	95
rect	230	97	231	98
rect	230	100	231	101
rect	230	103	231	104
rect	230	106	231	107
rect	230	109	231	110
rect	230	112	231	113
rect	230	115	231	116
rect	230	118	231	119
rect	230	121	231	122
rect	230	124	231	125
rect	230	127	231	128
rect	230	133	231	134
rect	230	136	231	137
rect	230	139	231	140
rect	230	142	231	143
rect	230	145	231	146
rect	230	148	231	149
rect	230	151	231	152
rect	230	154	231	155
rect	230	157	231	158
rect	230	160	231	161
rect	230	163	231	164
rect	230	166	231	167
rect	230	169	231	170
rect	230	172	231	173
rect	230	175	231	176
rect	230	178	231	179
rect	230	181	231	182
rect	230	184	231	185
rect	230	187	231	188
rect	230	190	231	191
rect	230	193	231	194
rect	230	196	231	197
rect	230	199	231	200
rect	230	202	231	203
rect	230	205	231	206
rect	230	208	231	209
rect	230	211	231	212
rect	230	214	231	215
rect	230	217	231	218
rect	230	220	231	221
rect	230	223	231	224
rect	230	226	231	227
rect	230	229	231	230
rect	230	232	231	233
rect	230	235	231	236
rect	230	238	231	239
rect	230	241	231	242
rect	230	244	231	245
rect	230	247	231	248
rect	230	250	231	251
rect	230	256	231	257
rect	230	259	231	260
rect	230	265	231	266
rect	230	274	231	275
rect	231	7	232	8
rect	231	10	232	11
rect	231	13	232	14
rect	231	16	232	17
rect	231	19	232	20
rect	231	22	232	23
rect	231	25	232	26
rect	231	28	232	29
rect	231	31	232	32
rect	231	34	232	35
rect	231	37	232	38
rect	231	40	232	41
rect	231	43	232	44
rect	231	46	232	47
rect	231	49	232	50
rect	231	52	232	53
rect	231	55	232	56
rect	231	58	232	59
rect	231	61	232	62
rect	231	64	232	65
rect	231	67	232	68
rect	231	70	232	71
rect	231	73	232	74
rect	231	76	232	77
rect	231	79	232	80
rect	231	82	232	83
rect	231	85	232	86
rect	231	88	232	89
rect	231	91	232	92
rect	231	94	232	95
rect	231	97	232	98
rect	231	100	232	101
rect	231	103	232	104
rect	231	106	232	107
rect	231	109	232	110
rect	231	112	232	113
rect	231	115	232	116
rect	231	118	232	119
rect	231	121	232	122
rect	231	124	232	125
rect	231	127	232	128
rect	231	133	232	134
rect	231	136	232	137
rect	231	142	232	143
rect	231	145	232	146
rect	231	148	232	149
rect	231	151	232	152
rect	231	154	232	155
rect	231	157	232	158
rect	231	160	232	161
rect	231	163	232	164
rect	231	166	232	167
rect	231	169	232	170
rect	231	172	232	173
rect	231	175	232	176
rect	231	178	232	179
rect	231	181	232	182
rect	231	184	232	185
rect	231	187	232	188
rect	231	190	232	191
rect	231	193	232	194
rect	231	196	232	197
rect	231	199	232	200
rect	231	202	232	203
rect	231	205	232	206
rect	231	208	232	209
rect	231	211	232	212
rect	231	214	232	215
rect	231	217	232	218
rect	231	220	232	221
rect	231	223	232	224
rect	231	226	232	227
rect	231	229	232	230
rect	231	232	232	233
rect	231	235	232	236
rect	231	238	232	239
rect	231	241	232	242
rect	231	244	232	245
rect	231	247	232	248
rect	231	250	232	251
rect	231	256	232	257
rect	231	259	232	260
rect	231	265	232	266
rect	231	274	232	275
rect	232	7	233	8
rect	232	10	233	11
rect	232	13	233	14
rect	232	16	233	17
rect	232	19	233	20
rect	232	22	233	23
rect	232	25	233	26
rect	232	28	233	29
rect	232	31	233	32
rect	232	34	233	35
rect	232	37	233	38
rect	232	40	233	41
rect	232	43	233	44
rect	232	46	233	47
rect	232	49	233	50
rect	232	52	233	53
rect	232	55	233	56
rect	232	58	233	59
rect	232	61	233	62
rect	232	64	233	65
rect	232	67	233	68
rect	232	70	233	71
rect	232	73	233	74
rect	232	76	233	77
rect	232	79	233	80
rect	232	82	233	83
rect	232	85	233	86
rect	232	88	233	89
rect	232	91	233	92
rect	232	94	233	95
rect	232	97	233	98
rect	232	100	233	101
rect	232	103	233	104
rect	232	106	233	107
rect	232	109	233	110
rect	232	112	233	113
rect	232	115	233	116
rect	232	118	233	119
rect	232	121	233	122
rect	232	124	233	125
rect	232	127	233	128
rect	232	133	233	134
rect	232	136	233	137
rect	232	139	233	140
rect	232	142	233	143
rect	232	145	233	146
rect	232	148	233	149
rect	232	151	233	152
rect	232	154	233	155
rect	232	157	233	158
rect	232	160	233	161
rect	232	163	233	164
rect	232	166	233	167
rect	232	169	233	170
rect	232	172	233	173
rect	232	175	233	176
rect	232	178	233	179
rect	232	181	233	182
rect	232	184	233	185
rect	232	187	233	188
rect	232	190	233	191
rect	232	193	233	194
rect	232	196	233	197
rect	232	199	233	200
rect	232	202	233	203
rect	232	205	233	206
rect	232	208	233	209
rect	232	211	233	212
rect	232	214	233	215
rect	232	217	233	218
rect	232	220	233	221
rect	232	223	233	224
rect	232	226	233	227
rect	232	229	233	230
rect	232	232	233	233
rect	232	235	233	236
rect	232	238	233	239
rect	232	241	233	242
rect	232	244	233	245
rect	232	247	233	248
rect	232	250	233	251
rect	232	256	233	257
rect	232	259	233	260
rect	232	265	233	266
rect	232	274	233	275
rect	233	7	234	8
rect	233	10	234	11
rect	233	13	234	14
rect	233	16	234	17
rect	233	19	234	20
rect	233	22	234	23
rect	233	25	234	26
rect	233	28	234	29
rect	233	31	234	32
rect	233	34	234	35
rect	233	37	234	38
rect	233	40	234	41
rect	233	43	234	44
rect	233	46	234	47
rect	233	49	234	50
rect	233	52	234	53
rect	233	55	234	56
rect	233	58	234	59
rect	233	61	234	62
rect	233	64	234	65
rect	233	67	234	68
rect	233	73	234	74
rect	233	76	234	77
rect	233	79	234	80
rect	233	82	234	83
rect	233	85	234	86
rect	233	88	234	89
rect	233	91	234	92
rect	233	94	234	95
rect	233	97	234	98
rect	233	100	234	101
rect	233	103	234	104
rect	233	106	234	107
rect	233	109	234	110
rect	233	112	234	113
rect	233	115	234	116
rect	233	118	234	119
rect	233	121	234	122
rect	233	124	234	125
rect	233	127	234	128
rect	233	133	234	134
rect	233	136	234	137
rect	233	139	234	140
rect	233	142	234	143
rect	233	145	234	146
rect	233	148	234	149
rect	233	151	234	152
rect	233	154	234	155
rect	233	157	234	158
rect	233	160	234	161
rect	233	163	234	164
rect	233	166	234	167
rect	233	169	234	170
rect	233	172	234	173
rect	233	175	234	176
rect	233	178	234	179
rect	233	181	234	182
rect	233	184	234	185
rect	233	187	234	188
rect	233	190	234	191
rect	233	193	234	194
rect	233	196	234	197
rect	233	199	234	200
rect	233	202	234	203
rect	233	205	234	206
rect	233	208	234	209
rect	233	211	234	212
rect	233	214	234	215
rect	233	217	234	218
rect	233	220	234	221
rect	233	223	234	224
rect	233	226	234	227
rect	233	229	234	230
rect	233	232	234	233
rect	233	235	234	236
rect	233	238	234	239
rect	233	244	234	245
rect	233	247	234	248
rect	233	250	234	251
rect	233	256	234	257
rect	233	259	234	260
rect	233	265	234	266
rect	233	274	234	275
rect	234	7	235	8
rect	234	10	235	11
rect	234	13	235	14
rect	234	16	235	17
rect	234	19	235	20
rect	234	22	235	23
rect	234	25	235	26
rect	234	28	235	29
rect	234	31	235	32
rect	234	34	235	35
rect	234	37	235	38
rect	234	40	235	41
rect	234	43	235	44
rect	234	46	235	47
rect	234	49	235	50
rect	234	52	235	53
rect	234	55	235	56
rect	234	58	235	59
rect	234	61	235	62
rect	234	64	235	65
rect	234	67	235	68
rect	234	70	235	71
rect	234	73	235	74
rect	234	76	235	77
rect	234	79	235	80
rect	234	82	235	83
rect	234	85	235	86
rect	234	88	235	89
rect	234	91	235	92
rect	234	94	235	95
rect	234	97	235	98
rect	234	100	235	101
rect	234	103	235	104
rect	234	106	235	107
rect	234	109	235	110
rect	234	112	235	113
rect	234	115	235	116
rect	234	118	235	119
rect	234	121	235	122
rect	234	124	235	125
rect	234	127	235	128
rect	234	133	235	134
rect	234	136	235	137
rect	234	139	235	140
rect	234	142	235	143
rect	234	145	235	146
rect	234	148	235	149
rect	234	151	235	152
rect	234	154	235	155
rect	234	157	235	158
rect	234	160	235	161
rect	234	163	235	164
rect	234	166	235	167
rect	234	169	235	170
rect	234	172	235	173
rect	234	175	235	176
rect	234	178	235	179
rect	234	181	235	182
rect	234	184	235	185
rect	234	187	235	188
rect	234	190	235	191
rect	234	193	235	194
rect	234	196	235	197
rect	234	199	235	200
rect	234	202	235	203
rect	234	205	235	206
rect	234	208	235	209
rect	234	211	235	212
rect	234	214	235	215
rect	234	217	235	218
rect	234	220	235	221
rect	234	223	235	224
rect	234	226	235	227
rect	234	229	235	230
rect	234	232	235	233
rect	234	235	235	236
rect	234	238	235	239
rect	234	241	235	242
rect	234	244	235	245
rect	234	247	235	248
rect	234	250	235	251
rect	234	256	235	257
rect	234	259	235	260
rect	234	265	235	266
rect	234	274	235	275
rect	235	7	236	8
rect	235	10	236	11
rect	235	13	236	14
rect	235	16	236	17
rect	235	19	236	20
rect	235	22	236	23
rect	235	25	236	26
rect	235	28	236	29
rect	235	31	236	32
rect	235	34	236	35
rect	235	37	236	38
rect	235	40	236	41
rect	235	43	236	44
rect	235	46	236	47
rect	235	49	236	50
rect	235	52	236	53
rect	235	55	236	56
rect	235	58	236	59
rect	235	61	236	62
rect	235	64	236	65
rect	235	67	236	68
rect	235	70	236	71
rect	235	73	236	74
rect	235	76	236	77
rect	235	79	236	80
rect	235	82	236	83
rect	235	85	236	86
rect	235	88	236	89
rect	235	94	236	95
rect	235	97	236	98
rect	235	100	236	101
rect	235	103	236	104
rect	235	106	236	107
rect	235	109	236	110
rect	235	112	236	113
rect	235	115	236	116
rect	235	118	236	119
rect	235	121	236	122
rect	235	124	236	125
rect	235	127	236	128
rect	235	133	236	134
rect	235	136	236	137
rect	235	139	236	140
rect	235	142	236	143
rect	235	145	236	146
rect	235	148	236	149
rect	235	151	236	152
rect	235	154	236	155
rect	235	157	236	158
rect	235	160	236	161
rect	235	163	236	164
rect	235	166	236	167
rect	235	169	236	170
rect	235	172	236	173
rect	235	175	236	176
rect	235	178	236	179
rect	235	181	236	182
rect	235	184	236	185
rect	235	187	236	188
rect	235	193	236	194
rect	235	196	236	197
rect	235	199	236	200
rect	235	202	236	203
rect	235	205	236	206
rect	235	208	236	209
rect	235	211	236	212
rect	235	214	236	215
rect	235	217	236	218
rect	235	220	236	221
rect	235	223	236	224
rect	235	226	236	227
rect	235	229	236	230
rect	235	232	236	233
rect	235	235	236	236
rect	235	238	236	239
rect	235	241	236	242
rect	235	244	236	245
rect	235	247	236	248
rect	235	250	236	251
rect	235	256	236	257
rect	235	259	236	260
rect	236	7	237	8
rect	236	10	237	11
rect	236	13	237	14
rect	236	16	237	17
rect	236	19	237	20
rect	236	22	237	23
rect	236	25	237	26
rect	236	28	237	29
rect	236	31	237	32
rect	236	34	237	35
rect	236	37	237	38
rect	236	40	237	41
rect	236	43	237	44
rect	236	46	237	47
rect	236	49	237	50
rect	236	52	237	53
rect	236	55	237	56
rect	236	58	237	59
rect	236	61	237	62
rect	236	64	237	65
rect	236	67	237	68
rect	236	70	237	71
rect	236	73	237	74
rect	236	76	237	77
rect	236	79	237	80
rect	236	82	237	83
rect	236	85	237	86
rect	236	88	237	89
rect	236	94	237	95
rect	236	97	237	98
rect	236	100	237	101
rect	236	103	237	104
rect	236	106	237	107
rect	236	109	237	110
rect	236	112	237	113
rect	236	115	237	116
rect	236	118	237	119
rect	236	121	237	122
rect	236	124	237	125
rect	236	127	237	128
rect	236	133	237	134
rect	236	136	237	137
rect	236	139	237	140
rect	236	142	237	143
rect	236	145	237	146
rect	236	148	237	149
rect	236	151	237	152
rect	236	154	237	155
rect	236	157	237	158
rect	236	160	237	161
rect	236	163	237	164
rect	236	166	237	167
rect	236	169	237	170
rect	236	172	237	173
rect	236	175	237	176
rect	236	178	237	179
rect	236	181	237	182
rect	236	184	237	185
rect	236	187	237	188
rect	236	193	237	194
rect	236	196	237	197
rect	236	199	237	200
rect	236	202	237	203
rect	236	205	237	206
rect	236	208	237	209
rect	236	211	237	212
rect	236	214	237	215
rect	236	217	237	218
rect	236	220	237	221
rect	236	223	237	224
rect	236	226	237	227
rect	236	229	237	230
rect	236	232	237	233
rect	236	235	237	236
rect	236	238	237	239
rect	236	241	237	242
rect	236	244	237	245
rect	236	247	237	248
rect	236	250	237	251
rect	236	256	237	257
rect	236	259	237	260
rect	237	7	238	8
rect	237	10	238	11
rect	237	13	238	14
rect	237	16	238	17
rect	237	19	238	20
rect	237	22	238	23
rect	237	25	238	26
rect	237	28	238	29
rect	237	31	238	32
rect	237	34	238	35
rect	237	37	238	38
rect	237	40	238	41
rect	237	43	238	44
rect	237	46	238	47
rect	237	49	238	50
rect	237	52	238	53
rect	237	55	238	56
rect	237	58	238	59
rect	237	61	238	62
rect	237	64	238	65
rect	237	67	238	68
rect	237	70	238	71
rect	237	73	238	74
rect	237	76	238	77
rect	237	79	238	80
rect	237	82	238	83
rect	237	85	238	86
rect	237	88	238	89
rect	237	94	238	95
rect	237	97	238	98
rect	237	100	238	101
rect	237	103	238	104
rect	237	106	238	107
rect	237	109	238	110
rect	237	112	238	113
rect	237	115	238	116
rect	237	118	238	119
rect	237	121	238	122
rect	237	124	238	125
rect	237	127	238	128
rect	237	133	238	134
rect	237	136	238	137
rect	237	139	238	140
rect	237	142	238	143
rect	237	145	238	146
rect	237	148	238	149
rect	237	151	238	152
rect	237	154	238	155
rect	237	157	238	158
rect	237	160	238	161
rect	237	163	238	164
rect	237	166	238	167
rect	237	169	238	170
rect	237	172	238	173
rect	237	175	238	176
rect	237	178	238	179
rect	237	181	238	182
rect	237	184	238	185
rect	237	187	238	188
rect	237	193	238	194
rect	237	196	238	197
rect	237	199	238	200
rect	237	202	238	203
rect	237	205	238	206
rect	237	208	238	209
rect	237	211	238	212
rect	237	214	238	215
rect	237	217	238	218
rect	237	220	238	221
rect	237	223	238	224
rect	237	226	238	227
rect	237	229	238	230
rect	237	232	238	233
rect	237	235	238	236
rect	237	238	238	239
rect	237	241	238	242
rect	237	244	238	245
rect	237	247	238	248
rect	237	250	238	251
rect	237	256	238	257
rect	237	259	238	260
rect	238	7	239	8
rect	238	10	239	11
rect	238	13	239	14
rect	238	16	239	17
rect	238	19	239	20
rect	238	22	239	23
rect	238	25	239	26
rect	238	28	239	29
rect	238	31	239	32
rect	238	34	239	35
rect	238	37	239	38
rect	238	40	239	41
rect	238	43	239	44
rect	238	46	239	47
rect	238	49	239	50
rect	238	52	239	53
rect	238	55	239	56
rect	238	58	239	59
rect	238	61	239	62
rect	238	64	239	65
rect	238	67	239	68
rect	238	70	239	71
rect	238	73	239	74
rect	238	76	239	77
rect	238	79	239	80
rect	238	82	239	83
rect	238	85	239	86
rect	238	88	239	89
rect	238	94	239	95
rect	238	97	239	98
rect	238	100	239	101
rect	238	103	239	104
rect	238	106	239	107
rect	238	109	239	110
rect	238	112	239	113
rect	238	115	239	116
rect	238	118	239	119
rect	238	121	239	122
rect	238	124	239	125
rect	238	127	239	128
rect	238	133	239	134
rect	238	136	239	137
rect	238	139	239	140
rect	238	142	239	143
rect	238	145	239	146
rect	238	148	239	149
rect	238	151	239	152
rect	238	154	239	155
rect	238	157	239	158
rect	238	160	239	161
rect	238	163	239	164
rect	238	166	239	167
rect	238	169	239	170
rect	238	172	239	173
rect	238	175	239	176
rect	238	178	239	179
rect	238	181	239	182
rect	238	184	239	185
rect	238	187	239	188
rect	238	193	239	194
rect	238	196	239	197
rect	238	199	239	200
rect	238	202	239	203
rect	238	205	239	206
rect	238	208	239	209
rect	238	211	239	212
rect	238	214	239	215
rect	238	217	239	218
rect	238	220	239	221
rect	238	223	239	224
rect	238	226	239	227
rect	238	229	239	230
rect	238	232	239	233
rect	238	235	239	236
rect	238	238	239	239
rect	238	241	239	242
rect	238	244	239	245
rect	238	247	239	248
rect	238	250	239	251
rect	238	256	239	257
rect	238	259	239	260
rect	239	7	240	8
rect	239	10	240	11
rect	239	13	240	14
rect	239	16	240	17
rect	239	19	240	20
rect	239	22	240	23
rect	239	25	240	26
rect	239	28	240	29
rect	239	31	240	32
rect	239	34	240	35
rect	239	37	240	38
rect	239	40	240	41
rect	239	43	240	44
rect	239	46	240	47
rect	239	49	240	50
rect	239	52	240	53
rect	239	55	240	56
rect	239	58	240	59
rect	239	61	240	62
rect	239	64	240	65
rect	239	67	240	68
rect	239	70	240	71
rect	239	73	240	74
rect	239	76	240	77
rect	239	79	240	80
rect	239	82	240	83
rect	239	85	240	86
rect	239	88	240	89
rect	239	94	240	95
rect	239	97	240	98
rect	239	100	240	101
rect	239	103	240	104
rect	239	106	240	107
rect	239	109	240	110
rect	239	112	240	113
rect	239	115	240	116
rect	239	118	240	119
rect	239	121	240	122
rect	239	124	240	125
rect	239	127	240	128
rect	239	133	240	134
rect	239	136	240	137
rect	239	139	240	140
rect	239	142	240	143
rect	239	145	240	146
rect	239	148	240	149
rect	239	151	240	152
rect	239	154	240	155
rect	239	157	240	158
rect	239	160	240	161
rect	239	163	240	164
rect	239	166	240	167
rect	239	169	240	170
rect	239	172	240	173
rect	239	175	240	176
rect	239	178	240	179
rect	239	181	240	182
rect	239	184	240	185
rect	239	187	240	188
rect	239	193	240	194
rect	239	196	240	197
rect	239	199	240	200
rect	239	202	240	203
rect	239	205	240	206
rect	239	208	240	209
rect	239	211	240	212
rect	239	214	240	215
rect	239	217	240	218
rect	239	220	240	221
rect	239	223	240	224
rect	239	226	240	227
rect	239	229	240	230
rect	239	232	240	233
rect	239	235	240	236
rect	239	238	240	239
rect	239	241	240	242
rect	239	244	240	245
rect	239	247	240	248
rect	239	250	240	251
rect	239	256	240	257
rect	239	259	240	260
rect	240	7	241	8
rect	240	10	241	11
rect	240	13	241	14
rect	240	16	241	17
rect	240	19	241	20
rect	240	22	241	23
rect	240	25	241	26
rect	240	28	241	29
rect	240	31	241	32
rect	240	34	241	35
rect	240	37	241	38
rect	240	40	241	41
rect	240	43	241	44
rect	240	46	241	47
rect	240	49	241	50
rect	240	52	241	53
rect	240	55	241	56
rect	240	58	241	59
rect	240	61	241	62
rect	240	64	241	65
rect	240	67	241	68
rect	240	70	241	71
rect	240	73	241	74
rect	240	76	241	77
rect	240	79	241	80
rect	240	82	241	83
rect	240	85	241	86
rect	240	88	241	89
rect	240	94	241	95
rect	240	97	241	98
rect	240	100	241	101
rect	240	103	241	104
rect	240	106	241	107
rect	240	109	241	110
rect	240	112	241	113
rect	240	115	241	116
rect	240	118	241	119
rect	240	121	241	122
rect	240	124	241	125
rect	240	127	241	128
rect	240	133	241	134
rect	240	136	241	137
rect	240	139	241	140
rect	240	142	241	143
rect	240	145	241	146
rect	240	148	241	149
rect	240	151	241	152
rect	240	154	241	155
rect	240	157	241	158
rect	240	160	241	161
rect	240	163	241	164
rect	240	166	241	167
rect	240	169	241	170
rect	240	172	241	173
rect	240	175	241	176
rect	240	178	241	179
rect	240	181	241	182
rect	240	184	241	185
rect	240	187	241	188
rect	240	193	241	194
rect	240	196	241	197
rect	240	199	241	200
rect	240	202	241	203
rect	240	205	241	206
rect	240	208	241	209
rect	240	211	241	212
rect	240	214	241	215
rect	240	217	241	218
rect	240	220	241	221
rect	240	223	241	224
rect	240	226	241	227
rect	240	229	241	230
rect	240	232	241	233
rect	240	235	241	236
rect	240	238	241	239
rect	240	241	241	242
rect	240	244	241	245
rect	240	247	241	248
rect	240	250	241	251
rect	240	256	241	257
rect	240	259	241	260
rect	241	7	242	8
rect	241	10	242	11
rect	241	13	242	14
rect	241	16	242	17
rect	241	19	242	20
rect	241	22	242	23
rect	241	25	242	26
rect	241	28	242	29
rect	241	31	242	32
rect	241	34	242	35
rect	241	37	242	38
rect	241	40	242	41
rect	241	43	242	44
rect	241	46	242	47
rect	241	49	242	50
rect	241	52	242	53
rect	241	55	242	56
rect	241	58	242	59
rect	241	61	242	62
rect	241	64	242	65
rect	241	67	242	68
rect	241	70	242	71
rect	241	73	242	74
rect	241	76	242	77
rect	241	79	242	80
rect	241	82	242	83
rect	241	85	242	86
rect	241	88	242	89
rect	241	94	242	95
rect	241	97	242	98
rect	241	100	242	101
rect	241	103	242	104
rect	241	106	242	107
rect	241	109	242	110
rect	241	112	242	113
rect	241	115	242	116
rect	241	118	242	119
rect	241	124	242	125
rect	241	127	242	128
rect	241	133	242	134
rect	241	136	242	137
rect	241	139	242	140
rect	241	142	242	143
rect	241	145	242	146
rect	241	148	242	149
rect	241	151	242	152
rect	241	154	242	155
rect	241	157	242	158
rect	241	160	242	161
rect	241	163	242	164
rect	241	166	242	167
rect	241	169	242	170
rect	241	172	242	173
rect	241	175	242	176
rect	241	178	242	179
rect	241	181	242	182
rect	241	184	242	185
rect	241	187	242	188
rect	241	193	242	194
rect	241	196	242	197
rect	241	199	242	200
rect	241	202	242	203
rect	241	205	242	206
rect	241	208	242	209
rect	241	211	242	212
rect	241	214	242	215
rect	241	217	242	218
rect	241	220	242	221
rect	241	223	242	224
rect	241	226	242	227
rect	241	229	242	230
rect	241	232	242	233
rect	241	235	242	236
rect	241	238	242	239
rect	241	244	242	245
rect	241	247	242	248
rect	241	250	242	251
rect	241	256	242	257
rect	241	259	242	260
rect	242	7	243	8
rect	242	10	243	11
rect	242	13	243	14
rect	242	16	243	17
rect	242	19	243	20
rect	242	22	243	23
rect	242	25	243	26
rect	242	28	243	29
rect	242	31	243	32
rect	242	34	243	35
rect	242	37	243	38
rect	242	40	243	41
rect	242	43	243	44
rect	242	46	243	47
rect	242	49	243	50
rect	242	52	243	53
rect	242	55	243	56
rect	242	58	243	59
rect	242	61	243	62
rect	242	64	243	65
rect	242	67	243	68
rect	242	70	243	71
rect	242	73	243	74
rect	242	76	243	77
rect	242	79	243	80
rect	242	82	243	83
rect	242	85	243	86
rect	242	88	243	89
rect	242	94	243	95
rect	242	97	243	98
rect	242	100	243	101
rect	242	103	243	104
rect	242	106	243	107
rect	242	109	243	110
rect	242	112	243	113
rect	242	115	243	116
rect	242	118	243	119
rect	242	124	243	125
rect	242	127	243	128
rect	242	133	243	134
rect	242	136	243	137
rect	242	139	243	140
rect	242	142	243	143
rect	242	145	243	146
rect	242	148	243	149
rect	242	151	243	152
rect	242	154	243	155
rect	242	157	243	158
rect	242	160	243	161
rect	242	163	243	164
rect	242	166	243	167
rect	242	169	243	170
rect	242	172	243	173
rect	242	175	243	176
rect	242	178	243	179
rect	242	181	243	182
rect	242	184	243	185
rect	242	187	243	188
rect	242	193	243	194
rect	242	196	243	197
rect	242	199	243	200
rect	242	202	243	203
rect	242	205	243	206
rect	242	208	243	209
rect	242	211	243	212
rect	242	214	243	215
rect	242	217	243	218
rect	242	220	243	221
rect	242	223	243	224
rect	242	226	243	227
rect	242	229	243	230
rect	242	232	243	233
rect	242	235	243	236
rect	242	238	243	239
rect	242	247	243	248
rect	242	250	243	251
rect	242	256	243	257
rect	242	259	243	260
rect	243	7	244	8
rect	243	10	244	11
rect	243	13	244	14
rect	243	16	244	17
rect	243	19	244	20
rect	243	22	244	23
rect	243	25	244	26
rect	243	28	244	29
rect	243	31	244	32
rect	243	34	244	35
rect	243	37	244	38
rect	243	40	244	41
rect	243	43	244	44
rect	243	46	244	47
rect	243	49	244	50
rect	243	52	244	53
rect	243	55	244	56
rect	243	58	244	59
rect	243	61	244	62
rect	243	64	244	65
rect	243	67	244	68
rect	243	70	244	71
rect	243	73	244	74
rect	243	76	244	77
rect	243	79	244	80
rect	243	82	244	83
rect	243	85	244	86
rect	243	88	244	89
rect	243	94	244	95
rect	243	97	244	98
rect	243	100	244	101
rect	243	103	244	104
rect	243	106	244	107
rect	243	109	244	110
rect	243	112	244	113
rect	243	115	244	116
rect	243	118	244	119
rect	243	124	244	125
rect	243	127	244	128
rect	243	133	244	134
rect	243	136	244	137
rect	243	139	244	140
rect	243	142	244	143
rect	243	145	244	146
rect	243	148	244	149
rect	243	151	244	152
rect	243	154	244	155
rect	243	157	244	158
rect	243	160	244	161
rect	243	163	244	164
rect	243	166	244	167
rect	243	169	244	170
rect	243	172	244	173
rect	243	175	244	176
rect	243	178	244	179
rect	243	181	244	182
rect	243	184	244	185
rect	243	187	244	188
rect	243	193	244	194
rect	243	196	244	197
rect	243	199	244	200
rect	243	202	244	203
rect	243	205	244	206
rect	243	208	244	209
rect	243	211	244	212
rect	243	214	244	215
rect	243	217	244	218
rect	243	220	244	221
rect	243	223	244	224
rect	243	226	244	227
rect	243	229	244	230
rect	243	232	244	233
rect	243	235	244	236
rect	243	238	244	239
rect	243	244	244	245
rect	243	247	244	248
rect	243	250	244	251
rect	243	256	244	257
rect	243	259	244	260
rect	244	7	245	8
rect	244	10	245	11
rect	244	13	245	14
rect	244	16	245	17
rect	244	19	245	20
rect	244	22	245	23
rect	244	25	245	26
rect	244	28	245	29
rect	244	31	245	32
rect	244	34	245	35
rect	244	37	245	38
rect	244	40	245	41
rect	244	43	245	44
rect	244	46	245	47
rect	244	49	245	50
rect	244	52	245	53
rect	244	55	245	56
rect	244	58	245	59
rect	244	61	245	62
rect	244	64	245	65
rect	244	67	245	68
rect	244	70	245	71
rect	244	73	245	74
rect	244	76	245	77
rect	244	79	245	80
rect	244	82	245	83
rect	244	85	245	86
rect	244	88	245	89
rect	244	94	245	95
rect	244	97	245	98
rect	244	100	245	101
rect	244	103	245	104
rect	244	106	245	107
rect	244	109	245	110
rect	244	112	245	113
rect	244	115	245	116
rect	244	118	245	119
rect	244	124	245	125
rect	244	127	245	128
rect	244	133	245	134
rect	244	136	245	137
rect	244	139	245	140
rect	244	142	245	143
rect	244	145	245	146
rect	244	148	245	149
rect	244	151	245	152
rect	244	154	245	155
rect	244	157	245	158
rect	244	160	245	161
rect	244	163	245	164
rect	244	166	245	167
rect	244	169	245	170
rect	244	172	245	173
rect	244	175	245	176
rect	244	178	245	179
rect	244	181	245	182
rect	244	184	245	185
rect	244	187	245	188
rect	244	193	245	194
rect	244	199	245	200
rect	244	202	245	203
rect	244	205	245	206
rect	244	208	245	209
rect	244	214	245	215
rect	244	217	245	218
rect	244	220	245	221
rect	244	223	245	224
rect	244	226	245	227
rect	244	229	245	230
rect	244	232	245	233
rect	244	235	245	236
rect	244	238	245	239
rect	244	244	245	245
rect	244	247	245	248
rect	244	250	245	251
rect	244	256	245	257
rect	244	259	245	260
rect	245	7	246	8
rect	245	10	246	11
rect	245	13	246	14
rect	245	16	246	17
rect	245	19	246	20
rect	245	22	246	23
rect	245	25	246	26
rect	245	28	246	29
rect	245	31	246	32
rect	245	34	246	35
rect	245	37	246	38
rect	245	40	246	41
rect	245	43	246	44
rect	245	46	246	47
rect	245	49	246	50
rect	245	52	246	53
rect	245	55	246	56
rect	245	58	246	59
rect	245	61	246	62
rect	245	64	246	65
rect	245	67	246	68
rect	245	70	246	71
rect	245	73	246	74
rect	245	76	246	77
rect	245	79	246	80
rect	245	82	246	83
rect	245	85	246	86
rect	245	88	246	89
rect	245	94	246	95
rect	245	97	246	98
rect	245	100	246	101
rect	245	103	246	104
rect	245	106	246	107
rect	245	109	246	110
rect	245	112	246	113
rect	245	115	246	116
rect	245	118	246	119
rect	245	121	246	122
rect	245	124	246	125
rect	245	127	246	128
rect	245	133	246	134
rect	245	136	246	137
rect	245	139	246	140
rect	245	142	246	143
rect	245	145	246	146
rect	245	148	246	149
rect	245	151	246	152
rect	245	154	246	155
rect	245	157	246	158
rect	245	160	246	161
rect	245	163	246	164
rect	245	166	246	167
rect	245	169	246	170
rect	245	172	246	173
rect	245	175	246	176
rect	245	178	246	179
rect	245	181	246	182
rect	245	184	246	185
rect	245	187	246	188
rect	245	193	246	194
rect	245	196	246	197
rect	245	199	246	200
rect	245	202	246	203
rect	245	205	246	206
rect	245	208	246	209
rect	245	211	246	212
rect	245	214	246	215
rect	245	217	246	218
rect	245	220	246	221
rect	245	223	246	224
rect	245	226	246	227
rect	245	229	246	230
rect	245	232	246	233
rect	245	235	246	236
rect	245	238	246	239
rect	245	241	246	242
rect	245	244	246	245
rect	245	247	246	248
rect	245	250	246	251
rect	245	256	246	257
rect	245	259	246	260
rect	246	7	247	8
rect	246	10	247	11
rect	246	13	247	14
rect	246	16	247	17
rect	246	19	247	20
rect	246	22	247	23
rect	246	25	247	26
rect	246	28	247	29
rect	246	31	247	32
rect	246	34	247	35
rect	246	37	247	38
rect	246	40	247	41
rect	246	43	247	44
rect	246	46	247	47
rect	246	49	247	50
rect	246	52	247	53
rect	246	55	247	56
rect	246	58	247	59
rect	246	61	247	62
rect	246	64	247	65
rect	246	67	247	68
rect	246	70	247	71
rect	246	73	247	74
rect	246	76	247	77
rect	246	79	247	80
rect	246	82	247	83
rect	246	85	247	86
rect	246	88	247	89
rect	246	94	247	95
rect	246	97	247	98
rect	246	100	247	101
rect	246	103	247	104
rect	246	106	247	107
rect	246	109	247	110
rect	246	115	247	116
rect	246	118	247	119
rect	246	124	247	125
rect	246	127	247	128
rect	246	133	247	134
rect	246	136	247	137
rect	246	139	247	140
rect	246	142	247	143
rect	246	145	247	146
rect	246	148	247	149
rect	246	151	247	152
rect	246	154	247	155
rect	246	157	247	158
rect	246	160	247	161
rect	246	163	247	164
rect	246	166	247	167
rect	246	169	247	170
rect	246	172	247	173
rect	246	175	247	176
rect	246	178	247	179
rect	246	181	247	182
rect	246	184	247	185
rect	246	187	247	188
rect	246	193	247	194
rect	246	196	247	197
rect	246	199	247	200
rect	246	202	247	203
rect	246	205	247	206
rect	246	208	247	209
rect	246	211	247	212
rect	246	214	247	215
rect	246	217	247	218
rect	246	220	247	221
rect	246	223	247	224
rect	246	226	247	227
rect	246	229	247	230
rect	246	238	247	239
rect	246	244	247	245
rect	246	247	247	248
rect	246	250	247	251
rect	247	7	248	8
rect	247	10	248	11
rect	247	13	248	14
rect	247	16	248	17
rect	247	19	248	20
rect	247	22	248	23
rect	247	25	248	26
rect	247	28	248	29
rect	247	31	248	32
rect	247	34	248	35
rect	247	37	248	38
rect	247	40	248	41
rect	247	43	248	44
rect	247	46	248	47
rect	247	49	248	50
rect	247	52	248	53
rect	247	55	248	56
rect	247	58	248	59
rect	247	61	248	62
rect	247	64	248	65
rect	247	67	248	68
rect	247	70	248	71
rect	247	73	248	74
rect	247	76	248	77
rect	247	79	248	80
rect	247	82	248	83
rect	247	85	248	86
rect	247	88	248	89
rect	247	94	248	95
rect	247	97	248	98
rect	247	100	248	101
rect	247	103	248	104
rect	247	106	248	107
rect	247	109	248	110
rect	247	115	248	116
rect	247	118	248	119
rect	247	124	248	125
rect	247	127	248	128
rect	247	133	248	134
rect	247	136	248	137
rect	247	139	248	140
rect	247	142	248	143
rect	247	145	248	146
rect	247	148	248	149
rect	247	151	248	152
rect	247	154	248	155
rect	247	157	248	158
rect	247	160	248	161
rect	247	163	248	164
rect	247	166	248	167
rect	247	169	248	170
rect	247	172	248	173
rect	247	175	248	176
rect	247	178	248	179
rect	247	181	248	182
rect	247	184	248	185
rect	247	187	248	188
rect	247	193	248	194
rect	247	196	248	197
rect	247	199	248	200
rect	247	202	248	203
rect	247	205	248	206
rect	247	208	248	209
rect	247	211	248	212
rect	247	214	248	215
rect	247	217	248	218
rect	247	220	248	221
rect	247	223	248	224
rect	247	226	248	227
rect	247	229	248	230
rect	247	238	248	239
rect	247	244	248	245
rect	247	247	248	248
rect	247	250	248	251
rect	248	7	249	8
rect	248	10	249	11
rect	248	13	249	14
rect	248	16	249	17
rect	248	19	249	20
rect	248	22	249	23
rect	248	25	249	26
rect	248	28	249	29
rect	248	31	249	32
rect	248	34	249	35
rect	248	37	249	38
rect	248	40	249	41
rect	248	43	249	44
rect	248	46	249	47
rect	248	49	249	50
rect	248	52	249	53
rect	248	55	249	56
rect	248	58	249	59
rect	248	61	249	62
rect	248	64	249	65
rect	248	67	249	68
rect	248	70	249	71
rect	248	73	249	74
rect	248	76	249	77
rect	248	79	249	80
rect	248	82	249	83
rect	248	85	249	86
rect	248	88	249	89
rect	248	94	249	95
rect	248	97	249	98
rect	248	100	249	101
rect	248	103	249	104
rect	248	106	249	107
rect	248	109	249	110
rect	248	115	249	116
rect	248	118	249	119
rect	248	124	249	125
rect	248	127	249	128
rect	248	133	249	134
rect	248	136	249	137
rect	248	139	249	140
rect	248	142	249	143
rect	248	145	249	146
rect	248	148	249	149
rect	248	151	249	152
rect	248	154	249	155
rect	248	157	249	158
rect	248	160	249	161
rect	248	163	249	164
rect	248	166	249	167
rect	248	169	249	170
rect	248	172	249	173
rect	248	175	249	176
rect	248	178	249	179
rect	248	181	249	182
rect	248	184	249	185
rect	248	187	249	188
rect	248	193	249	194
rect	248	196	249	197
rect	248	199	249	200
rect	248	202	249	203
rect	248	205	249	206
rect	248	208	249	209
rect	248	211	249	212
rect	248	214	249	215
rect	248	217	249	218
rect	248	220	249	221
rect	248	223	249	224
rect	248	226	249	227
rect	248	229	249	230
rect	248	238	249	239
rect	248	244	249	245
rect	248	247	249	248
rect	248	250	249	251
rect	249	7	250	8
rect	249	10	250	11
rect	249	13	250	14
rect	249	16	250	17
rect	249	19	250	20
rect	249	22	250	23
rect	249	25	250	26
rect	249	28	250	29
rect	249	31	250	32
rect	249	34	250	35
rect	249	37	250	38
rect	249	40	250	41
rect	249	43	250	44
rect	249	46	250	47
rect	249	49	250	50
rect	249	52	250	53
rect	249	55	250	56
rect	249	58	250	59
rect	249	61	250	62
rect	249	64	250	65
rect	249	67	250	68
rect	249	70	250	71
rect	249	73	250	74
rect	249	76	250	77
rect	249	79	250	80
rect	249	82	250	83
rect	249	85	250	86
rect	249	88	250	89
rect	249	94	250	95
rect	249	97	250	98
rect	249	100	250	101
rect	249	103	250	104
rect	249	106	250	107
rect	249	109	250	110
rect	249	115	250	116
rect	249	118	250	119
rect	249	124	250	125
rect	249	127	250	128
rect	249	133	250	134
rect	249	136	250	137
rect	249	139	250	140
rect	249	142	250	143
rect	249	145	250	146
rect	249	148	250	149
rect	249	151	250	152
rect	249	154	250	155
rect	249	157	250	158
rect	249	160	250	161
rect	249	163	250	164
rect	249	166	250	167
rect	249	169	250	170
rect	249	172	250	173
rect	249	175	250	176
rect	249	178	250	179
rect	249	181	250	182
rect	249	184	250	185
rect	249	187	250	188
rect	249	193	250	194
rect	249	196	250	197
rect	249	199	250	200
rect	249	202	250	203
rect	249	205	250	206
rect	249	208	250	209
rect	249	211	250	212
rect	249	214	250	215
rect	249	217	250	218
rect	249	220	250	221
rect	249	223	250	224
rect	249	226	250	227
rect	249	229	250	230
rect	249	238	250	239
rect	249	244	250	245
rect	249	247	250	248
rect	249	250	250	251
rect	250	7	251	8
rect	250	10	251	11
rect	250	13	251	14
rect	250	16	251	17
rect	250	19	251	20
rect	250	22	251	23
rect	250	25	251	26
rect	250	28	251	29
rect	250	31	251	32
rect	250	34	251	35
rect	250	37	251	38
rect	250	40	251	41
rect	250	43	251	44
rect	250	46	251	47
rect	250	49	251	50
rect	250	52	251	53
rect	250	55	251	56
rect	250	58	251	59
rect	250	61	251	62
rect	250	64	251	65
rect	250	67	251	68
rect	250	70	251	71
rect	250	73	251	74
rect	250	76	251	77
rect	250	79	251	80
rect	250	82	251	83
rect	250	85	251	86
rect	250	88	251	89
rect	250	94	251	95
rect	250	97	251	98
rect	250	100	251	101
rect	250	103	251	104
rect	250	106	251	107
rect	250	109	251	110
rect	250	115	251	116
rect	250	118	251	119
rect	250	124	251	125
rect	250	127	251	128
rect	250	133	251	134
rect	250	136	251	137
rect	250	139	251	140
rect	250	142	251	143
rect	250	145	251	146
rect	250	148	251	149
rect	250	151	251	152
rect	250	157	251	158
rect	250	160	251	161
rect	250	163	251	164
rect	250	166	251	167
rect	250	169	251	170
rect	250	172	251	173
rect	250	175	251	176
rect	250	178	251	179
rect	250	181	251	182
rect	250	184	251	185
rect	250	187	251	188
rect	250	193	251	194
rect	250	196	251	197
rect	250	199	251	200
rect	250	202	251	203
rect	250	205	251	206
rect	250	208	251	209
rect	250	211	251	212
rect	250	214	251	215
rect	250	217	251	218
rect	250	220	251	221
rect	250	223	251	224
rect	250	226	251	227
rect	250	229	251	230
rect	250	238	251	239
rect	250	247	251	248
rect	251	7	252	8
rect	251	10	252	11
rect	251	13	252	14
rect	251	16	252	17
rect	251	19	252	20
rect	251	22	252	23
rect	251	25	252	26
rect	251	28	252	29
rect	251	31	252	32
rect	251	34	252	35
rect	251	37	252	38
rect	251	40	252	41
rect	251	43	252	44
rect	251	46	252	47
rect	251	49	252	50
rect	251	52	252	53
rect	251	55	252	56
rect	251	58	252	59
rect	251	61	252	62
rect	251	64	252	65
rect	251	67	252	68
rect	251	70	252	71
rect	251	73	252	74
rect	251	76	252	77
rect	251	79	252	80
rect	251	82	252	83
rect	251	85	252	86
rect	251	88	252	89
rect	251	94	252	95
rect	251	97	252	98
rect	251	100	252	101
rect	251	103	252	104
rect	251	106	252	107
rect	251	109	252	110
rect	251	115	252	116
rect	251	118	252	119
rect	251	124	252	125
rect	251	127	252	128
rect	251	133	252	134
rect	251	136	252	137
rect	251	139	252	140
rect	251	142	252	143
rect	251	145	252	146
rect	251	148	252	149
rect	251	151	252	152
rect	251	157	252	158
rect	251	160	252	161
rect	251	163	252	164
rect	251	166	252	167
rect	251	169	252	170
rect	251	172	252	173
rect	251	175	252	176
rect	251	178	252	179
rect	251	181	252	182
rect	251	184	252	185
rect	251	187	252	188
rect	251	193	252	194
rect	251	196	252	197
rect	251	199	252	200
rect	251	202	252	203
rect	251	205	252	206
rect	251	208	252	209
rect	251	211	252	212
rect	251	214	252	215
rect	251	217	252	218
rect	251	220	252	221
rect	251	223	252	224
rect	251	226	252	227
rect	251	229	252	230
rect	251	235	252	236
rect	251	238	252	239
rect	251	247	252	248
rect	252	7	253	8
rect	252	10	253	11
rect	252	13	253	14
rect	252	16	253	17
rect	252	19	253	20
rect	252	22	253	23
rect	252	25	253	26
rect	252	28	253	29
rect	252	31	253	32
rect	252	34	253	35
rect	252	37	253	38
rect	252	40	253	41
rect	252	43	253	44
rect	252	46	253	47
rect	252	49	253	50
rect	252	52	253	53
rect	252	55	253	56
rect	252	58	253	59
rect	252	61	253	62
rect	252	64	253	65
rect	252	67	253	68
rect	252	70	253	71
rect	252	73	253	74
rect	252	76	253	77
rect	252	79	253	80
rect	252	82	253	83
rect	252	85	253	86
rect	252	88	253	89
rect	252	94	253	95
rect	252	97	253	98
rect	252	100	253	101
rect	252	103	253	104
rect	252	106	253	107
rect	252	109	253	110
rect	252	115	253	116
rect	252	118	253	119
rect	252	124	253	125
rect	252	127	253	128
rect	252	133	253	134
rect	252	136	253	137
rect	252	139	253	140
rect	252	142	253	143
rect	252	145	253	146
rect	252	148	253	149
rect	252	151	253	152
rect	252	157	253	158
rect	252	160	253	161
rect	252	163	253	164
rect	252	166	253	167
rect	252	169	253	170
rect	252	172	253	173
rect	252	175	253	176
rect	252	178	253	179
rect	252	181	253	182
rect	252	184	253	185
rect	252	187	253	188
rect	252	193	253	194
rect	252	196	253	197
rect	252	199	253	200
rect	252	202	253	203
rect	252	205	253	206
rect	252	208	253	209
rect	252	211	253	212
rect	252	214	253	215
rect	252	217	253	218
rect	252	220	253	221
rect	252	223	253	224
rect	252	226	253	227
rect	252	229	253	230
rect	252	235	253	236
rect	252	238	253	239
rect	252	247	253	248
rect	253	7	254	8
rect	253	10	254	11
rect	253	13	254	14
rect	253	16	254	17
rect	253	19	254	20
rect	253	22	254	23
rect	253	25	254	26
rect	253	28	254	29
rect	253	31	254	32
rect	253	34	254	35
rect	253	37	254	38
rect	253	40	254	41
rect	253	43	254	44
rect	253	46	254	47
rect	253	49	254	50
rect	253	52	254	53
rect	253	55	254	56
rect	253	58	254	59
rect	253	61	254	62
rect	253	64	254	65
rect	253	67	254	68
rect	253	70	254	71
rect	253	73	254	74
rect	253	76	254	77
rect	253	79	254	80
rect	253	82	254	83
rect	253	85	254	86
rect	253	88	254	89
rect	253	94	254	95
rect	253	97	254	98
rect	253	100	254	101
rect	253	103	254	104
rect	253	106	254	107
rect	253	109	254	110
rect	253	115	254	116
rect	253	118	254	119
rect	253	124	254	125
rect	253	127	254	128
rect	253	133	254	134
rect	253	136	254	137
rect	253	139	254	140
rect	253	142	254	143
rect	253	145	254	146
rect	253	148	254	149
rect	253	151	254	152
rect	253	157	254	158
rect	253	160	254	161
rect	253	163	254	164
rect	253	166	254	167
rect	253	169	254	170
rect	253	172	254	173
rect	253	175	254	176
rect	253	178	254	179
rect	253	181	254	182
rect	253	184	254	185
rect	253	187	254	188
rect	253	193	254	194
rect	253	196	254	197
rect	253	199	254	200
rect	253	202	254	203
rect	253	205	254	206
rect	253	208	254	209
rect	253	211	254	212
rect	253	214	254	215
rect	253	217	254	218
rect	253	220	254	221
rect	253	223	254	224
rect	253	226	254	227
rect	253	229	254	230
rect	253	238	254	239
rect	253	247	254	248
rect	254	7	255	8
rect	254	10	255	11
rect	254	13	255	14
rect	254	16	255	17
rect	254	19	255	20
rect	254	22	255	23
rect	254	25	255	26
rect	254	28	255	29
rect	254	31	255	32
rect	254	34	255	35
rect	254	37	255	38
rect	254	40	255	41
rect	254	43	255	44
rect	254	46	255	47
rect	254	49	255	50
rect	254	52	255	53
rect	254	55	255	56
rect	254	58	255	59
rect	254	61	255	62
rect	254	64	255	65
rect	254	67	255	68
rect	254	70	255	71
rect	254	73	255	74
rect	254	76	255	77
rect	254	79	255	80
rect	254	82	255	83
rect	254	85	255	86
rect	254	88	255	89
rect	254	94	255	95
rect	254	97	255	98
rect	254	100	255	101
rect	254	103	255	104
rect	254	106	255	107
rect	254	109	255	110
rect	254	115	255	116
rect	254	118	255	119
rect	254	124	255	125
rect	254	127	255	128
rect	254	133	255	134
rect	254	136	255	137
rect	254	139	255	140
rect	254	142	255	143
rect	254	145	255	146
rect	254	148	255	149
rect	254	151	255	152
rect	254	154	255	155
rect	254	157	255	158
rect	254	160	255	161
rect	254	163	255	164
rect	254	166	255	167
rect	254	169	255	170
rect	254	172	255	173
rect	254	175	255	176
rect	254	178	255	179
rect	254	181	255	182
rect	254	184	255	185
rect	254	187	255	188
rect	254	193	255	194
rect	254	196	255	197
rect	254	199	255	200
rect	254	202	255	203
rect	254	205	255	206
rect	254	208	255	209
rect	254	211	255	212
rect	254	214	255	215
rect	254	217	255	218
rect	254	220	255	221
rect	254	223	255	224
rect	254	226	255	227
rect	254	229	255	230
rect	254	238	255	239
rect	254	247	255	248
rect	254	250	255	251
rect	254	256	255	257
rect	255	7	256	8
rect	255	10	256	11
rect	255	13	256	14
rect	255	16	256	17
rect	255	19	256	20
rect	255	22	256	23
rect	255	25	256	26
rect	255	28	256	29
rect	255	31	256	32
rect	255	34	256	35
rect	255	37	256	38
rect	255	40	256	41
rect	255	43	256	44
rect	255	46	256	47
rect	255	49	256	50
rect	255	52	256	53
rect	255	55	256	56
rect	255	58	256	59
rect	255	61	256	62
rect	255	64	256	65
rect	255	67	256	68
rect	255	79	256	80
rect	255	82	256	83
rect	255	85	256	86
rect	255	88	256	89
rect	255	97	256	98
rect	255	100	256	101
rect	255	103	256	104
rect	255	109	256	110
rect	255	115	256	116
rect	255	118	256	119
rect	255	124	256	125
rect	255	127	256	128
rect	255	133	256	134
rect	255	136	256	137
rect	255	139	256	140
rect	255	142	256	143
rect	255	148	256	149
rect	255	151	256	152
rect	255	157	256	158
rect	255	160	256	161
rect	255	163	256	164
rect	255	166	256	167
rect	255	169	256	170
rect	255	172	256	173
rect	255	175	256	176
rect	255	178	256	179
rect	255	181	256	182
rect	255	184	256	185
rect	255	187	256	188
rect	255	193	256	194
rect	255	196	256	197
rect	255	199	256	200
rect	255	202	256	203
rect	255	205	256	206
rect	255	208	256	209
rect	255	211	256	212
rect	255	217	256	218
rect	255	220	256	221
rect	255	223	256	224
rect	255	238	256	239
rect	256	7	257	8
rect	256	10	257	11
rect	256	13	257	14
rect	256	16	257	17
rect	256	19	257	20
rect	256	22	257	23
rect	256	25	257	26
rect	256	28	257	29
rect	256	31	257	32
rect	256	34	257	35
rect	256	37	257	38
rect	256	40	257	41
rect	256	43	257	44
rect	256	46	257	47
rect	256	49	257	50
rect	256	52	257	53
rect	256	55	257	56
rect	256	58	257	59
rect	256	61	257	62
rect	256	64	257	65
rect	256	67	257	68
rect	256	79	257	80
rect	256	82	257	83
rect	256	85	257	86
rect	256	88	257	89
rect	256	97	257	98
rect	256	100	257	101
rect	256	103	257	104
rect	256	109	257	110
rect	256	115	257	116
rect	256	118	257	119
rect	256	124	257	125
rect	256	127	257	128
rect	256	133	257	134
rect	256	136	257	137
rect	256	139	257	140
rect	256	142	257	143
rect	256	148	257	149
rect	256	151	257	152
rect	256	157	257	158
rect	256	160	257	161
rect	256	163	257	164
rect	256	166	257	167
rect	256	169	257	170
rect	256	172	257	173
rect	256	175	257	176
rect	256	178	257	179
rect	256	181	257	182
rect	256	184	257	185
rect	256	187	257	188
rect	256	193	257	194
rect	256	196	257	197
rect	256	199	257	200
rect	256	202	257	203
rect	256	205	257	206
rect	256	208	257	209
rect	256	211	257	212
rect	256	217	257	218
rect	256	220	257	221
rect	256	223	257	224
rect	256	238	257	239
rect	257	7	258	8
rect	257	10	258	11
rect	257	13	258	14
rect	257	16	258	17
rect	257	19	258	20
rect	257	22	258	23
rect	257	25	258	26
rect	257	28	258	29
rect	257	31	258	32
rect	257	34	258	35
rect	257	37	258	38
rect	257	40	258	41
rect	257	43	258	44
rect	257	46	258	47
rect	257	49	258	50
rect	257	52	258	53
rect	257	55	258	56
rect	257	58	258	59
rect	257	61	258	62
rect	257	64	258	65
rect	257	67	258	68
rect	257	79	258	80
rect	257	82	258	83
rect	257	85	258	86
rect	257	88	258	89
rect	257	97	258	98
rect	257	100	258	101
rect	257	103	258	104
rect	257	109	258	110
rect	257	115	258	116
rect	257	118	258	119
rect	257	124	258	125
rect	257	127	258	128
rect	257	133	258	134
rect	257	136	258	137
rect	257	139	258	140
rect	257	142	258	143
rect	257	148	258	149
rect	257	151	258	152
rect	257	157	258	158
rect	257	160	258	161
rect	257	163	258	164
rect	257	166	258	167
rect	257	169	258	170
rect	257	172	258	173
rect	257	175	258	176
rect	257	178	258	179
rect	257	181	258	182
rect	257	184	258	185
rect	257	187	258	188
rect	257	193	258	194
rect	257	196	258	197
rect	257	199	258	200
rect	257	202	258	203
rect	257	205	258	206
rect	257	208	258	209
rect	257	211	258	212
rect	257	217	258	218
rect	257	220	258	221
rect	257	223	258	224
rect	257	238	258	239
rect	258	7	259	8
rect	258	10	259	11
rect	258	13	259	14
rect	258	16	259	17
rect	258	19	259	20
rect	258	22	259	23
rect	258	25	259	26
rect	258	28	259	29
rect	258	31	259	32
rect	258	34	259	35
rect	258	37	259	38
rect	258	40	259	41
rect	258	43	259	44
rect	258	46	259	47
rect	258	49	259	50
rect	258	52	259	53
rect	258	55	259	56
rect	258	58	259	59
rect	258	61	259	62
rect	258	64	259	65
rect	258	67	259	68
rect	258	79	259	80
rect	258	82	259	83
rect	258	85	259	86
rect	258	88	259	89
rect	258	97	259	98
rect	258	100	259	101
rect	258	103	259	104
rect	258	109	259	110
rect	258	115	259	116
rect	258	118	259	119
rect	258	124	259	125
rect	258	127	259	128
rect	258	133	259	134
rect	258	136	259	137
rect	258	139	259	140
rect	258	142	259	143
rect	258	148	259	149
rect	258	151	259	152
rect	258	157	259	158
rect	258	160	259	161
rect	258	163	259	164
rect	258	166	259	167
rect	258	169	259	170
rect	258	172	259	173
rect	258	175	259	176
rect	258	178	259	179
rect	258	181	259	182
rect	258	184	259	185
rect	258	187	259	188
rect	258	193	259	194
rect	258	196	259	197
rect	258	199	259	200
rect	258	202	259	203
rect	258	205	259	206
rect	258	208	259	209
rect	258	211	259	212
rect	258	217	259	218
rect	258	220	259	221
rect	258	223	259	224
rect	258	238	259	239
rect	259	7	260	8
rect	259	10	260	11
rect	259	13	260	14
rect	259	16	260	17
rect	259	19	260	20
rect	259	22	260	23
rect	259	25	260	26
rect	259	28	260	29
rect	259	31	260	32
rect	259	34	260	35
rect	259	37	260	38
rect	259	40	260	41
rect	259	43	260	44
rect	259	46	260	47
rect	259	49	260	50
rect	259	52	260	53
rect	259	55	260	56
rect	259	58	260	59
rect	259	61	260	62
rect	259	64	260	65
rect	259	67	260	68
rect	259	79	260	80
rect	259	82	260	83
rect	259	85	260	86
rect	259	88	260	89
rect	259	100	260	101
rect	259	103	260	104
rect	259	109	260	110
rect	259	115	260	116
rect	259	118	260	119
rect	259	124	260	125
rect	259	127	260	128
rect	259	133	260	134
rect	259	136	260	137
rect	259	139	260	140
rect	259	142	260	143
rect	259	148	260	149
rect	259	151	260	152
rect	259	157	260	158
rect	259	160	260	161
rect	259	163	260	164
rect	259	166	260	167
rect	259	169	260	170
rect	259	172	260	173
rect	259	175	260	176
rect	259	178	260	179
rect	259	181	260	182
rect	259	184	260	185
rect	259	187	260	188
rect	259	193	260	194
rect	259	196	260	197
rect	259	199	260	200
rect	259	202	260	203
rect	259	205	260	206
rect	259	208	260	209
rect	259	211	260	212
rect	259	217	260	218
rect	259	223	260	224
rect	259	238	260	239
rect	260	7	261	8
rect	260	10	261	11
rect	260	13	261	14
rect	260	16	261	17
rect	260	19	261	20
rect	260	22	261	23
rect	260	25	261	26
rect	260	28	261	29
rect	260	31	261	32
rect	260	34	261	35
rect	260	37	261	38
rect	260	40	261	41
rect	260	43	261	44
rect	260	46	261	47
rect	260	49	261	50
rect	260	52	261	53
rect	260	55	261	56
rect	260	58	261	59
rect	260	61	261	62
rect	260	64	261	65
rect	260	67	261	68
rect	260	79	261	80
rect	260	82	261	83
rect	260	85	261	86
rect	260	88	261	89
rect	260	100	261	101
rect	260	103	261	104
rect	260	109	261	110
rect	260	115	261	116
rect	260	118	261	119
rect	260	124	261	125
rect	260	127	261	128
rect	260	133	261	134
rect	260	136	261	137
rect	260	139	261	140
rect	260	142	261	143
rect	260	148	261	149
rect	260	151	261	152
rect	260	157	261	158
rect	260	160	261	161
rect	260	163	261	164
rect	260	166	261	167
rect	260	169	261	170
rect	260	172	261	173
rect	260	175	261	176
rect	260	178	261	179
rect	260	181	261	182
rect	260	184	261	185
rect	260	187	261	188
rect	260	193	261	194
rect	260	196	261	197
rect	260	199	261	200
rect	260	202	261	203
rect	260	205	261	206
rect	260	208	261	209
rect	260	211	261	212
rect	260	217	261	218
rect	260	223	261	224
rect	260	238	261	239
rect	261	7	262	8
rect	261	10	262	11
rect	261	13	262	14
rect	261	16	262	17
rect	261	19	262	20
rect	261	22	262	23
rect	261	25	262	26
rect	261	28	262	29
rect	261	31	262	32
rect	261	34	262	35
rect	261	37	262	38
rect	261	40	262	41
rect	261	43	262	44
rect	261	46	262	47
rect	261	49	262	50
rect	261	52	262	53
rect	261	55	262	56
rect	261	58	262	59
rect	261	61	262	62
rect	261	64	262	65
rect	261	67	262	68
rect	261	79	262	80
rect	261	82	262	83
rect	261	85	262	86
rect	261	88	262	89
rect	261	100	262	101
rect	261	103	262	104
rect	261	109	262	110
rect	261	115	262	116
rect	261	118	262	119
rect	261	124	262	125
rect	261	127	262	128
rect	261	133	262	134
rect	261	136	262	137
rect	261	139	262	140
rect	261	142	262	143
rect	261	148	262	149
rect	261	151	262	152
rect	261	157	262	158
rect	261	160	262	161
rect	261	163	262	164
rect	261	166	262	167
rect	261	169	262	170
rect	261	172	262	173
rect	261	175	262	176
rect	261	178	262	179
rect	261	181	262	182
rect	261	184	262	185
rect	261	187	262	188
rect	261	193	262	194
rect	261	196	262	197
rect	261	199	262	200
rect	261	202	262	203
rect	261	205	262	206
rect	261	208	262	209
rect	261	211	262	212
rect	261	217	262	218
rect	261	223	262	224
rect	261	238	262	239
rect	262	7	263	8
rect	262	10	263	11
rect	262	13	263	14
rect	262	16	263	17
rect	262	19	263	20
rect	262	22	263	23
rect	262	25	263	26
rect	262	28	263	29
rect	262	31	263	32
rect	262	34	263	35
rect	262	37	263	38
rect	262	40	263	41
rect	262	43	263	44
rect	262	46	263	47
rect	262	49	263	50
rect	262	52	263	53
rect	262	55	263	56
rect	262	58	263	59
rect	262	61	263	62
rect	262	64	263	65
rect	262	67	263	68
rect	262	79	263	80
rect	262	82	263	83
rect	262	85	263	86
rect	262	88	263	89
rect	262	100	263	101
rect	262	103	263	104
rect	262	109	263	110
rect	262	115	263	116
rect	262	118	263	119
rect	262	124	263	125
rect	262	127	263	128
rect	262	133	263	134
rect	262	136	263	137
rect	262	139	263	140
rect	262	142	263	143
rect	262	148	263	149
rect	262	151	263	152
rect	262	157	263	158
rect	262	160	263	161
rect	262	163	263	164
rect	262	166	263	167
rect	262	169	263	170
rect	262	172	263	173
rect	262	175	263	176
rect	262	178	263	179
rect	262	181	263	182
rect	262	184	263	185
rect	262	187	263	188
rect	262	193	263	194
rect	262	196	263	197
rect	262	199	263	200
rect	262	202	263	203
rect	262	205	263	206
rect	262	208	263	209
rect	262	211	263	212
rect	262	217	263	218
rect	262	223	263	224
rect	262	238	263	239
rect	263	7	264	8
rect	263	10	264	11
rect	263	13	264	14
rect	263	16	264	17
rect	263	19	264	20
rect	263	22	264	23
rect	263	25	264	26
rect	263	28	264	29
rect	263	31	264	32
rect	263	34	264	35
rect	263	37	264	38
rect	263	40	264	41
rect	263	43	264	44
rect	263	46	264	47
rect	263	49	264	50
rect	263	52	264	53
rect	263	55	264	56
rect	263	58	264	59
rect	263	61	264	62
rect	263	64	264	65
rect	263	67	264	68
rect	263	79	264	80
rect	263	82	264	83
rect	263	85	264	86
rect	263	88	264	89
rect	263	97	264	98
rect	263	100	264	101
rect	263	103	264	104
rect	263	106	264	107
rect	263	109	264	110
rect	263	115	264	116
rect	263	118	264	119
rect	263	124	264	125
rect	263	127	264	128
rect	263	133	264	134
rect	263	136	264	137
rect	263	139	264	140
rect	263	142	264	143
rect	263	148	264	149
rect	263	151	264	152
rect	263	157	264	158
rect	263	160	264	161
rect	263	163	264	164
rect	263	166	264	167
rect	263	169	264	170
rect	263	172	264	173
rect	263	175	264	176
rect	263	178	264	179
rect	263	181	264	182
rect	263	184	264	185
rect	263	187	264	188
rect	263	193	264	194
rect	263	196	264	197
rect	263	199	264	200
rect	263	202	264	203
rect	263	205	264	206
rect	263	208	264	209
rect	263	211	264	212
rect	263	217	264	218
rect	263	220	264	221
rect	263	223	264	224
rect	263	226	264	227
rect	263	238	264	239
rect	264	7	265	8
rect	264	10	265	11
rect	264	13	265	14
rect	264	16	265	17
rect	264	19	265	20
rect	264	22	265	23
rect	264	25	265	26
rect	264	28	265	29
rect	264	31	265	32
rect	264	34	265	35
rect	264	37	265	38
rect	264	40	265	41
rect	264	43	265	44
rect	264	46	265	47
rect	264	49	265	50
rect	264	52	265	53
rect	264	55	265	56
rect	264	58	265	59
rect	264	61	265	62
rect	264	64	265	65
rect	264	79	265	80
rect	264	82	265	83
rect	264	85	265	86
rect	264	88	265	89
rect	264	103	265	104
rect	264	109	265	110
rect	264	115	265	116
rect	264	118	265	119
rect	264	124	265	125
rect	264	127	265	128
rect	264	133	265	134
rect	264	136	265	137
rect	264	139	265	140
rect	264	142	265	143
rect	264	148	265	149
rect	264	151	265	152
rect	264	157	265	158
rect	264	160	265	161
rect	264	163	265	164
rect	264	166	265	167
rect	264	169	265	170
rect	264	172	265	173
rect	264	175	265	176
rect	264	178	265	179
rect	264	181	265	182
rect	264	184	265	185
rect	264	187	265	188
rect	264	193	265	194
rect	264	196	265	197
rect	264	199	265	200
rect	264	202	265	203
rect	264	211	265	212
rect	264	217	265	218
rect	264	238	265	239
rect	265	7	266	8
rect	265	10	266	11
rect	265	13	266	14
rect	265	16	266	17
rect	265	19	266	20
rect	265	22	266	23
rect	265	25	266	26
rect	265	28	266	29
rect	265	31	266	32
rect	265	34	266	35
rect	265	37	266	38
rect	265	40	266	41
rect	265	43	266	44
rect	265	46	266	47
rect	265	49	266	50
rect	265	52	266	53
rect	265	55	266	56
rect	265	58	266	59
rect	265	61	266	62
rect	265	64	266	65
rect	265	79	266	80
rect	265	82	266	83
rect	265	85	266	86
rect	265	88	266	89
rect	265	103	266	104
rect	265	109	266	110
rect	265	115	266	116
rect	265	118	266	119
rect	265	124	266	125
rect	265	127	266	128
rect	265	133	266	134
rect	265	136	266	137
rect	265	139	266	140
rect	265	142	266	143
rect	265	148	266	149
rect	265	151	266	152
rect	265	157	266	158
rect	265	160	266	161
rect	265	163	266	164
rect	265	166	266	167
rect	265	169	266	170
rect	265	172	266	173
rect	265	175	266	176
rect	265	178	266	179
rect	265	181	266	182
rect	265	184	266	185
rect	265	187	266	188
rect	265	193	266	194
rect	265	196	266	197
rect	265	199	266	200
rect	265	202	266	203
rect	265	211	266	212
rect	265	217	266	218
rect	265	238	266	239
rect	266	7	267	8
rect	266	10	267	11
rect	266	13	267	14
rect	266	16	267	17
rect	266	19	267	20
rect	266	22	267	23
rect	266	25	267	26
rect	266	28	267	29
rect	266	31	267	32
rect	266	34	267	35
rect	266	37	267	38
rect	266	40	267	41
rect	266	43	267	44
rect	266	46	267	47
rect	266	49	267	50
rect	266	52	267	53
rect	266	55	267	56
rect	266	58	267	59
rect	266	61	267	62
rect	266	64	267	65
rect	266	79	267	80
rect	266	82	267	83
rect	266	85	267	86
rect	266	88	267	89
rect	266	103	267	104
rect	266	109	267	110
rect	266	115	267	116
rect	266	118	267	119
rect	266	124	267	125
rect	266	127	267	128
rect	266	133	267	134
rect	266	136	267	137
rect	266	139	267	140
rect	266	142	267	143
rect	266	148	267	149
rect	266	151	267	152
rect	266	157	267	158
rect	266	160	267	161
rect	266	163	267	164
rect	266	166	267	167
rect	266	169	267	170
rect	266	172	267	173
rect	266	175	267	176
rect	266	178	267	179
rect	266	181	267	182
rect	266	184	267	185
rect	266	187	267	188
rect	266	193	267	194
rect	266	196	267	197
rect	266	199	267	200
rect	266	202	267	203
rect	266	211	267	212
rect	266	217	267	218
rect	266	238	267	239
rect	267	7	268	8
rect	267	10	268	11
rect	267	13	268	14
rect	267	16	268	17
rect	267	19	268	20
rect	267	22	268	23
rect	267	25	268	26
rect	267	28	268	29
rect	267	31	268	32
rect	267	34	268	35
rect	267	37	268	38
rect	267	40	268	41
rect	267	43	268	44
rect	267	46	268	47
rect	267	49	268	50
rect	267	52	268	53
rect	267	55	268	56
rect	267	58	268	59
rect	267	61	268	62
rect	267	64	268	65
rect	267	79	268	80
rect	267	82	268	83
rect	267	85	268	86
rect	267	88	268	89
rect	267	103	268	104
rect	267	109	268	110
rect	267	115	268	116
rect	267	118	268	119
rect	267	124	268	125
rect	267	127	268	128
rect	267	133	268	134
rect	267	136	268	137
rect	267	139	268	140
rect	267	142	268	143
rect	267	148	268	149
rect	267	151	268	152
rect	267	157	268	158
rect	267	160	268	161
rect	267	163	268	164
rect	267	166	268	167
rect	267	169	268	170
rect	267	172	268	173
rect	267	175	268	176
rect	267	178	268	179
rect	267	181	268	182
rect	267	184	268	185
rect	267	187	268	188
rect	267	193	268	194
rect	267	196	268	197
rect	267	199	268	200
rect	267	202	268	203
rect	267	211	268	212
rect	267	217	268	218
rect	267	238	268	239
rect	268	7	269	8
rect	268	10	269	11
rect	268	13	269	14
rect	268	16	269	17
rect	268	19	269	20
rect	268	22	269	23
rect	268	25	269	26
rect	268	28	269	29
rect	268	31	269	32
rect	268	34	269	35
rect	268	37	269	38
rect	268	40	269	41
rect	268	43	269	44
rect	268	46	269	47
rect	268	49	269	50
rect	268	52	269	53
rect	268	55	269	56
rect	268	58	269	59
rect	268	61	269	62
rect	268	64	269	65
rect	268	79	269	80
rect	268	82	269	83
rect	268	85	269	86
rect	268	88	269	89
rect	268	103	269	104
rect	268	109	269	110
rect	268	115	269	116
rect	268	118	269	119
rect	268	124	269	125
rect	268	127	269	128
rect	268	133	269	134
rect	268	136	269	137
rect	268	139	269	140
rect	268	142	269	143
rect	268	148	269	149
rect	268	151	269	152
rect	268	157	269	158
rect	268	160	269	161
rect	268	163	269	164
rect	268	166	269	167
rect	268	169	269	170
rect	268	172	269	173
rect	268	175	269	176
rect	268	178	269	179
rect	268	181	269	182
rect	268	184	269	185
rect	268	187	269	188
rect	268	193	269	194
rect	268	196	269	197
rect	268	199	269	200
rect	268	202	269	203
rect	268	211	269	212
rect	268	217	269	218
rect	268	238	269	239
rect	269	7	270	8
rect	269	10	270	11
rect	269	13	270	14
rect	269	16	270	17
rect	269	19	270	20
rect	269	22	270	23
rect	269	25	270	26
rect	269	28	270	29
rect	269	31	270	32
rect	269	34	270	35
rect	269	37	270	38
rect	269	40	270	41
rect	269	43	270	44
rect	269	46	270	47
rect	269	49	270	50
rect	269	52	270	53
rect	269	55	270	56
rect	269	58	270	59
rect	269	61	270	62
rect	269	64	270	65
rect	269	79	270	80
rect	269	82	270	83
rect	269	85	270	86
rect	269	88	270	89
rect	269	103	270	104
rect	269	109	270	110
rect	269	115	270	116
rect	269	118	270	119
rect	269	124	270	125
rect	269	127	270	128
rect	269	133	270	134
rect	269	136	270	137
rect	269	139	270	140
rect	269	142	270	143
rect	269	148	270	149
rect	269	151	270	152
rect	269	157	270	158
rect	269	160	270	161
rect	269	163	270	164
rect	269	166	270	167
rect	269	169	270	170
rect	269	172	270	173
rect	269	175	270	176
rect	269	178	270	179
rect	269	181	270	182
rect	269	184	270	185
rect	269	187	270	188
rect	269	193	270	194
rect	269	196	270	197
rect	269	199	270	200
rect	269	202	270	203
rect	269	211	270	212
rect	269	217	270	218
rect	269	238	270	239
rect	270	7	271	8
rect	270	10	271	11
rect	270	13	271	14
rect	270	16	271	17
rect	270	19	271	20
rect	270	22	271	23
rect	270	25	271	26
rect	270	28	271	29
rect	270	31	271	32
rect	270	34	271	35
rect	270	37	271	38
rect	270	40	271	41
rect	270	43	271	44
rect	270	46	271	47
rect	270	49	271	50
rect	270	55	271	56
rect	270	58	271	59
rect	270	61	271	62
rect	270	64	271	65
rect	270	79	271	80
rect	270	82	271	83
rect	270	85	271	86
rect	270	88	271	89
rect	270	103	271	104
rect	270	109	271	110
rect	270	115	271	116
rect	270	118	271	119
rect	270	124	271	125
rect	270	127	271	128
rect	270	133	271	134
rect	270	136	271	137
rect	270	139	271	140
rect	270	142	271	143
rect	270	148	271	149
rect	270	151	271	152
rect	270	157	271	158
rect	270	160	271	161
rect	270	163	271	164
rect	270	166	271	167
rect	270	169	271	170
rect	270	172	271	173
rect	270	175	271	176
rect	270	178	271	179
rect	270	181	271	182
rect	270	184	271	185
rect	270	187	271	188
rect	270	196	271	197
rect	270	199	271	200
rect	270	202	271	203
rect	270	217	271	218
rect	270	238	271	239
rect	271	7	272	8
rect	271	10	272	11
rect	271	13	272	14
rect	271	16	272	17
rect	271	19	272	20
rect	271	22	272	23
rect	271	25	272	26
rect	271	28	272	29
rect	271	31	272	32
rect	271	34	272	35
rect	271	37	272	38
rect	271	40	272	41
rect	271	43	272	44
rect	271	46	272	47
rect	271	49	272	50
rect	271	55	272	56
rect	271	58	272	59
rect	271	61	272	62
rect	271	64	272	65
rect	271	79	272	80
rect	271	82	272	83
rect	271	85	272	86
rect	271	88	272	89
rect	271	103	272	104
rect	271	109	272	110
rect	271	115	272	116
rect	271	118	272	119
rect	271	124	272	125
rect	271	127	272	128
rect	271	133	272	134
rect	271	136	272	137
rect	271	139	272	140
rect	271	142	272	143
rect	271	148	272	149
rect	271	151	272	152
rect	271	157	272	158
rect	271	160	272	161
rect	271	163	272	164
rect	271	166	272	167
rect	271	169	272	170
rect	271	172	272	173
rect	271	175	272	176
rect	271	178	272	179
rect	271	181	272	182
rect	271	184	272	185
rect	271	187	272	188
rect	271	196	272	197
rect	271	199	272	200
rect	271	202	272	203
rect	271	217	272	218
rect	271	238	272	239
rect	272	7	273	8
rect	272	10	273	11
rect	272	13	273	14
rect	272	16	273	17
rect	272	19	273	20
rect	272	22	273	23
rect	272	25	273	26
rect	272	28	273	29
rect	272	31	273	32
rect	272	34	273	35
rect	272	37	273	38
rect	272	40	273	41
rect	272	43	273	44
rect	272	46	273	47
rect	272	49	273	50
rect	272	55	273	56
rect	272	58	273	59
rect	272	61	273	62
rect	272	64	273	65
rect	272	79	273	80
rect	272	82	273	83
rect	272	85	273	86
rect	272	88	273	89
rect	272	103	273	104
rect	272	109	273	110
rect	272	115	273	116
rect	272	118	273	119
rect	272	124	273	125
rect	272	127	273	128
rect	272	133	273	134
rect	272	136	273	137
rect	272	139	273	140
rect	272	142	273	143
rect	272	148	273	149
rect	272	151	273	152
rect	272	157	273	158
rect	272	160	273	161
rect	272	163	273	164
rect	272	166	273	167
rect	272	169	273	170
rect	272	172	273	173
rect	272	175	273	176
rect	272	178	273	179
rect	272	181	273	182
rect	272	184	273	185
rect	272	187	273	188
rect	272	193	273	194
rect	272	196	273	197
rect	272	199	273	200
rect	272	202	273	203
rect	272	217	273	218
rect	272	238	273	239
rect	273	7	274	8
rect	273	10	274	11
rect	273	13	274	14
rect	273	16	274	17
rect	273	19	274	20
rect	273	22	274	23
rect	273	25	274	26
rect	273	28	274	29
rect	273	31	274	32
rect	273	34	274	35
rect	273	37	274	38
rect	273	40	274	41
rect	273	43	274	44
rect	273	46	274	47
rect	273	49	274	50
rect	273	55	274	56
rect	273	58	274	59
rect	273	61	274	62
rect	273	64	274	65
rect	273	79	274	80
rect	273	82	274	83
rect	273	85	274	86
rect	273	88	274	89
rect	273	103	274	104
rect	273	109	274	110
rect	273	115	274	116
rect	273	118	274	119
rect	273	124	274	125
rect	273	127	274	128
rect	273	133	274	134
rect	273	136	274	137
rect	273	139	274	140
rect	273	142	274	143
rect	273	148	274	149
rect	273	151	274	152
rect	273	157	274	158
rect	273	160	274	161
rect	273	163	274	164
rect	273	166	274	167
rect	273	169	274	170
rect	273	172	274	173
rect	273	175	274	176
rect	273	178	274	179
rect	273	181	274	182
rect	273	184	274	185
rect	273	187	274	188
rect	273	193	274	194
rect	273	196	274	197
rect	273	199	274	200
rect	273	202	274	203
rect	273	217	274	218
rect	273	238	274	239
rect	274	7	275	8
rect	274	10	275	11
rect	274	13	275	14
rect	274	16	275	17
rect	274	19	275	20
rect	274	22	275	23
rect	274	25	275	26
rect	274	28	275	29
rect	274	31	275	32
rect	274	34	275	35
rect	274	37	275	38
rect	274	40	275	41
rect	274	43	275	44
rect	274	46	275	47
rect	274	49	275	50
rect	274	52	275	53
rect	274	55	275	56
rect	274	58	275	59
rect	274	61	275	62
rect	274	64	275	65
rect	274	79	275	80
rect	274	82	275	83
rect	274	85	275	86
rect	274	88	275	89
rect	274	103	275	104
rect	274	109	275	110
rect	274	115	275	116
rect	274	118	275	119
rect	274	124	275	125
rect	274	127	275	128
rect	274	133	275	134
rect	274	136	275	137
rect	274	139	275	140
rect	274	142	275	143
rect	274	148	275	149
rect	274	151	275	152
rect	274	157	275	158
rect	274	160	275	161
rect	274	163	275	164
rect	274	166	275	167
rect	274	169	275	170
rect	274	172	275	173
rect	274	175	275	176
rect	274	178	275	179
rect	274	181	275	182
rect	274	184	275	185
rect	274	187	275	188
rect	274	190	275	191
rect	274	193	275	194
rect	274	196	275	197
rect	274	199	275	200
rect	274	202	275	203
rect	274	211	275	212
rect	274	217	275	218
rect	274	238	275	239
rect	275	7	276	8
rect	275	10	276	11
rect	275	13	276	14
rect	275	16	276	17
rect	275	19	276	20
rect	275	22	276	23
rect	275	25	276	26
rect	275	28	276	29
rect	275	31	276	32
rect	275	34	276	35
rect	275	37	276	38
rect	275	40	276	41
rect	275	43	276	44
rect	275	46	276	47
rect	275	49	276	50
rect	275	55	276	56
rect	275	61	276	62
rect	275	64	276	65
rect	275	79	276	80
rect	275	82	276	83
rect	275	85	276	86
rect	275	88	276	89
rect	275	109	276	110
rect	275	115	276	116
rect	275	118	276	119
rect	275	124	276	125
rect	275	133	276	134
rect	275	136	276	137
rect	275	139	276	140
rect	275	148	276	149
rect	275	151	276	152
rect	275	157	276	158
rect	275	160	276	161
rect	275	163	276	164
rect	275	166	276	167
rect	275	169	276	170
rect	275	172	276	173
rect	275	175	276	176
rect	275	178	276	179
rect	275	184	276	185
rect	275	187	276	188
rect	275	196	276	197
rect	275	217	276	218
rect	276	7	277	8
rect	276	10	277	11
rect	276	13	277	14
rect	276	16	277	17
rect	276	19	277	20
rect	276	22	277	23
rect	276	25	277	26
rect	276	28	277	29
rect	276	31	277	32
rect	276	34	277	35
rect	276	37	277	38
rect	276	40	277	41
rect	276	43	277	44
rect	276	46	277	47
rect	276	49	277	50
rect	276	55	277	56
rect	276	61	277	62
rect	276	64	277	65
rect	276	79	277	80
rect	276	82	277	83
rect	276	85	277	86
rect	276	88	277	89
rect	276	109	277	110
rect	276	115	277	116
rect	276	118	277	119
rect	276	124	277	125
rect	276	133	277	134
rect	276	136	277	137
rect	276	139	277	140
rect	276	148	277	149
rect	276	151	277	152
rect	276	157	277	158
rect	276	160	277	161
rect	276	163	277	164
rect	276	166	277	167
rect	276	169	277	170
rect	276	172	277	173
rect	276	175	277	176
rect	276	178	277	179
rect	276	184	277	185
rect	276	187	277	188
rect	276	196	277	197
rect	276	217	277	218
rect	277	7	278	8
rect	277	10	278	11
rect	277	13	278	14
rect	277	16	278	17
rect	277	19	278	20
rect	277	22	278	23
rect	277	25	278	26
rect	277	28	278	29
rect	277	31	278	32
rect	277	34	278	35
rect	277	37	278	38
rect	277	40	278	41
rect	277	43	278	44
rect	277	46	278	47
rect	277	49	278	50
rect	277	55	278	56
rect	277	61	278	62
rect	277	64	278	65
rect	277	79	278	80
rect	277	82	278	83
rect	277	85	278	86
rect	277	88	278	89
rect	277	109	278	110
rect	277	115	278	116
rect	277	118	278	119
rect	277	124	278	125
rect	277	133	278	134
rect	277	136	278	137
rect	277	139	278	140
rect	277	148	278	149
rect	277	151	278	152
rect	277	157	278	158
rect	277	160	278	161
rect	277	163	278	164
rect	277	166	278	167
rect	277	169	278	170
rect	277	172	278	173
rect	277	175	278	176
rect	277	178	278	179
rect	277	184	278	185
rect	277	187	278	188
rect	277	196	278	197
rect	277	217	278	218
rect	278	7	279	8
rect	278	10	279	11
rect	278	13	279	14
rect	278	16	279	17
rect	278	19	279	20
rect	278	22	279	23
rect	278	25	279	26
rect	278	28	279	29
rect	278	31	279	32
rect	278	34	279	35
rect	278	37	279	38
rect	278	40	279	41
rect	278	43	279	44
rect	278	46	279	47
rect	278	49	279	50
rect	278	55	279	56
rect	278	61	279	62
rect	278	64	279	65
rect	278	79	279	80
rect	278	82	279	83
rect	278	85	279	86
rect	278	88	279	89
rect	278	109	279	110
rect	278	115	279	116
rect	278	118	279	119
rect	278	124	279	125
rect	278	133	279	134
rect	278	136	279	137
rect	278	139	279	140
rect	278	148	279	149
rect	278	151	279	152
rect	278	157	279	158
rect	278	160	279	161
rect	278	163	279	164
rect	278	166	279	167
rect	278	169	279	170
rect	278	172	279	173
rect	278	175	279	176
rect	278	178	279	179
rect	278	184	279	185
rect	278	187	279	188
rect	278	196	279	197
rect	278	217	279	218
rect	279	7	280	8
rect	279	10	280	11
rect	279	13	280	14
rect	279	16	280	17
rect	279	19	280	20
rect	279	22	280	23
rect	279	25	280	26
rect	279	28	280	29
rect	279	31	280	32
rect	279	34	280	35
rect	279	37	280	38
rect	279	40	280	41
rect	279	43	280	44
rect	279	46	280	47
rect	279	49	280	50
rect	279	55	280	56
rect	279	61	280	62
rect	279	64	280	65
rect	279	79	280	80
rect	279	82	280	83
rect	279	85	280	86
rect	279	88	280	89
rect	279	109	280	110
rect	279	115	280	116
rect	279	118	280	119
rect	279	124	280	125
rect	279	133	280	134
rect	279	136	280	137
rect	279	139	280	140
rect	279	148	280	149
rect	279	151	280	152
rect	279	157	280	158
rect	279	160	280	161
rect	279	163	280	164
rect	279	166	280	167
rect	279	169	280	170
rect	279	172	280	173
rect	279	175	280	176
rect	279	178	280	179
rect	279	184	280	185
rect	279	187	280	188
rect	279	196	280	197
rect	279	217	280	218
rect	280	7	281	8
rect	280	10	281	11
rect	280	13	281	14
rect	280	16	281	17
rect	280	19	281	20
rect	280	22	281	23
rect	280	25	281	26
rect	280	28	281	29
rect	280	31	281	32
rect	280	34	281	35
rect	280	37	281	38
rect	280	40	281	41
rect	280	43	281	44
rect	280	46	281	47
rect	280	49	281	50
rect	280	55	281	56
rect	280	61	281	62
rect	280	64	281	65
rect	280	79	281	80
rect	280	82	281	83
rect	280	85	281	86
rect	280	88	281	89
rect	280	109	281	110
rect	280	115	281	116
rect	280	118	281	119
rect	280	124	281	125
rect	280	133	281	134
rect	280	136	281	137
rect	280	139	281	140
rect	280	148	281	149
rect	280	151	281	152
rect	280	157	281	158
rect	280	160	281	161
rect	280	163	281	164
rect	280	166	281	167
rect	280	169	281	170
rect	280	172	281	173
rect	280	175	281	176
rect	280	178	281	179
rect	280	184	281	185
rect	280	187	281	188
rect	280	196	281	197
rect	280	217	281	218
rect	281	7	282	8
rect	281	10	282	11
rect	281	13	282	14
rect	281	16	282	17
rect	281	19	282	20
rect	281	22	282	23
rect	281	25	282	26
rect	281	28	282	29
rect	281	31	282	32
rect	281	34	282	35
rect	281	37	282	38
rect	281	40	282	41
rect	281	43	282	44
rect	281	46	282	47
rect	281	49	282	50
rect	281	55	282	56
rect	281	61	282	62
rect	281	64	282	65
rect	281	79	282	80
rect	281	82	282	83
rect	281	85	282	86
rect	281	88	282	89
rect	281	109	282	110
rect	281	115	282	116
rect	281	118	282	119
rect	281	124	282	125
rect	281	133	282	134
rect	281	136	282	137
rect	281	139	282	140
rect	281	148	282	149
rect	281	151	282	152
rect	281	157	282	158
rect	281	160	282	161
rect	281	163	282	164
rect	281	166	282	167
rect	281	169	282	170
rect	281	172	282	173
rect	281	175	282	176
rect	281	178	282	179
rect	281	184	282	185
rect	281	187	282	188
rect	281	196	282	197
rect	281	217	282	218
rect	282	7	283	8
rect	282	10	283	11
rect	282	13	283	14
rect	282	16	283	17
rect	282	19	283	20
rect	282	22	283	23
rect	282	25	283	26
rect	282	28	283	29
rect	282	31	283	32
rect	282	34	283	35
rect	282	37	283	38
rect	282	40	283	41
rect	282	43	283	44
rect	282	46	283	47
rect	282	49	283	50
rect	282	55	283	56
rect	282	61	283	62
rect	282	64	283	65
rect	282	79	283	80
rect	282	82	283	83
rect	282	85	283	86
rect	282	88	283	89
rect	282	109	283	110
rect	282	115	283	116
rect	282	118	283	119
rect	282	124	283	125
rect	282	133	283	134
rect	282	136	283	137
rect	282	139	283	140
rect	282	148	283	149
rect	282	151	283	152
rect	282	157	283	158
rect	282	160	283	161
rect	282	166	283	167
rect	282	169	283	170
rect	282	172	283	173
rect	282	175	283	176
rect	282	178	283	179
rect	282	184	283	185
rect	282	187	283	188
rect	282	196	283	197
rect	282	217	283	218
rect	283	7	284	8
rect	283	10	284	11
rect	283	13	284	14
rect	283	16	284	17
rect	283	19	284	20
rect	283	22	284	23
rect	283	25	284	26
rect	283	28	284	29
rect	283	31	284	32
rect	283	37	284	38
rect	283	40	284	41
rect	283	43	284	44
rect	283	46	284	47
rect	283	49	284	50
rect	283	55	284	56
rect	283	61	284	62
rect	283	64	284	65
rect	283	79	284	80
rect	283	82	284	83
rect	283	85	284	86
rect	283	115	284	116
rect	283	118	284	119
rect	283	124	284	125
rect	283	133	284	134
rect	283	136	284	137
rect	283	139	284	140
rect	283	148	284	149
rect	283	151	284	152
rect	283	157	284	158
rect	283	160	284	161
rect	283	163	284	164
rect	283	166	284	167
rect	283	169	284	170
rect	283	172	284	173
rect	283	175	284	176
rect	283	178	284	179
rect	283	184	284	185
rect	283	187	284	188
rect	284	7	285	8
rect	284	10	285	11
rect	284	13	285	14
rect	284	16	285	17
rect	284	19	285	20
rect	284	22	285	23
rect	284	25	285	26
rect	284	28	285	29
rect	284	31	285	32
rect	284	37	285	38
rect	284	40	285	41
rect	284	43	285	44
rect	284	46	285	47
rect	284	49	285	50
rect	284	55	285	56
rect	284	61	285	62
rect	284	64	285	65
rect	284	79	285	80
rect	284	82	285	83
rect	284	85	285	86
rect	284	115	285	116
rect	284	118	285	119
rect	284	124	285	125
rect	284	133	285	134
rect	284	136	285	137
rect	284	139	285	140
rect	284	148	285	149
rect	284	151	285	152
rect	284	160	285	161
rect	284	163	285	164
rect	284	166	285	167
rect	284	169	285	170
rect	284	172	285	173
rect	284	175	285	176
rect	284	178	285	179
rect	284	184	285	185
rect	284	187	285	188
rect	285	7	286	8
rect	285	10	286	11
rect	285	13	286	14
rect	285	16	286	17
rect	285	19	286	20
rect	285	22	286	23
rect	285	25	286	26
rect	285	28	286	29
rect	285	31	286	32
rect	285	37	286	38
rect	285	40	286	41
rect	285	43	286	44
rect	285	46	286	47
rect	285	49	286	50
rect	285	55	286	56
rect	285	61	286	62
rect	285	64	286	65
rect	285	79	286	80
rect	285	82	286	83
rect	285	85	286	86
rect	285	88	286	89
rect	285	109	286	110
rect	285	115	286	116
rect	285	118	286	119
rect	285	124	286	125
rect	285	133	286	134
rect	285	136	286	137
rect	285	139	286	140
rect	285	148	286	149
rect	285	151	286	152
rect	285	157	286	158
rect	285	160	286	161
rect	285	163	286	164
rect	285	166	286	167
rect	285	169	286	170
rect	285	172	286	173
rect	285	175	286	176
rect	285	178	286	179
rect	285	184	286	185
rect	285	187	286	188
rect	285	196	286	197
rect	286	7	287	8
rect	286	10	287	11
rect	286	13	287	14
rect	286	16	287	17
rect	286	19	287	20
rect	286	22	287	23
rect	286	25	287	26
rect	286	28	287	29
rect	286	31	287	32
rect	286	37	287	38
rect	286	40	287	41
rect	286	43	287	44
rect	286	46	287	47
rect	286	49	287	50
rect	286	55	287	56
rect	286	61	287	62
rect	286	64	287	65
rect	286	79	287	80
rect	286	82	287	83
rect	286	85	287	86
rect	286	88	287	89
rect	286	109	287	110
rect	286	115	287	116
rect	286	118	287	119
rect	286	124	287	125
rect	286	133	287	134
rect	286	136	287	137
rect	286	139	287	140
rect	286	148	287	149
rect	286	151	287	152
rect	286	157	287	158
rect	286	160	287	161
rect	286	163	287	164
rect	286	166	287	167
rect	286	169	287	170
rect	286	172	287	173
rect	286	175	287	176
rect	286	178	287	179
rect	286	184	287	185
rect	286	187	287	188
rect	286	196	287	197
rect	287	7	288	8
rect	287	10	288	11
rect	287	13	288	14
rect	287	16	288	17
rect	287	19	288	20
rect	287	22	288	23
rect	287	25	288	26
rect	287	28	288	29
rect	287	31	288	32
rect	287	37	288	38
rect	287	40	288	41
rect	287	43	288	44
rect	287	46	288	47
rect	287	49	288	50
rect	287	52	288	53
rect	287	55	288	56
rect	287	61	288	62
rect	287	64	288	65
rect	287	79	288	80
rect	287	82	288	83
rect	287	85	288	86
rect	287	88	288	89
rect	287	109	288	110
rect	287	115	288	116
rect	287	118	288	119
rect	287	124	288	125
rect	287	133	288	134
rect	287	136	288	137
rect	287	139	288	140
rect	287	148	288	149
rect	287	151	288	152
rect	287	157	288	158
rect	287	160	288	161
rect	287	163	288	164
rect	287	166	288	167
rect	287	169	288	170
rect	287	172	288	173
rect	287	175	288	176
rect	287	178	288	179
rect	287	184	288	185
rect	287	187	288	188
rect	287	196	288	197
rect	287	217	288	218
rect	288	7	289	8
rect	288	10	289	11
rect	288	13	289	14
rect	288	19	289	20
rect	288	22	289	23
rect	288	28	289	29
rect	288	31	289	32
rect	288	37	289	38
rect	288	40	289	41
rect	288	46	289	47
rect	288	49	289	50
rect	288	55	289	56
rect	288	64	289	65
rect	288	82	289	83
rect	288	85	289	86
rect	288	115	289	116
rect	288	124	289	125
rect	288	136	289	137
rect	288	139	289	140
rect	288	148	289	149
rect	288	151	289	152
rect	288	157	289	158
rect	288	160	289	161
rect	288	166	289	167
rect	288	169	289	170
rect	288	175	289	176
rect	288	178	289	179
rect	289	7	290	8
rect	289	10	290	11
rect	289	13	290	14
rect	289	19	290	20
rect	289	22	290	23
rect	289	28	290	29
rect	289	31	290	32
rect	289	37	290	38
rect	289	40	290	41
rect	289	46	290	47
rect	289	49	290	50
rect	289	55	290	56
rect	289	64	290	65
rect	289	82	290	83
rect	289	85	290	86
rect	289	115	290	116
rect	289	124	290	125
rect	289	136	290	137
rect	289	139	290	140
rect	289	148	290	149
rect	289	151	290	152
rect	289	157	290	158
rect	289	160	290	161
rect	289	166	290	167
rect	289	169	290	170
rect	289	175	290	176
rect	289	178	290	179
rect	290	7	291	8
rect	290	10	291	11
rect	290	13	291	14
rect	290	19	291	20
rect	290	22	291	23
rect	290	28	291	29
rect	290	31	291	32
rect	290	37	291	38
rect	290	40	291	41
rect	290	46	291	47
rect	290	49	291	50
rect	290	55	291	56
rect	290	64	291	65
rect	290	82	291	83
rect	290	85	291	86
rect	290	115	291	116
rect	290	124	291	125
rect	290	136	291	137
rect	290	139	291	140
rect	290	148	291	149
rect	290	151	291	152
rect	290	157	291	158
rect	290	160	291	161
rect	290	166	291	167
rect	290	169	291	170
rect	290	175	291	176
rect	290	178	291	179
rect	291	7	292	8
rect	291	10	292	11
rect	291	13	292	14
rect	291	19	292	20
rect	291	22	292	23
rect	291	28	292	29
rect	291	31	292	32
rect	291	37	292	38
rect	291	40	292	41
rect	291	46	292	47
rect	291	49	292	50
rect	291	55	292	56
rect	291	64	292	65
rect	291	82	292	83
rect	291	85	292	86
rect	291	115	292	116
rect	291	124	292	125
rect	291	136	292	137
rect	291	139	292	140
rect	291	148	292	149
rect	291	151	292	152
rect	291	157	292	158
rect	291	160	292	161
rect	291	166	292	167
rect	291	169	292	170
rect	291	175	292	176
rect	291	178	292	179
rect	292	7	293	8
rect	292	10	293	11
rect	292	13	293	14
rect	292	22	293	23
rect	292	28	293	29
rect	292	31	293	32
rect	292	37	293	38
rect	292	49	293	50
rect	292	64	293	65
rect	292	82	293	83
rect	292	85	293	86
rect	292	115	293	116
rect	292	124	293	125
rect	292	136	293	137
rect	292	139	293	140
rect	292	151	293	152
rect	292	160	293	161
rect	292	166	293	167
rect	292	169	293	170
rect	293	7	294	8
rect	293	10	294	11
rect	293	13	294	14
rect	293	22	294	23
rect	293	28	294	29
rect	293	31	294	32
rect	293	37	294	38
rect	293	49	294	50
rect	293	64	294	65
rect	293	79	294	80
rect	293	82	294	83
rect	293	85	294	86
rect	293	115	294	116
rect	293	124	294	125
rect	293	136	294	137
rect	293	139	294	140
rect	293	151	294	152
rect	293	160	294	161
rect	293	166	294	167
rect	293	169	294	170
rect	294	7	295	8
rect	294	10	295	11
rect	294	13	295	14
rect	294	22	295	23
rect	294	28	295	29
rect	294	31	295	32
rect	294	37	295	38
rect	294	49	295	50
rect	294	64	295	65
rect	294	79	295	80
rect	294	82	295	83
rect	294	85	295	86
rect	294	115	295	116
rect	294	124	295	125
rect	294	136	295	137
rect	294	139	295	140
rect	294	151	295	152
rect	294	160	295	161
rect	294	166	295	167
rect	294	169	295	170
rect	295	7	296	8
rect	295	10	296	11
rect	295	13	296	14
rect	295	22	296	23
rect	295	28	296	29
rect	295	31	296	32
rect	295	37	296	38
rect	295	49	296	50
rect	295	64	296	65
rect	295	85	296	86
rect	295	115	296	116
rect	295	124	296	125
rect	295	136	296	137
rect	295	139	296	140
rect	295	151	296	152
rect	295	160	296	161
rect	295	166	296	167
rect	295	169	296	170
rect	296	4	297	5
rect	296	7	297	8
rect	296	10	297	11
rect	296	13	297	14
rect	296	19	297	20
rect	296	22	297	23
rect	296	28	297	29
rect	296	31	297	32
rect	296	37	297	38
rect	296	43	297	44
rect	296	46	297	47
rect	296	49	297	50
rect	296	64	297	65
rect	296	82	297	83
rect	296	85	297	86
rect	296	115	297	116
rect	296	124	297	125
rect	296	136	297	137
rect	296	139	297	140
rect	296	148	297	149
rect	296	151	297	152
rect	296	154	297	155
rect	296	160	297	161
rect	296	166	297	167
rect	296	169	297	170
rect	297	7	298	8
rect	297	13	298	14
rect	297	28	298	29
rect	297	31	298	32
rect	297	64	298	65
rect	297	85	298	86
rect	297	115	298	116
rect	297	124	298	125
rect	297	136	298	137
rect	297	139	298	140
rect	297	166	298	167
rect	298	7	299	8
rect	298	13	299	14
rect	298	28	299	29
rect	298	31	299	32
rect	298	64	299	65
rect	298	85	299	86
rect	298	115	299	116
rect	298	124	299	125
rect	298	136	299	137
rect	298	139	299	140
rect	298	166	299	167
rect	299	7	300	8
rect	299	13	300	14
rect	299	28	300	29
rect	299	31	300	32
rect	299	64	300	65
rect	299	85	300	86
rect	299	115	300	116
rect	299	124	300	125
rect	299	136	300	137
rect	299	139	300	140
rect	299	166	300	167
rect	300	7	301	8
rect	300	13	301	14
rect	300	28	301	29
rect	300	31	301	32
rect	300	64	301	65
rect	300	85	301	86
rect	300	115	301	116
rect	300	124	301	125
rect	300	136	301	137
rect	300	139	301	140
rect	300	166	301	167
rect	301	7	302	8
rect	301	13	302	14
rect	301	28	302	29
rect	301	31	302	32
rect	301	64	302	65
rect	301	85	302	86
rect	301	115	302	116
rect	301	124	302	125
rect	301	136	302	137
rect	301	139	302	140
rect	301	166	302	167
rect	302	7	303	8
rect	302	13	303	14
rect	302	28	303	29
rect	302	31	303	32
rect	302	64	303	65
rect	302	85	303	86
rect	302	115	303	116
rect	302	124	303	125
rect	302	136	303	137
rect	302	139	303	140
rect	302	166	303	167
rect	305	88	306	89
rect	305	115	306	116
rect	305	124	306	125
rect	305	130	306	131
rect	305	139	306	140
rect	305	142	306	143
rect	306	88	307	89
rect	306	115	307	116
rect	306	124	307	125
rect	306	130	307	131
rect	306	139	307	140
rect	306	142	307	143
rect	307	4	308	5
rect	307	7	308	8
rect	307	25	308	26
rect	307	28	308	29
rect	307	82	308	83
rect	307	88	308	89
rect	307	115	308	116
rect	307	124	308	125
rect	307	130	308	131
rect	307	139	308	140
rect	307	142	308	143
rect	307	166	308	167
